//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G58), .A2(G232), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(G50), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n218), .A2(KEYINPUT1), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NOR3_X1   g0026(.A1(new_n209), .A2(new_n220), .A3(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  XNOR2_X1  g0044(.A(KEYINPUT8), .B(G58), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NOR2_X1   g0046(.A1(G20), .A2(G33), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n246), .A2(new_n247), .B1(G20), .B2(G77), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n222), .A2(G33), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT15), .B(G87), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n221), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G13), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n253), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n257), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G77), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n254), .B1(G77), .B2(new_n257), .C1(new_n259), .C2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n267), .A3(G274), .ZN(new_n268));
  INV_X1    g0068(.A(G244), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n264), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(new_n271), .B(KEYINPUT70), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G107), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(new_n274), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n211), .A3(new_n275), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n273), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n272), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n263), .B1(new_n287), .B2(G190), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(G200), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n263), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n267), .B1(new_n283), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G222), .A2(G1698), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n275), .A2(G223), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n274), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G226), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n268), .B1(new_n302), .B2(new_n270), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n293), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(G179), .B2(new_n304), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT68), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n253), .B(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G50), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n222), .B1(new_n201), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT69), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G150), .ZN(new_n313));
  INV_X1    g0113(.A(new_n247), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n245), .A2(new_n249), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n308), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n253), .B(KEYINPUT68), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(G50), .A3(new_n257), .A4(new_n261), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n260), .A2(G13), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(new_n222), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n309), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n316), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n306), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n290), .A2(new_n295), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT9), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n304), .A2(G200), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n316), .A2(KEYINPUT9), .A3(new_n318), .A4(new_n321), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OR3_X1    g0131(.A1(new_n301), .A2(new_n331), .A3(new_n303), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT71), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n328), .A2(new_n334), .A3(new_n330), .A4(new_n332), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT10), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n333), .B1(new_n336), .B2(new_n335), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n229), .A2(G1698), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n274), .B(new_n341), .C1(G226), .C2(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n273), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT13), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n268), .B1(new_n211), .B2(new_n270), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n267), .B1(new_n342), .B2(new_n343), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT13), .B1(new_n350), .B2(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n293), .B1(new_n349), .B2(new_n351), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n353), .A2(G179), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n352), .A2(G169), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT74), .B1(new_n357), .B2(KEYINPUT14), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n354), .A2(new_n359), .A3(new_n355), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n356), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n210), .A2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n247), .A2(G50), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n362), .B(new_n363), .C1(new_n296), .C2(new_n249), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n308), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT11), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n258), .A2(new_n257), .A3(G68), .A4(new_n261), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT12), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n257), .B2(G68), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n210), .A2(KEYINPUT12), .A3(G20), .A4(new_n256), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n364), .A2(KEYINPUT11), .A3(new_n308), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n367), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT73), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n367), .A2(new_n372), .A3(new_n376), .A4(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n361), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n353), .A2(G190), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT72), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n352), .B2(G200), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  AOI211_X1 g0185(.A(KEYINPUT72), .B(new_n385), .C1(new_n349), .C2(new_n351), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n326), .A2(new_n340), .A3(new_n380), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT80), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT79), .ZN(new_n392));
  INV_X1    g0192(.A(G159), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n314), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G58), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n202), .B1(new_n210), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n394), .B1(new_n396), .B2(G20), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT7), .B1(new_n274), .B2(G20), .ZN(new_n398));
  AND2_X1   g0198(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n399));
  NOR2_X1   g0199(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n283), .A2(new_n401), .A3(new_n222), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n402), .A3(G68), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n403), .A3(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT76), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT76), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n397), .A2(new_n403), .A3(new_n406), .A4(KEYINPUT16), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(G20), .B1(new_n280), .B2(new_n282), .ZN(new_n409));
  XNOR2_X1  g0209(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT77), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n401), .B(new_n412), .C1(new_n274), .C2(G20), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT78), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n280), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n279), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n282), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n222), .A2(KEYINPUT7), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n411), .A2(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n397), .B1(new_n419), .B2(new_n210), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT16), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n408), .A2(new_n422), .A3(new_n253), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n308), .A2(new_n320), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n245), .B1(new_n260), .B2(G20), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n424), .A2(new_n425), .B1(new_n320), .B2(new_n245), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n302), .A2(G1698), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n274), .B(new_n427), .C1(G223), .C2(G1698), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n267), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n268), .B1(new_n229), .B2(new_n270), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n331), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G200), .B2(new_n432), .ZN(new_n434));
  AND4_X1   g0234(.A1(KEYINPUT17), .A2(new_n423), .A3(new_n426), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n426), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n258), .B1(new_n405), .B2(new_n407), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n437), .B2(new_n422), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT17), .B1(new_n438), .B2(new_n434), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n392), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n423), .A2(new_n426), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n432), .A2(new_n293), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(G179), .B2(new_n432), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT18), .B1(new_n438), .B2(new_n444), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n423), .A2(new_n426), .A3(new_n434), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n438), .A2(KEYINPUT17), .A3(new_n434), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(KEYINPUT79), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n440), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n390), .B1(new_n391), .B2(new_n454), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n454), .A2(new_n391), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n257), .A2(G97), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n279), .A2(G1), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n317), .A2(new_n257), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(G97), .B(G107), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT6), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n467), .A2(new_n464), .A3(G107), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(G20), .B1(G77), .B2(new_n247), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n419), .B2(new_n277), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n465), .B1(new_n473), .B2(new_n253), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n267), .A2(G274), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT83), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT5), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n477), .B1(new_n478), .B2(G41), .ZN(new_n479));
  INV_X1    g0279(.A(G45), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(G41), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n478), .A2(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT83), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n476), .A2(new_n479), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G257), .B(new_n267), .C1(new_n483), .C2(new_n485), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G1698), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n491), .A2(new_n280), .A3(new_n282), .A4(G244), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT82), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n274), .A2(new_n494), .A3(G244), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(new_n275), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n490), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n280), .A2(new_n282), .A3(G250), .A4(G1698), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n497), .A2(KEYINPUT81), .A3(new_n490), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n496), .A2(new_n500), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n489), .B1(new_n506), .B2(new_n273), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n497), .A2(new_n490), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(KEYINPUT81), .B1(new_n493), .B2(new_n495), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n503), .B1(new_n499), .B2(new_n498), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n267), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n512), .A2(G190), .A3(new_n489), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n474), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n308), .A2(new_n320), .A3(new_n461), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n459), .B1(new_n515), .B2(G97), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n469), .B1(new_n467), .B2(new_n466), .ZN(new_n517));
  OAI22_X1  g0317(.A1(new_n517), .A2(new_n222), .B1(new_n296), .B2(new_n314), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n411), .A2(new_n413), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n417), .A2(new_n418), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n521), .B2(G107), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n516), .B1(new_n522), .B2(new_n258), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n507), .A2(new_n293), .ZN(new_n524));
  AOI211_X1 g0324(.A(new_n291), .B(new_n489), .C1(new_n506), .C2(new_n273), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n280), .A2(new_n282), .A3(G244), .A4(G1698), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n280), .A2(new_n282), .A3(G238), .A4(new_n275), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n273), .ZN(new_n531));
  INV_X1    g0331(.A(G250), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n480), .B2(G1), .ZN(new_n533));
  INV_X1    g0333(.A(G274), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n260), .A2(new_n534), .A3(G45), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n267), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT84), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n267), .A2(new_n533), .A3(new_n535), .A4(KEYINPUT84), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(G87), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(new_n464), .A3(new_n277), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT85), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT85), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT19), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n343), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n549), .B2(G20), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n280), .A2(new_n282), .A3(new_n222), .A4(G68), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n546), .B(new_n548), .C1(new_n249), .C2(new_n464), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(new_n253), .B1(new_n320), .B2(new_n250), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n515), .A2(G87), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n531), .A2(new_n540), .A3(G190), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n542), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n250), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n317), .A2(new_n257), .A3(new_n558), .A4(new_n462), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n320), .A2(new_n250), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n552), .A2(new_n551), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n546), .A2(new_n548), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n222), .B1(new_n562), .B2(new_n343), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n561), .B1(new_n563), .B2(new_n544), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n559), .B(new_n560), .C1(new_n564), .C2(new_n258), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n531), .A2(new_n540), .A3(new_n291), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n541), .A2(new_n293), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n557), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n514), .A2(new_n526), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n320), .A2(new_n277), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT25), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n571), .B(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n463), .B2(new_n277), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n280), .A2(new_n282), .A3(new_n222), .A4(G87), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT22), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n274), .A2(KEYINPUT22), .A3(new_n222), .A4(G87), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n222), .A2(KEYINPUT23), .A3(G107), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n529), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n579), .A2(KEYINPUT87), .B1(new_n581), .B2(new_n222), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n277), .A3(G20), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT87), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n583), .A2(new_n584), .B1(KEYINPUT23), .B2(G107), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n577), .A2(new_n578), .A3(new_n582), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT24), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n579), .A2(KEYINPUT87), .B1(new_n580), .B2(new_n277), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n583), .A2(new_n584), .B1(new_n589), .B2(G20), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT24), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n578), .A4(new_n577), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n574), .B1(new_n253), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT90), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n280), .A2(new_n282), .A3(G257), .A4(G1698), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n280), .A2(new_n282), .A3(G250), .A4(new_n275), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G294), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n273), .ZN(new_n601));
  OAI211_X1 g0401(.A(G264), .B(new_n267), .C1(new_n483), .C2(new_n485), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n487), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n385), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G190), .B2(new_n603), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n595), .A2(new_n596), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n596), .B1(new_n595), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n570), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT21), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n280), .A2(new_n282), .A3(G264), .A4(G1698), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n280), .A2(new_n282), .A3(G257), .A4(new_n275), .ZN(new_n612));
  INV_X1    g0412(.A(G303), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n274), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n273), .ZN(new_n615));
  OAI211_X1 g0415(.A(G270), .B(new_n267), .C1(new_n483), .C2(new_n485), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n487), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G169), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n462), .A2(G116), .ZN(new_n619));
  INV_X1    g0419(.A(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G20), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n259), .A2(new_n619), .B1(new_n319), .B2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n253), .A2(new_n621), .ZN(new_n623));
  AOI21_X1  g0423(.A(G20), .B1(G33), .B2(G283), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n279), .A2(G97), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT86), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT86), .B1(new_n624), .B2(new_n625), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n623), .B(KEYINPUT20), .C1(new_n627), .C2(new_n626), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n622), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n610), .B1(new_n618), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  INV_X1    g0434(.A(new_n622), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(KEYINPUT21), .A3(G169), .A4(new_n617), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n615), .A2(G179), .A3(new_n487), .A4(new_n616), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n633), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n636), .B1(G200), .B2(new_n617), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n331), .B2(new_n617), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n594), .A2(new_n253), .ZN(new_n645));
  INV_X1    g0445(.A(new_n574), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n603), .A2(G169), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n648), .B(KEYINPUT88), .C1(new_n291), .C2(new_n603), .ZN(new_n649));
  OR3_X1    g0449(.A1(new_n603), .A2(KEYINPUT88), .A3(new_n291), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT89), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n647), .A2(new_n649), .A3(KEYINPUT89), .A4(new_n650), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND4_X1   g0455(.A1(new_n458), .A2(new_n609), .A3(new_n644), .A4(new_n655), .ZN(G372));
  OAI21_X1  g0456(.A(new_n380), .B1(new_n388), .B2(new_n295), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n440), .A3(new_n453), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n448), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT93), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n338), .B2(new_n339), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n335), .A2(new_n336), .ZN(new_n662));
  INV_X1    g0462(.A(new_n333), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(KEYINPUT93), .A3(new_n337), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n324), .B1(new_n659), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT91), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n524), .B2(new_n525), .ZN(new_n669));
  OAI21_X1  g0469(.A(G169), .B1(new_n512), .B2(new_n489), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n506), .A2(new_n273), .ZN(new_n671));
  INV_X1    g0471(.A(new_n489), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(G179), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(KEYINPUT91), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n669), .A2(new_n569), .A3(new_n674), .A4(new_n523), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n474), .B1(new_n670), .B2(new_n673), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(KEYINPUT26), .A3(new_n569), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n678), .A2(new_n569), .A3(KEYINPUT92), .A4(KEYINPUT26), .ZN(new_n682));
  AND3_X1   g0482(.A1(new_n677), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n507), .A2(new_n331), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n385), .B1(new_n512), .B2(new_n489), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n523), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n678), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n595), .A2(new_n605), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT90), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n595), .A2(new_n596), .A3(new_n605), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n618), .A2(new_n632), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n639), .B1(new_n692), .B2(KEYINPUT21), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n651), .A2(new_n693), .A3(new_n633), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n687), .A2(new_n691), .A3(new_n569), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n568), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n683), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n667), .B1(new_n457), .B2(new_n697), .ZN(G369));
  OR3_X1    g0498(.A1(new_n319), .A2(KEYINPUT27), .A3(G20), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT27), .B1(new_n319), .B2(G20), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT94), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G343), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n636), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n644), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n641), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n655), .A2(new_n691), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n595), .A2(new_n703), .ZN(new_n711));
  OAI22_X1  g0511(.A1(new_n710), .A2(new_n711), .B1(new_n651), .B2(new_n703), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n651), .A2(new_n704), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n641), .A2(new_n704), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n655), .A2(new_n715), .A3(new_n691), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n207), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  NOR4_X1   g0519(.A1(new_n719), .A2(new_n260), .A3(G116), .A4(new_n544), .ZN(new_n720));
  INV_X1    g0520(.A(new_n225), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT26), .B1(new_n678), .B2(new_n569), .ZN(new_n724));
  OAI22_X1  g0524(.A1(KEYINPUT97), .A2(new_n724), .B1(new_n675), .B2(new_n676), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n669), .A2(new_n523), .A3(new_n674), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(KEYINPUT26), .A3(new_n569), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n727), .B2(KEYINPUT97), .ZN(new_n728));
  INV_X1    g0528(.A(new_n568), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n653), .A2(new_n641), .A3(new_n654), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n609), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n704), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n609), .B2(new_n694), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n677), .A2(new_n681), .A3(new_n682), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n704), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n733), .B1(KEYINPUT29), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G330), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n609), .A2(new_n644), .A3(new_n655), .A4(new_n703), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n615), .A2(new_n487), .A3(new_n616), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n601), .A2(new_n602), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n531), .A2(new_n540), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n741), .A2(G179), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n671), .A2(new_n672), .ZN(new_n745));
  OAI211_X1 g0545(.A(KEYINPUT96), .B(new_n740), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n741), .A2(G179), .A3(new_n743), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n603), .A3(new_n745), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n742), .A2(new_n743), .ZN(new_n749));
  INV_X1    g0549(.A(new_n638), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n749), .A2(new_n750), .A3(new_n507), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n746), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n753), .A2(new_n704), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT31), .B1(new_n753), .B2(new_n704), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n738), .B1(new_n739), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n737), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n723), .B1(new_n761), .B2(G1), .ZN(G364));
  INV_X1    g0562(.A(new_n719), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n255), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n260), .B1(new_n764), .B2(G45), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n709), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G330), .B2(new_n707), .ZN(new_n769));
  INV_X1    g0569(.A(new_n767), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n221), .B1(G20), .B2(new_n293), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT101), .Z(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT102), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n718), .A2(new_n274), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT100), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n225), .A2(G45), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n243), .B2(G45), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n718), .A2(new_n283), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n782), .A2(G355), .B1(new_n620), .B2(new_n718), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n779), .A2(new_n781), .B1(new_n784), .B2(KEYINPUT99), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n784), .A2(KEYINPUT99), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n777), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n222), .A2(new_n291), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n331), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n291), .A2(new_n385), .A3(G190), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n790), .A2(G326), .B1(G294), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n788), .A2(G190), .A3(new_n385), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G322), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n788), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n274), .B1(new_n799), .B2(G311), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n793), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n789), .A2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(G317), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT33), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(KEYINPUT33), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n222), .A2(G179), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n808), .A2(new_n331), .A3(G200), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(G190), .A3(G200), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n806), .B1(new_n807), .B2(new_n809), .C1(new_n613), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n808), .A2(new_n797), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(KEYINPUT103), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(KEYINPUT103), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n801), .B(new_n811), .C1(G329), .C2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n802), .A2(G68), .B1(G97), .B2(new_n792), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n812), .A2(new_n393), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n819), .B1(KEYINPUT32), .B2(new_n821), .C1(new_n543), .C2(new_n810), .ZN(new_n822));
  INV_X1    g0622(.A(new_n809), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n821), .A2(KEYINPUT32), .B1(G107), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n790), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n309), .B2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n274), .B1(new_n798), .B2(new_n296), .C1(new_n395), .C2(new_n794), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n822), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n818), .A2(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n770), .B(new_n787), .C1(new_n774), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n773), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n830), .B1(new_n707), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n769), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(G396));
  NOR2_X1   g0634(.A1(new_n295), .A2(new_n704), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n288), .A2(new_n289), .B1(new_n263), .B2(new_n704), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(new_n837), .B2(new_n295), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n736), .B(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n767), .B1(new_n839), .B2(new_n760), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n760), .B2(new_n839), .ZN(new_n841));
  INV_X1    g0641(.A(new_n774), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n795), .A2(G143), .B1(new_n799), .B2(G159), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  INV_X1    g0644(.A(new_n802), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n843), .B1(new_n825), .B2(new_n844), .C1(new_n313), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT34), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n817), .A2(G132), .ZN(new_n850));
  INV_X1    g0650(.A(new_n792), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n851), .A2(new_n395), .B1(new_n810), .B2(new_n309), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n283), .B(new_n852), .C1(G68), .C2(new_n823), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n817), .A2(G311), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n810), .A2(new_n277), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n809), .A2(new_n543), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(G283), .C2(new_n802), .ZN(new_n858));
  INV_X1    g0658(.A(G294), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n283), .B1(new_n794), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n860), .B1(G116), .B2(new_n799), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n790), .A2(G303), .B1(G97), .B2(new_n792), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n855), .A2(new_n858), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n842), .B1(new_n854), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n842), .A2(new_n772), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n767), .B1(G77), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n838), .B2(new_n772), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n841), .A2(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n764), .A2(new_n260), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n755), .B1(new_n753), .B2(new_n704), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n753), .A2(new_n704), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n871), .B1(KEYINPUT31), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n739), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n458), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT107), .Z(new_n876));
  AND3_X1   g0676(.A1(new_n292), .A2(new_n263), .A3(new_n294), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n703), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n836), .B2(new_n877), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n380), .B(new_n389), .C1(new_n378), .C2(new_n703), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n379), .B(new_n704), .C1(new_n388), .C2(new_n361), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n882), .A2(new_n874), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n702), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n397), .A2(new_n403), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n408), .B(new_n308), .C1(KEYINPUT16), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n426), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n454), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n449), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n887), .A2(new_n426), .B1(new_n444), .B2(new_n885), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n441), .A2(new_n445), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n441), .A2(new_n702), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT37), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .A4(new_n449), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n889), .A2(KEYINPUT38), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT38), .B1(new_n889), .B2(new_n897), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n884), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n882), .A2(new_n874), .ZN(new_n901));
  XOR2_X1   g0701(.A(KEYINPUT105), .B(KEYINPUT38), .Z(new_n902));
  NAND2_X1  g0702(.A1(new_n446), .A2(new_n447), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n435), .A2(new_n439), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT106), .B1(new_n435), .B2(new_n439), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n894), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n893), .A2(new_n894), .A3(new_n449), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n896), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n902), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n454), .A2(new_n888), .B1(new_n896), .B2(new_n892), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT38), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n901), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n900), .B1(new_n916), .B2(new_n883), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n738), .B1(new_n876), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n876), .B2(new_n917), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  INV_X1    g0720(.A(new_n902), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n451), .A2(new_n905), .A3(new_n452), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n907), .A2(new_n448), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n894), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n921), .B1(new_n925), .B2(new_n911), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n920), .B1(new_n898), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n889), .A2(new_n897), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT38), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(KEYINPUT39), .A3(new_n915), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n380), .A2(new_n704), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n927), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n915), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n880), .A2(new_n881), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n703), .B(new_n838), .C1(new_n683), .C2(new_n696), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n835), .B(KEYINPUT104), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n934), .A2(new_n939), .B1(new_n903), .B2(new_n885), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n933), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n667), .B1(new_n737), .B2(new_n457), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n870), .B1(new_n919), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n919), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n620), .B(new_n224), .C1(new_n471), .C2(KEYINPUT35), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(KEYINPUT35), .B2(new_n471), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT36), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n721), .B(G77), .C1(new_n395), .C2(new_n210), .ZN(new_n949));
  INV_X1    g0749(.A(G68), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(G50), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(G1), .A3(new_n255), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n945), .A2(new_n948), .A3(new_n952), .ZN(G367));
  NAND2_X1  g0753(.A1(new_n523), .A2(new_n704), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n726), .A2(new_n704), .B1(new_n687), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n716), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT42), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n526), .B1(new_n955), .B2(new_n655), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n703), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n554), .A2(new_n555), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n704), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n569), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n729), .A2(new_n961), .A3(new_n704), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n965), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n967), .B(new_n970), .Z(new_n971));
  NOR2_X1   g0771(.A1(new_n713), .A2(new_n955), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n719), .B(KEYINPUT41), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n716), .A2(new_n714), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n955), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT44), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n975), .A2(new_n955), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT45), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n980), .A2(new_n709), .A3(new_n712), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n977), .A2(new_n713), .A3(new_n979), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n716), .B1(new_n712), .B2(new_n715), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n709), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n761), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n974), .B1(new_n988), .B2(new_n761), .ZN(new_n989));
  INV_X1    g0789(.A(new_n765), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n973), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n776), .ZN(new_n992));
  INV_X1    g0792(.A(new_n779), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n992), .B1(new_n207), .B2(new_n250), .C1(new_n993), .C2(new_n235), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n994), .A2(new_n767), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n283), .B1(new_n798), .B2(new_n807), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n794), .A2(new_n613), .B1(new_n812), .B2(new_n803), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n810), .A2(new_n620), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n997), .C1(KEYINPUT46), .C2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(KEYINPUT46), .B2(new_n998), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n845), .A2(new_n859), .B1(new_n809), .B2(new_n464), .ZN(new_n1001));
  INV_X1    g0801(.A(G311), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n825), .A2(new_n1002), .B1(new_n277), .B2(new_n851), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n851), .A2(new_n950), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G150), .B2(new_n795), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT108), .Z(new_n1007));
  INV_X1    g0807(.A(G143), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1008), .A2(new_n825), .B1(new_n845), .B2(new_n393), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n274), .B1(new_n812), .B2(new_n844), .C1(new_n309), .C2(new_n798), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n809), .A2(new_n296), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n810), .A2(new_n395), .ZN(new_n1012));
  NOR4_X1   g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1004), .B1(new_n1007), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n995), .B1(new_n831), .B2(new_n965), .C1(new_n1016), .C2(new_n842), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n991), .A2(new_n1017), .ZN(G387));
  OR2_X1    g0818(.A1(new_n712), .A2(new_n831), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n782), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n544), .A2(G116), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(G107), .B2(new_n207), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n232), .A2(new_n480), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT110), .Z(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n480), .C1(new_n950), .C2(new_n296), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n245), .B2(G50), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n246), .A2(KEYINPUT50), .A3(new_n309), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1025), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n993), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1022), .B1(new_n1024), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n767), .B1(new_n1031), .B2(new_n777), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n795), .A2(G317), .B1(new_n799), .B2(G303), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n790), .A2(G322), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n1002), .C2(new_n845), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n807), .B2(new_n851), .C1(new_n859), .C2(new_n810), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT49), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n809), .A2(new_n620), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n274), .B(new_n1043), .C1(G326), .C2(new_n813), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n845), .A2(new_n245), .B1(new_n296), .B2(new_n810), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n851), .A2(new_n250), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(KEYINPUT111), .B(G150), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n798), .A2(new_n950), .B1(new_n812), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n283), .B(new_n1050), .C1(G50), .C2(new_n795), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n790), .A2(G159), .B1(new_n823), .B2(G97), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1048), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1032), .B1(new_n1054), .B2(new_n774), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n985), .A2(new_n990), .B1(new_n1019), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n986), .A2(new_n719), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n761), .A2(new_n985), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(G393));
  AOI21_X1  g0859(.A(new_n763), .B1(new_n983), .B2(new_n987), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n981), .A2(new_n982), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n986), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n955), .A2(new_n773), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n992), .B1(new_n464), .B2(new_n207), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n240), .B2(new_n779), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n825), .A2(new_n313), .B1(new_n393), .B2(new_n794), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n283), .B(new_n857), .C1(new_n246), .C2(new_n799), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n851), .A2(new_n296), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G50), .B2(new_n802), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n810), .A2(new_n210), .B1(new_n812), .B2(new_n1008), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT112), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n845), .A2(new_n613), .B1(new_n809), .B2(new_n277), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n274), .B1(new_n813), .B2(G322), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n859), .B2(new_n798), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n851), .A2(new_n620), .B1(new_n810), .B2(new_n807), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G317), .A2(new_n790), .B1(new_n795), .B2(G311), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1072), .A2(new_n1074), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1066), .B(new_n770), .C1(new_n774), .C2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1064), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1061), .B2(new_n765), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1063), .A2(new_n1086), .ZN(G390));
  AOI21_X1  g0887(.A(new_n738), .B1(new_n873), .B2(new_n739), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n936), .B1(new_n1089), .B2(new_n879), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n837), .A2(new_n295), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n835), .B1(new_n732), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n738), .B(new_n879), .C1(new_n739), .C2(new_n758), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n935), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n739), .A2(new_n758), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(G330), .A3(new_n838), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1097), .A2(new_n936), .B1(new_n882), .B2(new_n1088), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n938), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n736), .B2(new_n838), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1098), .A2(KEYINPUT115), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT115), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1088), .A2(new_n882), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n1093), .B2(new_n935), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n937), .A2(new_n938), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1095), .B1(new_n1101), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n455), .A2(new_n456), .A3(new_n1088), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n667), .B(new_n1108), .C1(new_n737), .C2(new_n457), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1100), .A2(new_n936), .B1(new_n380), .B2(new_n704), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n898), .A2(new_n899), .A3(new_n920), .ZN(new_n1115));
  AOI21_X1  g0915(.A(KEYINPUT39), .B1(new_n913), .B2(new_n915), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n932), .B(KEYINPUT114), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n898), .B2(new_n926), .C1(new_n1092), .C2(new_n936), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1117), .A2(new_n1119), .A3(new_n1094), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1103), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1113), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1111), .B(new_n1112), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n719), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n771), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n767), .B1(new_n246), .B2(new_n865), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n816), .A2(new_n859), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n283), .B1(new_n798), .B2(new_n464), .C1(new_n620), .C2(new_n794), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n950), .A2(new_n809), .B1(new_n810), .B2(new_n543), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1070), .B1(G283), .B2(new_n790), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n277), .C2(new_n845), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n810), .A2(new_n1049), .ZN(new_n1134));
  XOR2_X1   g0934(.A(new_n1134), .B(KEYINPUT53), .Z(new_n1135));
  NAND2_X1  g0935(.A1(new_n817), .A2(G125), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n845), .A2(new_n844), .B1(new_n809), .B2(new_n309), .ZN(new_n1137));
  INV_X1    g0937(.A(G128), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n825), .A2(new_n1138), .B1(new_n393), .B2(new_n851), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n274), .B1(new_n798), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G132), .B2(new_n795), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1133), .B1(new_n1135), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1127), .B1(new_n774), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1122), .A2(new_n990), .B1(new_n1126), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1125), .A2(new_n1147), .ZN(G378));
  NAND3_X1  g0948(.A1(new_n661), .A2(new_n665), .A3(new_n325), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n323), .A2(new_n885), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1150), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n661), .A2(new_n665), .A3(new_n325), .A4(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n925), .A2(new_n911), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(new_n902), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n1159));
  OAI21_X1  g0959(.A(KEYINPUT40), .B1(new_n1159), .B2(new_n901), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n738), .B(new_n1157), .C1(new_n1160), .C2(new_n900), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1157), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n917), .B2(G330), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n941), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n901), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n898), .B2(new_n926), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1166), .A2(KEYINPUT40), .B1(new_n934), .B2(new_n884), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1157), .B1(new_n1167), .B2(new_n738), .ZN(new_n1168));
  AND2_X1   g0968(.A1(new_n933), .A2(new_n940), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n917), .A2(G330), .A3(new_n1162), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1164), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1157), .A2(new_n771), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n767), .B1(G50), .B2(new_n865), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n274), .A2(G41), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n309), .B1(G33), .B2(G41), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n825), .A2(new_n620), .B1(new_n809), .B2(new_n395), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G97), .B2(new_n802), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1175), .B1(new_n798), .B2(new_n250), .C1(new_n277), .C2(new_n794), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n810), .A2(new_n296), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1180), .A2(new_n1005), .A3(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1179), .B(new_n1182), .C1(new_n807), .C2(new_n816), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1177), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT117), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n802), .A2(G132), .B1(new_n799), .B2(G137), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT118), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n794), .A2(new_n1138), .B1(new_n810), .B2(new_n1141), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT119), .Z(new_n1191));
  AOI22_X1  g0991(.A1(new_n790), .A2(G125), .B1(G150), .B2(new_n792), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OR2_X1    g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n823), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n813), .C2(G124), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .A4(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1187), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1174), .B1(new_n1201), .B2(new_n774), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1172), .A2(new_n990), .B1(new_n1173), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1103), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n932), .B1(new_n1105), .B2(new_n935), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n927), .B2(new_n931), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n675), .A2(KEYINPUT97), .A3(new_n676), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n724), .A2(KEYINPUT97), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n727), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n609), .A2(new_n730), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n568), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n703), .B(new_n1091), .C1(new_n1209), .C2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n936), .B1(new_n1212), .B2(new_n878), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1118), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1213), .A2(new_n1159), .A3(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1204), .B1(new_n1206), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1117), .A2(new_n1119), .A3(new_n1094), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n1107), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n1164), .A2(new_n1171), .B1(new_n1218), .B2(new_n1110), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n719), .B1(new_n1219), .B2(KEYINPUT57), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT120), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1164), .A2(new_n1221), .A3(new_n1171), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(new_n1218), .B2(new_n1110), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1168), .A2(new_n1169), .A3(KEYINPUT120), .A4(new_n1170), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1203), .B1(new_n1220), .B2(new_n1226), .ZN(G375));
  AND2_X1   g1027(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT115), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1104), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1092), .A2(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1109), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n974), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n1111), .A3(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1234), .B(KEYINPUT121), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n936), .A2(new_n771), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n767), .B1(G68), .B2(new_n865), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n790), .A2(G132), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n393), .B2(new_n810), .C1(new_n845), .C2(new_n1141), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n816), .A2(new_n1138), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n274), .B1(new_n798), .B2(new_n313), .C1(new_n844), .C2(new_n794), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n851), .A2(new_n309), .B1(new_n809), .B2(new_n395), .ZN(new_n1242));
  OR4_X1    g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n816), .A2(new_n613), .B1(new_n464), .B2(new_n810), .ZN(new_n1244));
  XOR2_X1   g1044(.A(new_n1244), .B(KEYINPUT122), .Z(new_n1245));
  OAI22_X1  g1045(.A1(new_n620), .A2(new_n845), .B1(new_n825), .B2(new_n859), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n283), .B1(new_n798), .B2(new_n277), .C1(new_n807), .C2(new_n794), .ZN(new_n1247));
  OR4_X1    g1047(.A1(new_n1011), .A2(new_n1246), .A3(new_n1047), .A4(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1243), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1237), .B1(new_n1249), .B2(new_n774), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1107), .A2(new_n990), .B1(new_n1236), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1235), .A2(new_n1251), .ZN(G381));
  NOR3_X1   g1052(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n1253), .B(KEYINPUT123), .Z(new_n1254));
  NOR2_X1   g1054(.A1(new_n1063), .A2(new_n1086), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n991), .A3(new_n1017), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1254), .A2(new_n1256), .A3(G381), .A4(G378), .ZN(new_n1257));
  INV_X1    g1057(.A(G375), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(G407));
  AND2_X1   g1059(.A1(new_n1125), .A2(new_n1147), .ZN(new_n1260));
  INV_X1    g1060(.A(G213), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G343), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1258), .A2(new_n1260), .A3(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(G407), .A2(G213), .A3(new_n1263), .ZN(G409));
  NAND2_X1  g1064(.A1(new_n1262), .A2(G2897), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1111), .A2(KEYINPUT60), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1232), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1268), .A2(KEYINPUT60), .A3(new_n1109), .A4(new_n1095), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n719), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G384), .B1(new_n1272), .B2(new_n1251), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1270), .B1(new_n1266), .B2(new_n1232), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1251), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1265), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT124), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1272), .A2(G384), .A3(new_n1251), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1275), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(G2897), .A4(new_n1262), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1278), .A2(new_n1279), .A3(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G378), .B(new_n1203), .C1(new_n1220), .C2(new_n1226), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1222), .A2(new_n990), .A3(new_n1225), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1173), .A2(new_n1202), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1218), .A2(new_n1110), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1172), .A2(new_n1233), .A3(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1285), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1260), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1262), .B1(new_n1284), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1279), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1292));
  OR3_X1    g1092(.A1(new_n1283), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(G393), .B(new_n833), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1256), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1255), .B1(new_n991), .B2(new_n1017), .ZN(new_n1296));
  OAI211_X1 g1096(.A(KEYINPUT125), .B(new_n1294), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(G387), .A2(G390), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1294), .A2(KEYINPUT125), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(KEYINPUT125), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1298), .A2(new_n1256), .A3(new_n1299), .A4(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1297), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n1262), .B(new_n1304), .C1(new_n1284), .C2(new_n1290), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT63), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1304), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1291), .A2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1293), .A2(new_n1303), .A3(new_n1306), .A4(new_n1310), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1302), .B1(new_n1312), .B2(new_n1291), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1305), .B2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1308), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1313), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1311), .B1(new_n1320), .B2(new_n1321), .ZN(G405));
  NAND2_X1  g1122(.A1(G375), .A2(new_n1260), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1323), .A2(KEYINPUT127), .A3(new_n1284), .ZN(new_n1324));
  AOI21_X1  g1124(.A(KEYINPUT127), .B1(new_n1323), .B2(new_n1284), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1307), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1284), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1329));
  OAI211_X1 g1129(.A(new_n1329), .B(new_n719), .C1(KEYINPUT57), .C2(new_n1219), .ZN(new_n1330));
  AOI21_X1  g1130(.A(G378), .B1(new_n1330), .B2(new_n1203), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1327), .B1(new_n1328), .B2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1323), .A2(KEYINPUT127), .A3(new_n1284), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1304), .A3(new_n1333), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1326), .A2(new_n1321), .A3(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1321), .B1(new_n1326), .B2(new_n1334), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(G402));
endmodule


