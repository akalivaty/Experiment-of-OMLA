//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G122), .Z(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT8), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G104), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n192), .A2(G107), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n193), .A2(new_n196), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(G107), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n195), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(G101), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n199), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G119), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G116), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n204), .A2(KEYINPUT65), .A3(G119), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT2), .A2(G113), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT2), .ZN(new_n213));
  INV_X1    g027(.A(G113), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n211), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n210), .A2(new_n217), .A3(KEYINPUT66), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT5), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n214), .B1(new_n205), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n203), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n210), .A2(new_n217), .A3(KEYINPUT66), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT66), .B1(new_n210), .B2(new_n217), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n226), .B(new_n203), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n191), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT0), .B(G128), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G125), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n235), .A2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n233), .A2(G143), .ZN(new_n245));
  OAI211_X1 g059(.A(G128), .B(new_n243), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G128), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n234), .B(new_n236), .C1(KEYINPUT1), .C2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n242), .B1(new_n249), .B2(G125), .ZN(new_n250));
  INV_X1    g064(.A(G224), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT7), .B1(new_n251), .B2(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n252), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n242), .B(new_n254), .C1(new_n249), .C2(G125), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n232), .A2(new_n257), .A3(KEYINPUT84), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT84), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n226), .B1(new_n228), .B2(new_n229), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n199), .A2(new_n202), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n190), .B1(new_n262), .B2(new_n230), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n263), .B2(new_n256), .ZN(new_n264));
  INV_X1    g078(.A(new_n189), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n210), .A2(new_n217), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n220), .B2(new_n221), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n193), .A2(new_n196), .A3(new_n198), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G101), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n271), .A3(G101), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n230), .B(new_n265), .C1(new_n267), .C2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n258), .A2(new_n264), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n275), .A2(KEYINPUT85), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT85), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n230), .B1(new_n267), .B2(new_n273), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n189), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT6), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n251), .A2(G953), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n250), .B(new_n283), .Z(new_n284));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(KEYINPUT82), .A3(new_n189), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT6), .A3(new_n274), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT82), .B1(new_n280), .B2(new_n189), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n285), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n288), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n274), .A2(KEYINPUT6), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT83), .A4(new_n286), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n282), .B(new_n284), .C1(new_n289), .C2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n188), .B1(new_n279), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT86), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n275), .A2(new_n276), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT85), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n275), .A2(KEYINPUT85), .A3(new_n276), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n289), .A2(new_n292), .ZN(new_n301));
  INV_X1    g115(.A(new_n282), .ZN(new_n302));
  INV_X1    g116(.A(new_n284), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n187), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n294), .A2(new_n295), .A3(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n300), .A2(KEYINPUT86), .A3(new_n187), .A4(new_n304), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G140), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n312), .A2(G227), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n246), .A2(new_n248), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n246), .A2(KEYINPUT67), .A3(new_n248), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n317), .A2(KEYINPUT10), .A3(new_n318), .A4(new_n203), .ZN(new_n319));
  INV_X1    g133(.A(new_n241), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n270), .A2(new_n320), .A3(new_n272), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n249), .A2(new_n203), .A3(KEYINPUT78), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n315), .B2(new_n261), .ZN(new_n326));
  AOI21_X1  g140(.A(KEYINPUT10), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT11), .ZN(new_n329));
  INV_X1    g143(.A(G134), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(G137), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(G137), .ZN(new_n332));
  INV_X1    g146(.A(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT11), .A3(G134), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G131), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n334), .A3(new_n337), .A4(new_n332), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n323), .A2(new_n328), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT12), .B1(new_n339), .B2(KEYINPUT79), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n324), .A2(new_n326), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n315), .A2(new_n261), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n344), .B1(new_n347), .B2(new_n339), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n324), .A2(new_n326), .B1(new_n315), .B2(new_n261), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n349), .A2(new_n340), .A3(new_n343), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n341), .B(new_n342), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(new_n339), .A3(new_n344), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n343), .B1(new_n349), .B2(new_n340), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n342), .B1(new_n355), .B2(new_n341), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n314), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n340), .B1(new_n323), .B2(new_n328), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n322), .A2(new_n327), .A3(new_n339), .ZN(new_n359));
  OR3_X1    g173(.A1(new_n358), .A2(new_n359), .A3(new_n314), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(G469), .A3(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n314), .B1(new_n358), .B2(new_n359), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n359), .B2(new_n314), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n355), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n359), .A2(new_n363), .A3(new_n314), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G469), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT73), .B(G902), .Z(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n276), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n361), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G221), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT9), .B(G234), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n376), .B2(new_n276), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(G237), .A2(G953), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(G143), .A3(G214), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G143), .B1(new_n380), .B2(G214), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G237), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n312), .A3(G214), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n235), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n337), .A3(new_n381), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G125), .B(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT16), .ZN(new_n391));
  INV_X1    g205(.A(G125), .ZN(new_n392));
  OR3_X1    g206(.A1(new_n392), .A2(KEYINPUT16), .A3(G140), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(G146), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT88), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(KEYINPUT19), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n390), .B2(new_n397), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n389), .B(new_n394), .C1(new_n399), .C2(G146), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n387), .A2(new_n381), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT87), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT18), .B(G131), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT18), .A2(G131), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n387), .A2(KEYINPUT87), .A3(new_n404), .A4(new_n381), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n390), .B(new_n233), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(G113), .B(G122), .Z(new_n409));
  XOR2_X1   g223(.A(KEYINPUT89), .B(G104), .Z(new_n410));
  XOR2_X1   g224(.A(new_n409), .B(new_n410), .Z(new_n411));
  NOR2_X1   g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n384), .A2(new_n413), .A3(new_n388), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n391), .A2(new_n393), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n233), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n401), .A2(KEYINPUT17), .A3(G131), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n414), .A2(new_n416), .A3(new_n394), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n407), .A3(new_n411), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n418), .A2(new_n407), .A3(KEYINPUT90), .A4(new_n411), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n412), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G475), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n276), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT20), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n422), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n408), .A2(new_n411), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT20), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n424), .A4(new_n276), .ZN(new_n431));
  INV_X1    g245(.A(new_n427), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n411), .B1(new_n418), .B2(new_n407), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n276), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n426), .A2(new_n431), .B1(new_n434), .B2(G475), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n204), .A2(G122), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n195), .B1(new_n436), .B2(KEYINPUT14), .ZN(new_n437));
  XNOR2_X1  g251(.A(G116), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n235), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n247), .A2(G143), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT94), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT94), .B1(new_n440), .B2(new_n441), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n330), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n443), .A2(new_n330), .A3(new_n444), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n439), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n441), .B1(new_n449), .B2(new_n440), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n440), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT93), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT93), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n453), .A3(new_n440), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(new_n330), .ZN(new_n456));
  XNOR2_X1  g270(.A(KEYINPUT91), .B(G107), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n438), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n445), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n448), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G217), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n375), .A2(new_n461), .A3(G953), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n448), .B(new_n462), .C1(new_n456), .C2(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n369), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n467), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT95), .B(G952), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G953), .ZN(new_n473));
  NAND2_X1  g287(.A1(G234), .A2(G237), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n369), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n477), .A2(G953), .A3(new_n474), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n435), .A2(new_n471), .A3(new_n481), .ZN(new_n482));
  NOR4_X1   g296(.A1(new_n308), .A2(new_n310), .A3(new_n379), .A4(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n461), .B1(new_n369), .B2(G234), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n416), .A2(new_n394), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n247), .B(G119), .C1(KEYINPUT75), .C2(KEYINPUT23), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n487), .B1(new_n207), .B2(G128), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n207), .B2(G128), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G119), .B(G128), .ZN(new_n492));
  XOR2_X1   g306(.A(KEYINPUT24), .B(G110), .Z(new_n493));
  AOI22_X1  g307(.A1(new_n491), .A2(G110), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n485), .A2(new_n494), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n491), .A2(G110), .B1(new_n492), .B2(new_n493), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n390), .A2(new_n233), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n394), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT22), .B(G137), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n500), .B(new_n501), .Z(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n498), .A3(new_n502), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT25), .A3(new_n369), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT25), .B1(new_n506), .B2(new_n369), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n484), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n484), .A2(G902), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT76), .Z(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT77), .Z(new_n515));
  NOR2_X1   g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n332), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n330), .A2(G137), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n520), .A2(new_n338), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n317), .A2(new_n521), .A3(new_n318), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n241), .B1(new_n338), .B2(new_n336), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n267), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT71), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n525), .ZN(new_n532));
  AND4_X1   g346(.A1(new_n520), .A2(new_n246), .A3(new_n338), .A4(new_n248), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n267), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT28), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(KEYINPUT26), .B(G101), .Z(new_n538));
  NAND2_X1  g352(.A1(new_n380), .A2(G210), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT31), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n522), .A2(new_n524), .A3(new_n546), .A4(KEYINPUT30), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT30), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT30), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n523), .B2(new_n533), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT68), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n547), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n267), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n525), .A3(new_n542), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n532), .B1(new_n552), .B2(new_n553), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT70), .A3(new_n542), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n545), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n545), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n544), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT32), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n544), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT70), .B1(new_n558), .B2(new_n542), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT30), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT68), .A3(new_n550), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n267), .B1(new_n570), .B2(new_n547), .ZN(new_n571));
  NOR4_X1   g385(.A1(new_n571), .A2(new_n556), .A3(new_n532), .A4(new_n543), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT31), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n567), .B1(new_n573), .B2(new_n561), .ZN(new_n574));
  INV_X1    g388(.A(new_n565), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT32), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT72), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n529), .B2(new_n530), .ZN(new_n579));
  INV_X1    g393(.A(new_n530), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(KEYINPUT72), .A3(new_n528), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n267), .B1(new_n522), .B2(new_n524), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n532), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT28), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n579), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n542), .A2(KEYINPUT29), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n369), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT74), .ZN(new_n588));
  INV_X1    g402(.A(new_n558), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n543), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT29), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n590), .B(new_n591), .C1(new_n537), .C2(new_n543), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n587), .A2(KEYINPUT74), .ZN(new_n594));
  OAI21_X1  g408(.A(G472), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n517), .B1(new_n577), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n483), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n599));
  INV_X1    g413(.A(new_n379), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n516), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n574), .B2(new_n477), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n563), .A2(new_n565), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n599), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n602), .A2(new_n603), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n606), .A2(KEYINPUT96), .A3(new_n516), .A4(new_n600), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n279), .A2(new_n293), .A3(new_n188), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n187), .B1(new_n300), .B2(new_n304), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n309), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT97), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n426), .A2(new_n431), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n434), .A2(G475), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n615), .B1(new_n463), .B2(KEYINPUT98), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n464), .A2(new_n465), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n464), .B2(new_n465), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n477), .A2(new_n468), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n467), .A2(new_n468), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n613), .A2(new_n614), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n294), .A2(new_n305), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n309), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n612), .A2(new_n481), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n608), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT99), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT34), .B(G104), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  NAND2_X1  g446(.A1(new_n435), .A2(new_n470), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n612), .A2(new_n481), .A3(new_n626), .A4(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n608), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NOR2_X1   g453(.A1(new_n503), .A2(KEYINPUT36), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n499), .B(new_n640), .Z(new_n641));
  INV_X1    g455(.A(new_n513), .ZN(new_n642));
  OR2_X1    g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n510), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n604), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n483), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  AOI21_X1  g463(.A(new_n625), .B1(new_n624), .B2(new_n309), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT97), .B(new_n310), .C1(new_n294), .C2(new_n305), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n379), .B1(new_n577), .B2(new_n595), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n476), .B1(new_n478), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n634), .A2(KEYINPUT100), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n658), .B1(new_n633), .B2(new_n655), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n645), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  NOR4_X1   g477(.A1(new_n644), .A2(new_n471), .A3(new_n435), .A4(new_n310), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT102), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n655), .B(KEYINPUT39), .Z(new_n666));
  NAND2_X1  g480(.A1(new_n600), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n665), .B1(KEYINPUT40), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n308), .B(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n671));
  AOI211_X1 g485(.A(new_n572), .B(new_n568), .C1(new_n543), .C2(new_n583), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n672), .B2(G902), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n577), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR4_X1   g489(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n235), .ZN(G45));
  NAND2_X1  g491(.A1(new_n623), .A2(new_n656), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n645), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n652), .A2(new_n653), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  AOI21_X1  g495(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n574), .A2(KEYINPUT32), .A3(new_n575), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n595), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n367), .A2(new_n369), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G469), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n370), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n377), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n684), .A2(new_n516), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n627), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT41), .B(G113), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT103), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n690), .B(new_n692), .ZN(G15));
  NOR2_X1   g507(.A1(new_n689), .A2(new_n635), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n204), .ZN(G18));
  NOR2_X1   g509(.A1(new_n482), .A2(new_n645), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n652), .A2(new_n684), .A3(new_n688), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  NOR2_X1   g512(.A1(new_n471), .A2(new_n435), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n560), .A2(new_n562), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n585), .A2(new_n543), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n565), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n702), .A2(new_n602), .A3(new_n516), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n687), .A2(new_n377), .A3(new_n480), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n652), .A2(new_n699), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND3_X1  g520(.A1(new_n702), .A2(new_n602), .A3(new_n644), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n623), .B2(new_n656), .ZN(new_n709));
  AOI22_X1  g523(.A1(new_n619), .A2(new_n620), .B1(new_n468), .B2(new_n467), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n435), .A2(new_n710), .A3(KEYINPUT104), .A4(new_n655), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n707), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n652), .A3(new_n688), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n310), .B1(new_n306), .B2(new_n307), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n684), .A2(new_n717), .A3(new_n516), .A4(new_n600), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n718), .B2(new_n712), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n310), .B(new_n379), .C1(new_n306), .C2(new_n307), .ZN(new_n720));
  INV_X1    g534(.A(new_n712), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n596), .A3(KEYINPUT42), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  NOR2_X1   g538(.A1(new_n718), .A2(new_n660), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n330), .ZN(G36));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT46), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n357), .A2(KEYINPUT45), .A3(new_n360), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n357), .A2(KEYINPUT105), .A3(KEYINPUT45), .A4(new_n360), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT45), .B1(new_n357), .B2(new_n360), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n368), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n727), .B(new_n728), .C1(new_n736), .C2(new_n371), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n371), .B1(new_n733), .B2(new_n735), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT106), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n739));
  INV_X1    g553(.A(new_n370), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n378), .A3(new_n666), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n613), .A2(new_n614), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n710), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n606), .A2(new_n749), .A3(new_n645), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n750), .A2(KEYINPUT44), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n717), .B1(new_n750), .B2(KEYINPUT44), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n742), .A2(KEYINPUT107), .A3(new_n378), .A4(new_n666), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n745), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  INV_X1    g570(.A(new_n717), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n757), .A2(new_n684), .A3(new_n516), .A4(new_n678), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n742), .A2(new_n378), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n759), .B1(new_n742), .B2(new_n378), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  NOR2_X1   g577(.A1(new_n749), .A2(new_n475), .ZN(new_n764));
  INV_X1    g578(.A(new_n688), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n309), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n670), .A2(new_n703), .A3(new_n764), .A4(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT50), .Z(new_n768));
  NOR2_X1   g582(.A1(new_n757), .A2(new_n765), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(new_n516), .A3(new_n476), .A4(new_n675), .ZN(new_n770));
  INV_X1    g584(.A(new_n710), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n770), .A2(new_n746), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n764), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n707), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n768), .A2(KEYINPUT51), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n742), .A2(new_n378), .ZN(new_n777));
  INV_X1    g591(.A(new_n759), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n742), .A2(new_n378), .A3(new_n759), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n779), .B(new_n780), .C1(new_n378), .C2(new_n687), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT116), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n764), .A2(new_n703), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n783), .A2(new_n757), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT114), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n781), .A2(KEYINPUT116), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n776), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n596), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n773), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(KEYINPUT48), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n612), .A2(new_n626), .A3(new_n688), .ZN(new_n792));
  INV_X1    g606(.A(new_n623), .ZN(new_n793));
  OAI221_X1 g607(.A(new_n473), .B1(new_n792), .B2(new_n783), .C1(new_n770), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n790), .A2(KEYINPUT48), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n791), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n768), .A2(new_n775), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n781), .A2(new_n785), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT115), .B1(new_n768), .B2(new_n775), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n788), .B(new_n796), .C1(new_n802), .C2(KEYINPUT51), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n652), .B(new_n653), .C1(new_n661), .C2(new_n679), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n805), .B1(new_n644), .B2(new_n655), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n645), .A2(KEYINPUT111), .A3(new_n656), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n379), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n652), .A2(new_n699), .A3(new_n674), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n804), .A2(new_n809), .A3(new_n714), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n804), .A2(new_n809), .A3(new_n714), .A4(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n684), .A2(new_n696), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n612), .A2(new_n626), .A3(new_n699), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n704), .A2(new_n516), .A3(new_n602), .A4(new_n702), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n816), .A2(new_n792), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n819), .A2(new_n690), .A3(new_n694), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n308), .A2(new_n310), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n634), .A2(KEYINPUT109), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT109), .B1(new_n634), .B2(new_n623), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n480), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n605), .A2(new_n607), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n483), .B1(new_n596), .B2(new_n646), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n725), .B1(new_n719), .B2(new_n722), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n645), .A2(new_n746), .A3(new_n470), .A4(new_n655), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n684), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n717), .A2(new_n600), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT110), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n720), .A2(new_n833), .A3(new_n684), .A4(new_n829), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n832), .A2(new_n834), .B1(new_n713), .B2(new_n720), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n820), .A2(new_n827), .A3(new_n828), .A4(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT53), .B1(new_n815), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT112), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n814), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n812), .A2(KEYINPUT112), .A3(new_n813), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n828), .A2(new_n835), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n697), .B(new_n705), .C1(new_n627), .C2(new_n689), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n825), .A2(new_n826), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n844), .A3(new_n694), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n837), .B(KEYINPUT54), .C1(new_n841), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n846), .B1(new_n815), .B2(new_n836), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n819), .A2(new_n690), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n689), .A2(new_n635), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT113), .B1(new_n843), .B2(new_n694), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n844), .A2(new_n846), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n842), .A2(new_n853), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n849), .B1(new_n841), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n848), .B1(new_n857), .B2(KEYINPUT54), .ZN(new_n858));
  OAI22_X1  g672(.A1(new_n803), .A2(new_n858), .B1(G952), .B2(G953), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n687), .A2(KEYINPUT49), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n516), .A2(new_n747), .A3(new_n309), .A4(new_n378), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n687), .A2(KEYINPUT49), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n670), .A2(new_n675), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n859), .A2(new_n864), .ZN(G75));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n857), .A2(new_n866), .A3(new_n477), .A4(new_n188), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT56), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n301), .A2(new_n302), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(new_n303), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n854), .A2(new_n853), .A3(new_n855), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(new_n842), .A3(new_n839), .A4(new_n840), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n369), .B1(new_n874), .B2(new_n849), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n866), .B1(new_n875), .B2(new_n188), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n312), .A2(G952), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT56), .B1(new_n875), .B2(new_n188), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n871), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n877), .A2(new_n881), .ZN(G51));
  NOR2_X1   g696(.A1(new_n857), .A2(KEYINPUT54), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n874), .B2(new_n849), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n371), .B(KEYINPUT57), .Z(new_n887));
  OAI21_X1  g701(.A(new_n367), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n875), .A2(new_n736), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(G54));
  AND2_X1   g704(.A1(KEYINPUT58), .A2(G475), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n857), .A2(new_n477), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n423), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n857), .A2(new_n477), .A3(new_n429), .A4(new_n891), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n879), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n893), .A2(KEYINPUT118), .A3(new_n879), .A4(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(G60));
  XOR2_X1   g713(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n900));
  NOR2_X1   g714(.A1(new_n468), .A2(new_n276), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n619), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n879), .B1(new_n886), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n619), .B1(new_n858), .B2(new_n903), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(G63));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT120), .Z(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT60), .Z(new_n910));
  NAND2_X1  g724(.A1(new_n857), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(new_n641), .ZN(new_n912));
  INV_X1    g726(.A(new_n506), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n878), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n912), .B(new_n914), .C1(new_n915), .C2(KEYINPUT61), .ZN(new_n916));
  INV_X1    g730(.A(new_n910), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n874), .B2(new_n849), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n915), .B(new_n879), .C1(new_n918), .C2(new_n506), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n879), .B1(new_n918), .B2(new_n506), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n911), .A2(new_n641), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n919), .B(new_n920), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n916), .A2(new_n923), .ZN(G66));
  OAI21_X1  g738(.A(G953), .B1(new_n479), .B2(new_n251), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT122), .Z(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n845), .B2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n869), .B1(G898), .B2(new_n312), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  XNOR2_X1  g743(.A(new_n552), .B(new_n399), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT124), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n804), .A2(new_n932), .A3(new_n714), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n932), .B1(new_n804), .B2(new_n714), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n828), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n758), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n779), .B2(new_n780), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n789), .A2(new_n817), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n745), .A2(new_n754), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n938), .A2(new_n312), .A3(new_n755), .A4(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n654), .B2(new_n312), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n822), .A2(new_n823), .ZN(new_n943));
  OR4_X1    g757(.A1(new_n789), .A2(new_n757), .A3(new_n667), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n755), .A2(new_n762), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n933), .A2(new_n934), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n676), .ZN(new_n948));
  INV_X1    g762(.A(new_n676), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(KEYINPUT62), .C1(new_n934), .C2(new_n933), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n951), .A2(G953), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n931), .B(new_n942), .C1(new_n952), .C2(KEYINPUT123), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n930), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n312), .B1(G227), .B2(G900), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n953), .A2(new_n957), .A3(new_n955), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G72));
  NAND2_X1  g775(.A1(new_n948), .A2(new_n950), .ZN(new_n962));
  INV_X1    g776(.A(new_n945), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(new_n845), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n967), .A2(KEYINPUT125), .A3(new_n542), .A4(new_n589), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n969));
  INV_X1    g783(.A(new_n966), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n951), .B2(new_n845), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n589), .A2(new_n542), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n938), .A2(new_n755), .A3(new_n845), .A4(new_n940), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n966), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n589), .A2(new_n542), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n975), .B(new_n879), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n976), .B2(new_n966), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT126), .B1(new_n981), .B2(new_n878), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n568), .A2(new_n572), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n970), .B1(new_n984), .B2(new_n590), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n837), .B(new_n985), .C1(new_n841), .C2(new_n847), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n974), .A2(new_n983), .A3(new_n986), .ZN(G57));
endmodule


