

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775;

  NOR2_X1 U379 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U380 ( .A1(n602), .A2(n775), .ZN(n401) );
  XOR2_X1 U381 ( .A(n606), .B(KEYINPUT79), .Z(n357) );
  XNOR2_X1 U382 ( .A(n465), .B(n464), .ZN(n546) );
  XNOR2_X2 U383 ( .A(n552), .B(KEYINPUT22), .ZN(n584) );
  XNOR2_X1 U384 ( .A(n399), .B(n523), .ZN(n545) );
  INV_X1 U385 ( .A(n702), .ZN(n615) );
  NOR2_X1 U386 ( .A1(n383), .A2(n673), .ZN(n576) );
  NOR2_X1 U387 ( .A1(n545), .A2(n607), .ZN(n448) );
  AND2_X1 U388 ( .A1(n616), .A2(n615), .ZN(n691) );
  AND2_X1 U389 ( .A1(n522), .A2(n521), .ZN(n621) );
  AND2_X1 U390 ( .A1(n569), .A2(n565), .ZN(n675) );
  AND2_X1 U391 ( .A1(n686), .A2(n611), .ZN(n624) );
  XNOR2_X1 U392 ( .A(n607), .B(KEYINPUT105), .ZN(n686) );
  NAND2_X1 U393 ( .A1(n544), .A2(n543), .ZN(n607) );
  NAND2_X1 U394 ( .A1(n546), .A2(n717), .ZN(n422) );
  XNOR2_X1 U395 ( .A(n390), .B(G113), .ZN(n392) );
  XNOR2_X1 U396 ( .A(n496), .B(G119), .ZN(n478) );
  INV_X2 U397 ( .A(G104), .ZN(n390) );
  NOR2_X1 U398 ( .A1(n647), .A2(n646), .ZN(n358) );
  INV_X1 U399 ( .A(n610), .ZN(n359) );
  NOR2_X2 U400 ( .A1(n694), .A2(n636), .ZN(n647) );
  XNOR2_X1 U401 ( .A(n558), .B(n554), .ZN(n608) );
  XNOR2_X2 U402 ( .A(n563), .B(n562), .ZN(n689) );
  NAND2_X1 U403 ( .A1(n643), .A2(n429), .ZN(n428) );
  NOR2_X1 U404 ( .A1(n431), .A2(n430), .ZN(n429) );
  XNOR2_X1 U405 ( .A(n401), .B(KEYINPUT46), .ZN(n400) );
  XNOR2_X1 U406 ( .A(n497), .B(n744), .ZN(n516) );
  INV_X1 U407 ( .A(n675), .ZN(n377) );
  NAND2_X1 U408 ( .A1(n716), .A2(KEYINPUT103), .ZN(n381) );
  AND2_X1 U409 ( .A1(n404), .A2(n427), .ZN(n426) );
  INV_X1 U410 ( .A(n630), .ZN(n427) );
  NAND2_X1 U411 ( .A1(n431), .A2(n430), .ZN(n404) );
  OR2_X1 U412 ( .A1(n774), .A2(n638), .ZN(n431) );
  NAND2_X1 U413 ( .A1(n380), .A2(n378), .ZN(n383) );
  NAND2_X1 U414 ( .A1(n400), .A2(n402), .ZN(n370) );
  OR2_X1 U415 ( .A1(n664), .A2(G902), .ZN(n517) );
  XNOR2_X1 U416 ( .A(n494), .B(G122), .ZN(n536) );
  XNOR2_X1 U417 ( .A(n407), .B(n405), .ZN(n535) );
  XNOR2_X1 U418 ( .A(n406), .B(G134), .ZN(n405) );
  XNOR2_X1 U419 ( .A(n449), .B(n408), .ZN(n407) );
  INV_X1 U420 ( .A(G116), .ZN(n406) );
  NAND2_X1 U421 ( .A1(n469), .A2(G234), .ZN(n471) );
  XNOR2_X1 U422 ( .A(n433), .B(n432), .ZN(n412) );
  INV_X1 U423 ( .A(KEYINPUT106), .ZN(n432) );
  NAND2_X1 U424 ( .A1(n624), .A2(n717), .ZN(n433) );
  NAND2_X1 U425 ( .A1(n621), .A2(n718), .ZN(n399) );
  XNOR2_X1 U426 ( .A(n416), .B(n415), .ZN(n568) );
  XNOR2_X1 U427 ( .A(G478), .B(KEYINPUT102), .ZN(n415) );
  OR2_X1 U428 ( .A1(n740), .A2(G902), .ZN(n416) );
  INV_X1 U429 ( .A(KEYINPUT71), .ZN(n430) );
  NAND2_X1 U430 ( .A1(n381), .A2(n363), .ZN(n374) );
  OR2_X1 U431 ( .A1(n675), .A2(n382), .ZN(n379) );
  AND2_X1 U432 ( .A1(n403), .A2(n620), .ZN(n402) );
  NOR2_X1 U433 ( .A1(n357), .A2(n773), .ZN(n403) );
  INV_X1 U434 ( .A(G237), .ZN(n462) );
  INV_X1 U435 ( .A(G119), .ZN(n508) );
  XNOR2_X1 U436 ( .A(G134), .B(G131), .ZN(n758) );
  XNOR2_X1 U437 ( .A(n537), .B(KEYINPUT4), .ZN(n760) );
  INV_X1 U438 ( .A(KEYINPUT44), .ZN(n585) );
  XNOR2_X1 U439 ( .A(n391), .B(G140), .ZN(n491) );
  INV_X1 U440 ( .A(G137), .ZN(n391) );
  XNOR2_X1 U441 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n408) );
  XNOR2_X1 U442 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n449) );
  NOR2_X1 U443 ( .A1(G953), .A2(G237), .ZN(n524) );
  XNOR2_X1 U444 ( .A(n491), .B(n390), .ZN(n492) );
  XOR2_X1 U445 ( .A(KEYINPUT74), .B(KEYINPUT90), .Z(n490) );
  XNOR2_X1 U446 ( .A(n760), .B(G101), .ZN(n497) );
  NOR2_X1 U447 ( .A1(n643), .A2(KEYINPUT71), .ZN(n445) );
  INV_X1 U448 ( .A(KEYINPUT81), .ZN(n447) );
  INV_X1 U449 ( .A(KEYINPUT18), .ZN(n453) );
  XNOR2_X1 U450 ( .A(n452), .B(n451), .ZN(n456) );
  XOR2_X1 U451 ( .A(KEYINPUT89), .B(KEYINPUT17), .Z(n452) );
  INV_X1 U452 ( .A(n431), .ZN(n629) );
  XNOR2_X1 U453 ( .A(KEYINPUT68), .B(KEYINPUT88), .ZN(n459) );
  INV_X1 U454 ( .A(KEYINPUT3), .ZN(n458) );
  XNOR2_X1 U455 ( .A(n425), .B(n423), .ZN(n746) );
  XNOR2_X1 U456 ( .A(n536), .B(n424), .ZN(n423) );
  XNOR2_X1 U457 ( .A(n392), .B(n478), .ZN(n425) );
  INV_X1 U458 ( .A(KEYINPUT16), .ZN(n424) );
  INV_X2 U459 ( .A(G953), .ZN(n469) );
  XNOR2_X1 U460 ( .A(G143), .B(G122), .ZN(n436) );
  XNOR2_X1 U461 ( .A(G140), .B(KEYINPUT11), .ZN(n528) );
  XOR2_X1 U462 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n529) );
  INV_X1 U463 ( .A(KEYINPUT10), .ZN(n467) );
  XNOR2_X1 U464 ( .A(n461), .B(n516), .ZN(n651) );
  XNOR2_X1 U465 ( .A(n746), .B(n457), .ZN(n461) );
  XNOR2_X1 U466 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U467 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n501) );
  INV_X1 U469 ( .A(KEYINPUT33), .ZN(n396) );
  OR2_X2 U470 ( .A1(n571), .A2(n702), .ZN(n397) );
  OR2_X1 U471 ( .A1(n702), .A2(n625), .ZN(n413) );
  INV_X1 U472 ( .A(KEYINPUT96), .ZN(n560) );
  NAND2_X1 U473 ( .A1(n621), .A2(n626), .ZN(n389) );
  INV_X1 U474 ( .A(KEYINPUT110), .ZN(n388) );
  INV_X1 U475 ( .A(KEYINPUT19), .ZN(n547) );
  XNOR2_X1 U476 ( .A(n597), .B(n596), .ZN(n600) );
  XNOR2_X1 U477 ( .A(n595), .B(KEYINPUT113), .ZN(n596) );
  XNOR2_X1 U478 ( .A(n558), .B(KEYINPUT104), .ZN(n591) );
  AND2_X1 U479 ( .A1(n589), .A2(n360), .ZN(n367) );
  XNOR2_X1 U480 ( .A(n539), .B(n538), .ZN(n740) );
  XNOR2_X1 U481 ( .A(n535), .B(n534), .ZN(n539) );
  XNOR2_X1 U482 ( .A(n437), .B(n434), .ZN(n659) );
  XNOR2_X1 U483 ( .A(n527), .B(n435), .ZN(n434) );
  XNOR2_X1 U484 ( .A(n530), .B(n438), .ZN(n437) );
  XNOR2_X1 U485 ( .A(n525), .B(n436), .ZN(n435) );
  BUF_X1 U486 ( .A(n669), .Z(n739) );
  XNOR2_X1 U487 ( .A(n655), .B(KEYINPUT87), .ZN(n743) );
  XNOR2_X1 U488 ( .A(n698), .B(KEYINPUT82), .ZN(n368) );
  XNOR2_X1 U489 ( .A(n448), .B(KEYINPUT40), .ZN(n602) );
  XNOR2_X1 U490 ( .A(n385), .B(KEYINPUT111), .ZN(n773) );
  NAND2_X1 U491 ( .A1(n387), .A2(n386), .ZN(n385) );
  INV_X1 U492 ( .A(n622), .ZN(n386) );
  XNOR2_X1 U493 ( .A(n389), .B(n388), .ZN(n387) );
  XOR2_X1 U494 ( .A(n488), .B(KEYINPUT21), .Z(n360) );
  INV_X1 U495 ( .A(n716), .ZN(n384) );
  XOR2_X1 U496 ( .A(n514), .B(G107), .Z(n361) );
  AND2_X1 U497 ( .A1(n413), .A2(n627), .ZN(n362) );
  NAND2_X1 U498 ( .A1(n384), .A2(n382), .ZN(n363) );
  NOR2_X1 U499 ( .A1(n712), .A2(n372), .ZN(n364) );
  INV_X1 U500 ( .A(G107), .ZN(n494) );
  INV_X1 U501 ( .A(G902), .ZN(n463) );
  XOR2_X1 U502 ( .A(KEYINPUT65), .B(KEYINPUT0), .Z(n365) );
  XNOR2_X1 U503 ( .A(KEYINPUT15), .B(G902), .ZN(n630) );
  XNOR2_X1 U504 ( .A(n623), .B(KEYINPUT48), .ZN(n366) );
  NAND2_X1 U505 ( .A1(n377), .A2(n381), .ZN(n376) );
  NAND2_X1 U506 ( .A1(n569), .A2(n367), .ZN(n552) );
  NAND2_X1 U507 ( .A1(n368), .A2(n700), .ZN(n731) );
  XNOR2_X1 U508 ( .A(n442), .B(n369), .ZN(n441) );
  XNOR2_X1 U509 ( .A(n481), .B(n480), .ZN(n369) );
  XNOR2_X2 U510 ( .A(n370), .B(n366), .ZN(n643) );
  XNOR2_X1 U511 ( .A(n371), .B(n668), .ZN(G57) );
  NOR2_X2 U512 ( .A1(n667), .A2(n743), .ZN(n371) );
  XNOR2_X1 U513 ( .A(n443), .B(n447), .ZN(n633) );
  NAND2_X1 U514 ( .A1(n428), .A2(n426), .ZN(n446) );
  AND2_X2 U515 ( .A1(n372), .A2(n569), .ZN(n562) );
  XNOR2_X1 U516 ( .A(n561), .B(n560), .ZN(n372) );
  NOR2_X1 U517 ( .A1(n733), .A2(G902), .ZN(n500) );
  XNOR2_X1 U518 ( .A(n498), .B(n373), .ZN(n733) );
  XNOR2_X1 U519 ( .A(n495), .B(n361), .ZN(n373) );
  NAND2_X1 U520 ( .A1(n375), .A2(n374), .ZN(n380) );
  OR2_X2 U521 ( .A1(n689), .A2(n376), .ZN(n375) );
  OR2_X1 U522 ( .A1(n689), .A2(n379), .ZN(n378) );
  INV_X1 U523 ( .A(KEYINPUT103), .ZN(n382) );
  XNOR2_X1 U524 ( .A(n526), .B(n392), .ZN(n438) );
  XNOR2_X2 U525 ( .A(n393), .B(n365), .ZN(n569) );
  NOR2_X2 U526 ( .A1(n604), .A2(n551), .ZN(n393) );
  XNOR2_X2 U527 ( .A(n613), .B(n547), .ZN(n604) );
  XNOR2_X2 U528 ( .A(n422), .B(KEYINPUT86), .ZN(n613) );
  XNOR2_X2 U529 ( .A(G143), .B(G128), .ZN(n537) );
  XNOR2_X1 U530 ( .A(n394), .B(KEYINPUT34), .ZN(n572) );
  NAND2_X1 U531 ( .A1(n395), .A2(n569), .ZN(n394) );
  INV_X1 U532 ( .A(n724), .ZN(n395) );
  XNOR2_X2 U533 ( .A(n397), .B(n396), .ZN(n724) );
  NAND2_X1 U534 ( .A1(n706), .A2(n360), .ZN(n440) );
  XNOR2_X2 U535 ( .A(n398), .B(n486), .ZN(n706) );
  NAND2_X1 U536 ( .A1(n441), .A2(n463), .ZN(n398) );
  NAND2_X1 U537 ( .A1(n412), .A2(n414), .ZN(n410) );
  NOR2_X1 U538 ( .A1(n411), .A2(n409), .ZN(n628) );
  NAND2_X1 U539 ( .A1(n410), .A2(n362), .ZN(n409) );
  NOR2_X1 U540 ( .A1(n412), .A2(n625), .ZN(n411) );
  AND2_X1 U541 ( .A1(n702), .A2(n625), .ZN(n414) );
  XNOR2_X2 U542 ( .A(n417), .B(KEYINPUT45), .ZN(n753) );
  NAND2_X1 U543 ( .A1(n419), .A2(n418), .ZN(n417) );
  XNOR2_X1 U544 ( .A(n421), .B(KEYINPUT85), .ZN(n418) );
  NAND2_X1 U545 ( .A1(n420), .A2(n588), .ZN(n419) );
  XNOR2_X1 U546 ( .A(n587), .B(n585), .ZN(n420) );
  NAND2_X1 U547 ( .A1(n576), .A2(n575), .ZN(n421) );
  NOR2_X1 U548 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X2 U549 ( .A1(n656), .A2(n743), .ZN(n658) );
  NOR2_X2 U550 ( .A1(n662), .A2(n743), .ZN(n663) );
  NOR2_X2 U551 ( .A1(n572), .A2(n622), .ZN(n574) );
  NOR2_X1 U552 ( .A1(n446), .A2(n445), .ZN(n444) );
  XNOR2_X1 U553 ( .A(n439), .B(KEYINPUT72), .ZN(n522) );
  NOR2_X2 U554 ( .A1(n701), .A2(n507), .ZN(n439) );
  XNOR2_X2 U555 ( .A(n440), .B(KEYINPUT66), .ZN(n701) );
  XNOR2_X1 U556 ( .A(n441), .B(KEYINPUT123), .ZN(n670) );
  INV_X1 U557 ( .A(n762), .ZN(n442) );
  NAND2_X1 U558 ( .A1(n444), .A2(n753), .ZN(n443) );
  NAND2_X1 U559 ( .A1(n643), .A2(n629), .ZN(n763) );
  NOR2_X1 U560 ( .A1(n699), .A2(G953), .ZN(n700) );
  NAND2_X1 U561 ( .A1(n619), .A2(n618), .ZN(n450) );
  NOR2_X1 U562 ( .A1(n691), .A2(n450), .ZN(n620) );
  XNOR2_X1 U563 ( .A(n493), .B(n492), .ZN(n495) );
  INV_X1 U564 ( .A(KEYINPUT28), .ZN(n595) );
  INV_X1 U565 ( .A(KEYINPUT6), .ZN(n554) );
  XNOR2_X1 U566 ( .A(KEYINPUT35), .B(KEYINPUT75), .ZN(n573) );
  XOR2_X1 U567 ( .A(G134), .B(KEYINPUT117), .Z(n541) );
  XNOR2_X1 U568 ( .A(G146), .B(G125), .ZN(n468) );
  INV_X1 U569 ( .A(n468), .ZN(n451) );
  NAND2_X1 U570 ( .A1(G224), .A2(n469), .ZN(n454) );
  XNOR2_X1 U571 ( .A(n458), .B(G116), .ZN(n460) );
  XNOR2_X1 U572 ( .A(n460), .B(n459), .ZN(n744) );
  NAND2_X1 U573 ( .A1(n651), .A2(n630), .ZN(n465) );
  NAND2_X1 U574 ( .A1(n463), .A2(n462), .ZN(n518) );
  AND2_X1 U575 ( .A1(n518), .A2(G210), .ZN(n464) );
  BUF_X1 U576 ( .A(n546), .Z(n626) );
  INV_X1 U577 ( .A(KEYINPUT38), .ZN(n466) );
  XNOR2_X1 U578 ( .A(n626), .B(n466), .ZN(n718) );
  XNOR2_X1 U579 ( .A(n468), .B(n467), .ZN(n527) );
  XNOR2_X1 U580 ( .A(n527), .B(n491), .ZN(n762) );
  INV_X1 U581 ( .A(KEYINPUT8), .ZN(n470) );
  XNOR2_X2 U582 ( .A(n471), .B(n470), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n533), .A2(G221), .ZN(n475) );
  XNOR2_X1 U584 ( .A(KEYINPUT93), .B(KEYINPUT24), .ZN(n473) );
  XNOR2_X1 U585 ( .A(KEYINPUT73), .B(KEYINPUT80), .ZN(n472) );
  XNOR2_X1 U586 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U587 ( .A(n475), .B(n474), .ZN(n481) );
  XNOR2_X1 U588 ( .A(G128), .B(KEYINPUT92), .ZN(n477) );
  XNOR2_X1 U589 ( .A(KEYINPUT23), .B(KEYINPUT91), .ZN(n476) );
  XNOR2_X1 U590 ( .A(n477), .B(n476), .ZN(n479) );
  XNOR2_X1 U591 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U592 ( .A1(n630), .A2(G234), .ZN(n483) );
  XNOR2_X1 U593 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n482) );
  XNOR2_X1 U594 ( .A(n483), .B(n482), .ZN(n487) );
  NAND2_X1 U595 ( .A1(n487), .A2(G217), .ZN(n485) );
  XNOR2_X1 U596 ( .A(KEYINPUT95), .B(KEYINPUT25), .ZN(n484) );
  XNOR2_X1 U597 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U598 ( .A1(n487), .A2(G221), .ZN(n488) );
  NAND2_X1 U599 ( .A1(G227), .A2(n469), .ZN(n489) );
  XNOR2_X1 U600 ( .A(n490), .B(n489), .ZN(n493) );
  XNOR2_X1 U601 ( .A(n758), .B(G146), .ZN(n514) );
  INV_X2 U602 ( .A(G110), .ZN(n496) );
  XNOR2_X1 U603 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U604 ( .A(KEYINPUT67), .B(G469), .ZN(n499) );
  XNOR2_X2 U605 ( .A(n500), .B(n499), .ZN(n598) );
  XOR2_X1 U606 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n502) );
  XOR2_X1 U607 ( .A(n502), .B(n501), .Z(n503) );
  NAND2_X1 U608 ( .A1(G952), .A2(n503), .ZN(n729) );
  NOR2_X1 U609 ( .A1(n729), .A2(G953), .ZN(n550) );
  INV_X1 U610 ( .A(n550), .ZN(n506) );
  AND2_X1 U611 ( .A1(n503), .A2(G953), .ZN(n504) );
  NAND2_X1 U612 ( .A1(G902), .A2(n504), .ZN(n548) );
  OR2_X1 U613 ( .A1(n548), .A2(G900), .ZN(n505) );
  NAND2_X1 U614 ( .A1(n506), .A2(n505), .ZN(n592) );
  NAND2_X1 U615 ( .A1(n598), .A2(n592), .ZN(n507) );
  NAND2_X1 U616 ( .A1(n524), .A2(G210), .ZN(n510) );
  XNOR2_X1 U617 ( .A(n508), .B(G137), .ZN(n509) );
  XNOR2_X1 U618 ( .A(n510), .B(n509), .ZN(n512) );
  XNOR2_X1 U619 ( .A(G113), .B(KEYINPUT5), .ZN(n511) );
  XNOR2_X1 U620 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U621 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n516), .B(n515), .ZN(n664) );
  XNOR2_X2 U623 ( .A(n517), .B(G472), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n518), .A2(G214), .ZN(n717) );
  NAND2_X1 U625 ( .A1(n591), .A2(n717), .ZN(n520) );
  XNOR2_X1 U626 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n519) );
  XNOR2_X1 U627 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U628 ( .A(KEYINPUT69), .B(KEYINPUT39), .ZN(n523) );
  INV_X1 U629 ( .A(n545), .ZN(n540) );
  XNOR2_X1 U630 ( .A(KEYINPUT13), .B(G475), .ZN(n532) );
  XOR2_X1 U631 ( .A(G131), .B(KEYINPUT98), .Z(n526) );
  NAND2_X1 U632 ( .A1(G214), .A2(n524), .ZN(n525) );
  XNOR2_X1 U633 ( .A(n529), .B(n528), .ZN(n530) );
  NOR2_X1 U634 ( .A1(G902), .A2(n659), .ZN(n531) );
  XNOR2_X1 U635 ( .A(n532), .B(n531), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n567), .B(KEYINPUT99), .ZN(n542) );
  NAND2_X1 U637 ( .A1(G217), .A2(n533), .ZN(n534) );
  XOR2_X1 U638 ( .A(n537), .B(n536), .Z(n538) );
  AND2_X1 U639 ( .A1(n542), .A2(n568), .ZN(n688) );
  AND2_X1 U640 ( .A1(n540), .A2(n688), .ZN(n638) );
  XOR2_X1 U641 ( .A(n541), .B(n638), .Z(G36) );
  INV_X1 U642 ( .A(n568), .ZN(n544) );
  INV_X1 U643 ( .A(n542), .ZN(n543) );
  XOR2_X1 U644 ( .A(n602), .B(G131), .Z(G33) );
  NOR2_X1 U645 ( .A1(n548), .A2(G898), .ZN(n549) );
  NOR2_X1 U646 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U647 ( .A1(n567), .A2(n568), .ZN(n589) );
  INV_X1 U648 ( .A(KEYINPUT1), .ZN(n553) );
  XNOR2_X2 U649 ( .A(n598), .B(n553), .ZN(n702) );
  INV_X1 U650 ( .A(n706), .ZN(n555) );
  NOR2_X1 U651 ( .A1(n359), .A2(n555), .ZN(n556) );
  NAND2_X1 U652 ( .A1(n702), .A2(n556), .ZN(n557) );
  NOR2_X1 U653 ( .A1(n584), .A2(n557), .ZN(n673) );
  INV_X1 U654 ( .A(KEYINPUT31), .ZN(n563) );
  INV_X1 U655 ( .A(n558), .ZN(n708) );
  NOR2_X1 U656 ( .A1(n701), .A2(n708), .ZN(n559) );
  NAND2_X1 U657 ( .A1(n615), .A2(n559), .ZN(n561) );
  NAND2_X1 U658 ( .A1(n598), .A2(n708), .ZN(n564) );
  NOR2_X1 U659 ( .A1(n701), .A2(n564), .ZN(n565) );
  INV_X1 U660 ( .A(n688), .ZN(n566) );
  AND2_X1 U661 ( .A1(n566), .A2(n607), .ZN(n716) );
  NAND2_X1 U662 ( .A1(n568), .A2(n567), .ZN(n622) );
  INV_X1 U663 ( .A(n701), .ZN(n570) );
  NAND2_X1 U664 ( .A1(n570), .A2(n608), .ZN(n571) );
  XNOR2_X2 U665 ( .A(n574), .B(n573), .ZN(n586) );
  NAND2_X1 U666 ( .A1(KEYINPUT44), .A2(n586), .ZN(n575) );
  XNOR2_X1 U667 ( .A(n608), .B(KEYINPUT76), .ZN(n577) );
  OR2_X1 U668 ( .A1(n577), .A2(n706), .ZN(n578) );
  OR2_X1 U669 ( .A1(n702), .A2(n578), .ZN(n579) );
  NOR2_X1 U670 ( .A1(n584), .A2(n579), .ZN(n581) );
  XNOR2_X1 U671 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n580) );
  XNOR2_X1 U672 ( .A(n581), .B(n580), .ZN(n772) );
  NOR2_X1 U673 ( .A1(n591), .A2(n706), .ZN(n582) );
  NAND2_X1 U674 ( .A1(n702), .A2(n582), .ZN(n583) );
  NOR2_X1 U675 ( .A1(n584), .A2(n583), .ZN(n679) );
  NOR2_X2 U676 ( .A1(n772), .A2(n679), .ZN(n587) );
  NAND2_X1 U677 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U678 ( .A1(n718), .A2(n717), .ZN(n715) );
  INV_X1 U679 ( .A(n589), .ZN(n720) );
  NOR2_X1 U680 ( .A1(n715), .A2(n720), .ZN(n590) );
  XNOR2_X1 U681 ( .A(n590), .B(KEYINPUT41), .ZN(n714) );
  INV_X1 U682 ( .A(n591), .ZN(n594) );
  NAND2_X1 U683 ( .A1(n360), .A2(n592), .ZN(n593) );
  OR2_X1 U684 ( .A1(n706), .A2(n593), .ZN(n609) );
  NOR2_X1 U685 ( .A1(n594), .A2(n609), .ZN(n597) );
  XNOR2_X1 U686 ( .A(n598), .B(KEYINPUT112), .ZN(n599) );
  NAND2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n603) );
  NOR2_X1 U688 ( .A1(n714), .A2(n603), .ZN(n601) );
  XNOR2_X1 U689 ( .A(n601), .B(KEYINPUT42), .ZN(n775) );
  NOR2_X2 U690 ( .A1(n604), .A2(n603), .ZN(n683) );
  INV_X1 U691 ( .A(KEYINPUT47), .ZN(n605) );
  NOR2_X1 U692 ( .A1(n683), .A2(n605), .ZN(n606) );
  INV_X1 U693 ( .A(n608), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U695 ( .A(KEYINPUT114), .B(n624), .Z(n612) );
  NOR2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U697 ( .A(n614), .B(KEYINPUT36), .ZN(n616) );
  NOR2_X1 U698 ( .A1(n716), .A2(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n683), .A2(n617), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n716), .A2(KEYINPUT47), .ZN(n618) );
  INV_X1 U701 ( .A(KEYINPUT84), .ZN(n623) );
  XOR2_X1 U702 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n625) );
  INV_X1 U703 ( .A(n626), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n628), .B(KEYINPUT108), .ZN(n774) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT83), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n631), .A2(KEYINPUT2), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n648) );
  INV_X1 U708 ( .A(n763), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n753), .A2(n634), .ZN(n694) );
  INV_X1 U710 ( .A(KEYINPUT77), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n635), .A2(KEYINPUT2), .ZN(n636) );
  INV_X1 U712 ( .A(n774), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n637), .A2(KEYINPUT77), .ZN(n641) );
  INV_X1 U714 ( .A(n638), .ZN(n639) );
  AND2_X1 U715 ( .A1(n639), .A2(KEYINPUT2), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n753), .A2(n642), .ZN(n645) );
  INV_X1 U718 ( .A(n643), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n697) );
  AND2_X2 U720 ( .A1(n648), .A2(n697), .ZN(n669) );
  NAND2_X1 U721 ( .A1(n669), .A2(G210), .ZN(n653) );
  XNOR2_X1 U722 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n649) );
  XNOR2_X1 U723 ( .A(n649), .B(KEYINPUT55), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n656) );
  INV_X1 U726 ( .A(G952), .ZN(n654) );
  NAND2_X1 U727 ( .A1(n654), .A2(G953), .ZN(n655) );
  XOR2_X1 U728 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n657) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(G51) );
  NAND2_X1 U730 ( .A1(n669), .A2(G475), .ZN(n661) );
  XOR2_X1 U731 ( .A(KEYINPUT59), .B(n659), .Z(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U734 ( .A(KEYINPUT63), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(G472), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n664), .B(KEYINPUT62), .ZN(n665) );
  XNOR2_X1 U737 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n739), .A2(G217), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U740 ( .A1(n672), .A2(n743), .ZN(G66) );
  XOR2_X1 U741 ( .A(G101), .B(n673), .Z(G3) );
  NAND2_X1 U742 ( .A1(n675), .A2(n686), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n674), .B(G104), .ZN(G6) );
  XOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n677) );
  NAND2_X1 U745 ( .A1(n675), .A2(n688), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U747 ( .A(G107), .B(n678), .ZN(G9) );
  XOR2_X1 U748 ( .A(G110), .B(n679), .Z(G12) );
  XOR2_X1 U749 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n681) );
  NAND2_X1 U750 ( .A1(n683), .A2(n688), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U752 ( .A(G128), .B(n682), .Z(G30) );
  NAND2_X1 U753 ( .A1(n683), .A2(n686), .ZN(n684) );
  XNOR2_X1 U754 ( .A(n684), .B(KEYINPUT116), .ZN(n685) );
  XNOR2_X1 U755 ( .A(G146), .B(n685), .ZN(G48) );
  NAND2_X1 U756 ( .A1(n686), .A2(n689), .ZN(n687) );
  XNOR2_X1 U757 ( .A(n687), .B(G113), .ZN(G15) );
  NAND2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U759 ( .A(n690), .B(G116), .ZN(G18) );
  XNOR2_X1 U760 ( .A(G125), .B(n691), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U762 ( .A(KEYINPUT2), .ZN(n693) );
  NAND2_X1 U763 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U764 ( .A(n695), .B(KEYINPUT78), .ZN(n696) );
  NAND2_X1 U765 ( .A1(n358), .A2(n696), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n724), .A2(n714), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n705) );
  XNOR2_X1 U768 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n703) );
  XNOR2_X1 U769 ( .A(n703), .B(KEYINPUT118), .ZN(n704) );
  XNOR2_X1 U770 ( .A(n705), .B(n704), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n706), .A2(n360), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT49), .ZN(n709) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U775 ( .A(KEYINPUT51), .B(n364), .Z(n713) );
  NOR2_X1 U776 ( .A1(n714), .A2(n713), .ZN(n726) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U781 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U783 ( .A(n727), .B(KEYINPUT52), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U785 ( .A(n732), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U786 ( .A1(n739), .A2(G469), .ZN(n737) );
  XOR2_X1 U787 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n735) );
  XNOR2_X1 U788 ( .A(n733), .B(KEYINPUT122), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(n736) );
  XNOR2_X1 U790 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U791 ( .A1(n743), .A2(n738), .ZN(G54) );
  NAND2_X1 U792 ( .A1(n739), .A2(G478), .ZN(n741) );
  XNOR2_X1 U793 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(G63) );
  XOR2_X1 U795 ( .A(G101), .B(n744), .Z(n745) );
  XNOR2_X1 U796 ( .A(n746), .B(n745), .ZN(n748) );
  NOR2_X1 U797 ( .A1(G898), .A2(n469), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U799 ( .A(KEYINPUT125), .B(n749), .Z(n757) );
  NAND2_X1 U800 ( .A1(G953), .A2(G224), .ZN(n750) );
  XNOR2_X1 U801 ( .A(KEYINPUT61), .B(n750), .ZN(n751) );
  NAND2_X1 U802 ( .A1(n751), .A2(G898), .ZN(n752) );
  XNOR2_X1 U803 ( .A(n752), .B(KEYINPUT124), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n753), .A2(n469), .ZN(n754) );
  NAND2_X1 U805 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(G69) );
  XOR2_X1 U807 ( .A(n758), .B(KEYINPUT90), .Z(n759) );
  XOR2_X1 U808 ( .A(n760), .B(n759), .Z(n761) );
  XNOR2_X1 U809 ( .A(n762), .B(n761), .ZN(n765) );
  XNOR2_X1 U810 ( .A(n763), .B(n765), .ZN(n764) );
  NOR2_X1 U811 ( .A1(n764), .A2(G953), .ZN(n770) );
  XOR2_X1 U812 ( .A(G227), .B(n765), .Z(n766) );
  NAND2_X1 U813 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U814 ( .A1(G953), .A2(n767), .ZN(n768) );
  XOR2_X1 U815 ( .A(KEYINPUT126), .B(n768), .Z(n769) );
  NOR2_X1 U816 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U817 ( .A(KEYINPUT127), .B(n771), .ZN(G72) );
  XOR2_X1 U818 ( .A(n772), .B(G119), .Z(G21) );
  XOR2_X1 U819 ( .A(G122), .B(n586), .Z(G24) );
  XOR2_X1 U820 ( .A(G143), .B(n773), .Z(G45) );
  XOR2_X1 U821 ( .A(G140), .B(n774), .Z(G42) );
  XOR2_X1 U822 ( .A(G137), .B(n775), .Z(G39) );
endmodule

