

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U560 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U561 ( .A1(G1384), .A2(G164), .ZN(n722) );
  NOR2_X1 U562 ( .A1(n540), .A2(n539), .ZN(G160) );
  BUF_X2 U563 ( .A(n898), .Z(n527) );
  XOR2_X1 U564 ( .A(KEYINPUT17), .B(n535), .Z(n898) );
  AND2_X1 U565 ( .A1(n700), .A2(n688), .ZN(n691) );
  INV_X4 U566 ( .A(n669), .ZN(n607) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n801) );
  AND2_X1 U568 ( .A1(n646), .A2(n645), .ZN(n528) );
  AND2_X1 U569 ( .A1(G8), .A2(n656), .ZN(n529) );
  NOR2_X1 U570 ( .A1(n666), .A2(n665), .ZN(n530) );
  XNOR2_X1 U571 ( .A(n608), .B(KEYINPUT27), .ZN(n609) );
  XNOR2_X1 U572 ( .A(n610), .B(n609), .ZN(n612) );
  NAND2_X1 U573 ( .A1(G8), .A2(n669), .ZN(n705) );
  AND2_X1 U574 ( .A1(n536), .A2(G2104), .ZN(n899) );
  XNOR2_X1 U575 ( .A(n624), .B(KEYINPUT15), .ZN(n988) );
  INV_X1 U576 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U577 ( .A1(G101), .A2(n899), .ZN(n531) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n531), .Z(n534) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n902) );
  NAND2_X1 U580 ( .A1(G113), .A2(n902), .ZN(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT65), .B(n532), .Z(n533) );
  NAND2_X1 U582 ( .A1(n534), .A2(n533), .ZN(n540) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  NAND2_X1 U584 ( .A1(G137), .A2(n527), .ZN(n538) );
  NOR2_X2 U585 ( .A1(G2104), .A2(n536), .ZN(n903) );
  NAND2_X1 U586 ( .A1(G125), .A2(n903), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U588 ( .A1(G138), .A2(n527), .ZN(n546) );
  AND2_X1 U589 ( .A1(G102), .A2(n899), .ZN(n544) );
  NAND2_X1 U590 ( .A1(G114), .A2(n902), .ZN(n542) );
  NAND2_X1 U591 ( .A1(G126), .A2(n903), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U593 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n546), .A2(n545), .ZN(n548) );
  INV_X1 U595 ( .A(KEYINPUT90), .ZN(n547) );
  XNOR2_X1 U596 ( .A(n548), .B(n547), .ZN(G164) );
  INV_X1 U597 ( .A(G651), .ZN(n554) );
  NOR2_X1 U598 ( .A1(G543), .A2(n554), .ZN(n549) );
  XOR2_X1 U599 ( .A(KEYINPUT66), .B(n549), .Z(n550) );
  XNOR2_X1 U600 ( .A(KEYINPUT1), .B(n550), .ZN(n802) );
  NAND2_X1 U601 ( .A1(G61), .A2(n802), .ZN(n553) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n586) );
  NOR2_X1 U603 ( .A1(G651), .A2(n586), .ZN(n551) );
  XNOR2_X1 U604 ( .A(KEYINPUT64), .B(n551), .ZN(n798) );
  NAND2_X1 U605 ( .A1(G48), .A2(n798), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n557) );
  NOR2_X2 U607 ( .A1(n586), .A2(n554), .ZN(n796) );
  NAND2_X1 U608 ( .A1(n796), .A2(G73), .ZN(n555) );
  XOR2_X1 U609 ( .A(KEYINPUT2), .B(n555), .Z(n556) );
  NOR2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n801), .A2(G86), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n559), .A2(n558), .ZN(G305) );
  NAND2_X1 U613 ( .A1(G64), .A2(n802), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G52), .A2(n798), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n567) );
  NAND2_X1 U616 ( .A1(n801), .A2(G90), .ZN(n562) );
  XOR2_X1 U617 ( .A(KEYINPUT69), .B(n562), .Z(n564) );
  NAND2_X1 U618 ( .A1(n796), .A2(G77), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U621 ( .A1(n567), .A2(n566), .ZN(G171) );
  INV_X1 U622 ( .A(G171), .ZN(G301) );
  NAND2_X1 U623 ( .A1(n801), .A2(G89), .ZN(n568) );
  XNOR2_X1 U624 ( .A(n568), .B(KEYINPUT4), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G76), .A2(n796), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U627 ( .A(n571), .B(KEYINPUT5), .ZN(n577) );
  XNOR2_X1 U628 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n575) );
  NAND2_X1 U629 ( .A1(G63), .A2(n802), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G51), .A2(n798), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U632 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U633 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U634 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  NAND2_X1 U635 ( .A1(G88), .A2(n801), .ZN(n580) );
  NAND2_X1 U636 ( .A1(G75), .A2(n796), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n580), .A2(n579), .ZN(n585) );
  NAND2_X1 U638 ( .A1(G62), .A2(n802), .ZN(n582) );
  NAND2_X1 U639 ( .A1(G50), .A2(n798), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U641 ( .A(KEYINPUT83), .B(n583), .Z(n584) );
  NOR2_X1 U642 ( .A1(n585), .A2(n584), .ZN(G166) );
  INV_X1 U643 ( .A(G166), .ZN(G303) );
  XOR2_X1 U644 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U645 ( .A1(G87), .A2(n586), .ZN(n588) );
  NAND2_X1 U646 ( .A1(G74), .A2(G651), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U648 ( .A1(n802), .A2(n589), .ZN(n591) );
  NAND2_X1 U649 ( .A1(G49), .A2(n798), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n591), .A2(n590), .ZN(G288) );
  NAND2_X1 U651 ( .A1(G60), .A2(n802), .ZN(n598) );
  NAND2_X1 U652 ( .A1(G85), .A2(n801), .ZN(n593) );
  NAND2_X1 U653 ( .A1(G72), .A2(n796), .ZN(n592) );
  NAND2_X1 U654 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U655 ( .A1(G47), .A2(n798), .ZN(n594) );
  XNOR2_X1 U656 ( .A(KEYINPUT67), .B(n594), .ZN(n595) );
  NOR2_X1 U657 ( .A1(n596), .A2(n595), .ZN(n597) );
  NAND2_X1 U658 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U659 ( .A(n599), .B(KEYINPUT68), .ZN(G290) );
  XNOR2_X1 U660 ( .A(G1981), .B(G305), .ZN(n985) );
  NAND2_X1 U661 ( .A1(G65), .A2(n802), .ZN(n601) );
  NAND2_X1 U662 ( .A1(G53), .A2(n798), .ZN(n600) );
  NAND2_X1 U663 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U664 ( .A1(G91), .A2(n801), .ZN(n603) );
  NAND2_X1 U665 ( .A1(G78), .A2(n796), .ZN(n602) );
  NAND2_X1 U666 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U667 ( .A1(n605), .A2(n604), .ZN(n989) );
  NAND2_X1 U668 ( .A1(G160), .A2(G40), .ZN(n721) );
  INV_X1 U669 ( .A(n721), .ZN(n606) );
  NAND2_X2 U670 ( .A1(n722), .A2(n606), .ZN(n669) );
  NAND2_X1 U671 ( .A1(G2072), .A2(n607), .ZN(n610) );
  INV_X1 U672 ( .A(KEYINPUT99), .ZN(n608) );
  INV_X1 U673 ( .A(G1956), .ZN(n1010) );
  NOR2_X1 U674 ( .A1(n607), .A2(n1010), .ZN(n611) );
  NOR2_X1 U675 ( .A1(n612), .A2(n611), .ZN(n644) );
  NOR2_X1 U676 ( .A1(n989), .A2(n644), .ZN(n614) );
  INV_X1 U677 ( .A(KEYINPUT28), .ZN(n613) );
  XNOR2_X1 U678 ( .A(n614), .B(n613), .ZN(n649) );
  NOR2_X1 U679 ( .A1(n607), .A2(G1348), .ZN(n616) );
  NOR2_X1 U680 ( .A1(G2067), .A2(n669), .ZN(n615) );
  NOR2_X1 U681 ( .A1(n616), .A2(n615), .ZN(n625) );
  NAND2_X1 U682 ( .A1(n798), .A2(G54), .ZN(n623) );
  NAND2_X1 U683 ( .A1(G92), .A2(n801), .ZN(n618) );
  NAND2_X1 U684 ( .A1(G66), .A2(n802), .ZN(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G79), .A2(n796), .ZN(n619) );
  XNOR2_X1 U687 ( .A(KEYINPUT75), .B(n619), .ZN(n620) );
  NOR2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n624) );
  INV_X1 U690 ( .A(n988), .ZN(n770) );
  OR2_X1 U691 ( .A1(n625), .A2(n770), .ZN(n647) );
  NAND2_X1 U692 ( .A1(n770), .A2(n625), .ZN(n643) );
  NAND2_X1 U693 ( .A1(G81), .A2(n801), .ZN(n626) );
  XOR2_X1 U694 ( .A(KEYINPUT12), .B(n626), .Z(n627) );
  XNOR2_X1 U695 ( .A(n627), .B(KEYINPUT73), .ZN(n629) );
  NAND2_X1 U696 ( .A1(G68), .A2(n796), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U698 ( .A(KEYINPUT13), .B(n630), .ZN(n636) );
  NAND2_X1 U699 ( .A1(n802), .A2(G56), .ZN(n631) );
  XOR2_X1 U700 ( .A(KEYINPUT14), .B(n631), .Z(n634) );
  NAND2_X1 U701 ( .A1(n798), .A2(G43), .ZN(n632) );
  XOR2_X1 U702 ( .A(KEYINPUT74), .B(n632), .Z(n633) );
  NOR2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n987) );
  XNOR2_X1 U705 ( .A(G1996), .B(KEYINPUT100), .ZN(n965) );
  NAND2_X1 U706 ( .A1(n607), .A2(n965), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT26), .ZN(n640) );
  NAND2_X1 U708 ( .A1(n669), .A2(G1341), .ZN(n638) );
  XOR2_X1 U709 ( .A(KEYINPUT101), .B(n638), .Z(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U711 ( .A1(n987), .A2(n641), .ZN(n642) );
  NAND2_X1 U712 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U713 ( .A1(n989), .A2(n644), .ZN(n645) );
  NAND2_X1 U714 ( .A1(n647), .A2(n528), .ZN(n648) );
  NAND2_X1 U715 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U716 ( .A(KEYINPUT102), .B(KEYINPUT29), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n655) );
  XOR2_X1 U718 ( .A(KEYINPUT25), .B(G2078), .Z(n966) );
  NOR2_X1 U719 ( .A1(n966), .A2(n669), .ZN(n653) );
  NOR2_X1 U720 ( .A1(n607), .A2(G1961), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n660) );
  NOR2_X1 U722 ( .A1(n660), .A2(G301), .ZN(n654) );
  NOR2_X2 U723 ( .A1(n655), .A2(n654), .ZN(n678) );
  NOR2_X1 U724 ( .A1(G1966), .A2(n705), .ZN(n666) );
  INV_X1 U725 ( .A(n666), .ZN(n657) );
  NOR2_X1 U726 ( .A1(G2084), .A2(n669), .ZN(n664) );
  INV_X1 U727 ( .A(n664), .ZN(n656) );
  NAND2_X1 U728 ( .A1(n657), .A2(n529), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT30), .B(n658), .ZN(n659) );
  NOR2_X1 U730 ( .A1(n659), .A2(G168), .ZN(n662) );
  AND2_X1 U731 ( .A1(G301), .A2(n660), .ZN(n661) );
  NOR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT31), .ZN(n676) );
  OR2_X1 U734 ( .A1(n678), .A2(n676), .ZN(n667) );
  AND2_X1 U735 ( .A1(G8), .A2(n664), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n667), .A2(n530), .ZN(n668) );
  XNOR2_X1 U737 ( .A(KEYINPUT103), .B(n668), .ZN(n685) );
  INV_X1 U738 ( .A(G8), .ZN(n675) );
  NOR2_X1 U739 ( .A1(G1971), .A2(n705), .ZN(n671) );
  NOR2_X1 U740 ( .A1(G2090), .A2(n669), .ZN(n670) );
  NOR2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(KEYINPUT104), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n673), .A2(G303), .ZN(n674) );
  NOR2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n680) );
  OR2_X1 U745 ( .A1(n676), .A2(n680), .ZN(n677) );
  AND2_X1 U746 ( .A1(G286), .A2(G8), .ZN(n679) );
  OR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U749 ( .A(n683), .B(KEYINPUT32), .Z(n684) );
  NOR2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U751 ( .A(n686), .B(KEYINPUT105), .ZN(n700) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n993), .A2(n687), .ZN(n688) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n994) );
  INV_X1 U756 ( .A(n705), .ZN(n689) );
  NAND2_X1 U757 ( .A1(n994), .A2(n689), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U759 ( .A1(n692), .A2(KEYINPUT33), .ZN(n693) );
  XNOR2_X1 U760 ( .A(n693), .B(KEYINPUT106), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n985), .A2(n694), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n993), .A2(KEYINPUT33), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n705), .A2(n695), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n696), .B(KEYINPUT107), .ZN(n697) );
  AND2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n709) );
  NOR2_X1 U766 ( .A1(G2090), .A2(G303), .ZN(n699) );
  NAND2_X1 U767 ( .A1(G8), .A2(n699), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U769 ( .A1(n702), .A2(n705), .ZN(n707) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U771 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  OR2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n745) );
  XNOR2_X1 U775 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  XNOR2_X1 U776 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n720) );
  NAND2_X1 U777 ( .A1(G116), .A2(n902), .ZN(n711) );
  NAND2_X1 U778 ( .A1(G128), .A2(n903), .ZN(n710) );
  NAND2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U780 ( .A(KEYINPUT35), .B(n712), .ZN(n718) );
  NAND2_X1 U781 ( .A1(G140), .A2(n527), .ZN(n714) );
  NAND2_X1 U782 ( .A1(G104), .A2(n899), .ZN(n713) );
  NAND2_X1 U783 ( .A1(n714), .A2(n713), .ZN(n716) );
  XOR2_X1 U784 ( .A(KEYINPUT34), .B(KEYINPUT92), .Z(n715) );
  XNOR2_X1 U785 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U786 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U787 ( .A(n720), .B(n719), .ZN(n896) );
  NOR2_X1 U788 ( .A1(n758), .A2(n896), .ZN(n941) );
  NOR2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n760) );
  NAND2_X1 U790 ( .A1(n941), .A2(n760), .ZN(n723) );
  XNOR2_X1 U791 ( .A(n723), .B(KEYINPUT94), .ZN(n756) );
  XOR2_X1 U792 ( .A(KEYINPUT98), .B(G1991), .Z(n962) );
  NAND2_X1 U793 ( .A1(G131), .A2(n527), .ZN(n725) );
  NAND2_X1 U794 ( .A1(G95), .A2(n899), .ZN(n724) );
  NAND2_X1 U795 ( .A1(n725), .A2(n724), .ZN(n732) );
  NAND2_X1 U796 ( .A1(n903), .A2(G119), .ZN(n726) );
  XNOR2_X1 U797 ( .A(KEYINPUT95), .B(n726), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n902), .A2(G107), .ZN(n727) );
  XOR2_X1 U799 ( .A(KEYINPUT96), .B(n727), .Z(n728) );
  NOR2_X1 U800 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U801 ( .A(n730), .B(KEYINPUT97), .ZN(n731) );
  NOR2_X1 U802 ( .A1(n732), .A2(n731), .ZN(n895) );
  NOR2_X1 U803 ( .A1(n962), .A2(n895), .ZN(n741) );
  NAND2_X1 U804 ( .A1(G141), .A2(n527), .ZN(n734) );
  NAND2_X1 U805 ( .A1(G117), .A2(n902), .ZN(n733) );
  NAND2_X1 U806 ( .A1(n734), .A2(n733), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n899), .A2(G105), .ZN(n735) );
  XOR2_X1 U808 ( .A(KEYINPUT38), .B(n735), .Z(n736) );
  NOR2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n739) );
  NAND2_X1 U810 ( .A1(n903), .A2(G129), .ZN(n738) );
  NAND2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n914) );
  AND2_X1 U812 ( .A1(n914), .A2(G1996), .ZN(n740) );
  NOR2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n938) );
  INV_X1 U814 ( .A(n760), .ZN(n742) );
  NOR2_X1 U815 ( .A1(n938), .A2(n742), .ZN(n752) );
  INV_X1 U816 ( .A(n752), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n756), .A2(n743), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n748) );
  XOR2_X1 U819 ( .A(G1986), .B(G290), .Z(n746) );
  XNOR2_X1 U820 ( .A(KEYINPUT91), .B(n746), .ZN(n1002) );
  NAND2_X1 U821 ( .A1(n1002), .A2(n760), .ZN(n747) );
  NAND2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n763) );
  XOR2_X1 U823 ( .A(KEYINPUT39), .B(KEYINPUT109), .Z(n755) );
  NOR2_X1 U824 ( .A1(G1996), .A2(n914), .ZN(n945) );
  NAND2_X1 U825 ( .A1(n962), .A2(n895), .ZN(n749) );
  XOR2_X1 U826 ( .A(KEYINPUT108), .B(n749), .Z(n952) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U828 ( .A1(n952), .A2(n750), .ZN(n751) );
  NOR2_X1 U829 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U830 ( .A1(n945), .A2(n753), .ZN(n754) );
  XNOR2_X1 U831 ( .A(n755), .B(n754), .ZN(n757) );
  NAND2_X1 U832 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U833 ( .A1(n758), .A2(n896), .ZN(n943) );
  NAND2_X1 U834 ( .A1(n759), .A2(n943), .ZN(n761) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U836 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U837 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n764) );
  XNOR2_X1 U838 ( .A(n765), .B(n764), .ZN(G329) );
  INV_X1 U839 ( .A(G120), .ZN(G236) );
  INV_X1 U840 ( .A(G69), .ZN(G235) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  NAND2_X1 U843 ( .A1(G94), .A2(G452), .ZN(n766) );
  XOR2_X1 U844 ( .A(KEYINPUT70), .B(n766), .Z(G173) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U846 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U847 ( .A(G567), .ZN(n834) );
  NOR2_X1 U848 ( .A1(G223), .A2(n834), .ZN(n769) );
  XNOR2_X1 U849 ( .A(KEYINPUT72), .B(KEYINPUT11), .ZN(n768) );
  XNOR2_X1 U850 ( .A(n769), .B(n768), .ZN(G234) );
  INV_X1 U851 ( .A(G860), .ZN(n778) );
  OR2_X1 U852 ( .A1(n987), .A2(n778), .ZN(G153) );
  INV_X1 U853 ( .A(G868), .ZN(n820) );
  NAND2_X1 U854 ( .A1(n770), .A2(n820), .ZN(n771) );
  XNOR2_X1 U855 ( .A(n771), .B(KEYINPUT76), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(G284) );
  INV_X1 U858 ( .A(n989), .ZN(G299) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n774) );
  XOR2_X1 U860 ( .A(KEYINPUT79), .B(n774), .Z(n777) );
  NOR2_X1 U861 ( .A1(G286), .A2(n820), .ZN(n775) );
  XNOR2_X1 U862 ( .A(KEYINPUT78), .B(n775), .ZN(n776) );
  NOR2_X1 U863 ( .A1(n777), .A2(n776), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n778), .A2(G559), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n779), .A2(n988), .ZN(n780) );
  XNOR2_X1 U866 ( .A(n780), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U867 ( .A1(G868), .A2(n987), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G868), .A2(n988), .ZN(n781) );
  NOR2_X1 U869 ( .A1(G559), .A2(n781), .ZN(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(G282) );
  NAND2_X1 U871 ( .A1(G99), .A2(n899), .ZN(n790) );
  NAND2_X1 U872 ( .A1(G135), .A2(n527), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G111), .A2(n902), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n903), .A2(G123), .ZN(n786) );
  XOR2_X1 U876 ( .A(KEYINPUT18), .B(n786), .Z(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U878 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U879 ( .A(n791), .B(KEYINPUT80), .ZN(n937) );
  XNOR2_X1 U880 ( .A(n937), .B(G2096), .ZN(n792) );
  XNOR2_X1 U881 ( .A(n792), .B(KEYINPUT81), .ZN(n794) );
  INV_X1 U882 ( .A(G2100), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(G156) );
  NAND2_X1 U884 ( .A1(G559), .A2(n988), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n795), .B(n987), .ZN(n817) );
  NOR2_X1 U886 ( .A1(n817), .A2(G860), .ZN(n807) );
  NAND2_X1 U887 ( .A1(n796), .A2(G80), .ZN(n797) );
  XNOR2_X1 U888 ( .A(n797), .B(KEYINPUT82), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G93), .A2(n801), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G67), .A2(n802), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n819) );
  XOR2_X1 U895 ( .A(n807), .B(n819), .Z(G145) );
  XNOR2_X1 U896 ( .A(G166), .B(G299), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n808), .B(G305), .ZN(n814) );
  XNOR2_X1 U898 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n809) );
  XNOR2_X1 U899 ( .A(n809), .B(KEYINPUT19), .ZN(n810) );
  XNOR2_X1 U900 ( .A(KEYINPUT84), .B(n810), .ZN(n812) );
  XNOR2_X1 U901 ( .A(G288), .B(KEYINPUT87), .ZN(n811) );
  XNOR2_X1 U902 ( .A(n812), .B(n811), .ZN(n813) );
  XOR2_X1 U903 ( .A(n814), .B(n813), .Z(n816) );
  XOR2_X1 U904 ( .A(G290), .B(n819), .Z(n815) );
  XNOR2_X1 U905 ( .A(n816), .B(n815), .ZN(n921) );
  XNOR2_X1 U906 ( .A(n817), .B(n921), .ZN(n818) );
  NAND2_X1 U907 ( .A1(n818), .A2(G868), .ZN(n822) );
  NAND2_X1 U908 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U909 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U910 ( .A(KEYINPUT88), .B(n823), .ZN(G295) );
  NAND2_X1 U911 ( .A1(G2078), .A2(G2084), .ZN(n824) );
  XOR2_X1 U912 ( .A(KEYINPUT20), .B(n824), .Z(n825) );
  NAND2_X1 U913 ( .A1(G2090), .A2(n825), .ZN(n826) );
  XNOR2_X1 U914 ( .A(KEYINPUT21), .B(n826), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n827), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U916 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U917 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NOR2_X1 U918 ( .A1(G220), .A2(G219), .ZN(n828) );
  XOR2_X1 U919 ( .A(KEYINPUT22), .B(n828), .Z(n829) );
  NOR2_X1 U920 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U921 ( .A1(G96), .A2(n830), .ZN(n856) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n856), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n831), .B(KEYINPUT89), .ZN(n836) );
  NOR2_X1 U924 ( .A1(G237), .A2(G236), .ZN(n832) );
  NAND2_X1 U925 ( .A1(G108), .A2(n832), .ZN(n833) );
  NOR2_X1 U926 ( .A1(G235), .A2(n833), .ZN(n858) );
  NOR2_X1 U927 ( .A1(n834), .A2(n858), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G319) );
  INV_X1 U929 ( .A(G319), .ZN(n838) );
  NAND2_X1 U930 ( .A1(G483), .A2(G661), .ZN(n837) );
  NOR2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n855) );
  NAND2_X1 U932 ( .A1(n855), .A2(G36), .ZN(G176) );
  XOR2_X1 U933 ( .A(G2435), .B(G2454), .Z(n840) );
  XNOR2_X1 U934 ( .A(G1348), .B(G1341), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n850) );
  XOR2_X1 U936 ( .A(KEYINPUT114), .B(KEYINPUT111), .Z(n842) );
  XNOR2_X1 U937 ( .A(G2427), .B(G2451), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U939 ( .A(G2430), .B(G2443), .Z(n844) );
  XNOR2_X1 U940 ( .A(G2438), .B(KEYINPUT113), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U943 ( .A(KEYINPUT112), .B(G2446), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  NAND2_X1 U946 ( .A1(n851), .A2(G14), .ZN(n926) );
  XNOR2_X1 U947 ( .A(KEYINPUT115), .B(n926), .ZN(G401) );
  INV_X1 U948 ( .A(G223), .ZN(n852) );
  NAND2_X1 U949 ( .A1(G2106), .A2(n852), .ZN(G217) );
  AND2_X1 U950 ( .A1(G15), .A2(G2), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G661), .A2(n853), .ZN(G259) );
  NAND2_X1 U952 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U953 ( .A1(n855), .A2(n854), .ZN(G188) );
  INV_X1 U955 ( .A(G96), .ZN(G221) );
  INV_X1 U956 ( .A(n856), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(G261) );
  INV_X1 U958 ( .A(G261), .ZN(G325) );
  XOR2_X1 U959 ( .A(G2096), .B(KEYINPUT43), .Z(n860) );
  XNOR2_X1 U960 ( .A(G2090), .B(KEYINPUT42), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U962 ( .A(n861), .B(G2678), .Z(n863) );
  XNOR2_X1 U963 ( .A(G2067), .B(G2072), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U965 ( .A(KEYINPUT116), .B(G2100), .Z(n865) );
  XNOR2_X1 U966 ( .A(G2078), .B(G2084), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(G227) );
  XOR2_X1 U969 ( .A(G1976), .B(G1956), .Z(n869) );
  XNOR2_X1 U970 ( .A(G1986), .B(G1961), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U972 ( .A(n870), .B(G2474), .Z(n872) );
  XNOR2_X1 U973 ( .A(G1996), .B(G1991), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U975 ( .A(KEYINPUT41), .B(G1981), .Z(n874) );
  XNOR2_X1 U976 ( .A(G1966), .B(G1971), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(G229) );
  NAND2_X1 U979 ( .A1(n903), .A2(G124), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G136), .A2(n527), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(n880), .B(KEYINPUT117), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G112), .A2(n902), .ZN(n882) );
  NAND2_X1 U985 ( .A1(G100), .A2(n899), .ZN(n881) );
  NAND2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U987 ( .A(KEYINPUT118), .B(n883), .Z(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U989 ( .A(n886), .B(KEYINPUT119), .ZN(G162) );
  NAND2_X1 U990 ( .A1(G118), .A2(n902), .ZN(n888) );
  NAND2_X1 U991 ( .A1(G130), .A2(n903), .ZN(n887) );
  NAND2_X1 U992 ( .A1(n888), .A2(n887), .ZN(n893) );
  NAND2_X1 U993 ( .A1(G142), .A2(n527), .ZN(n890) );
  NAND2_X1 U994 ( .A1(G106), .A2(n899), .ZN(n889) );
  NAND2_X1 U995 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U996 ( .A(KEYINPUT45), .B(n891), .Z(n892) );
  NOR2_X1 U997 ( .A1(n893), .A2(n892), .ZN(n894) );
  XNOR2_X1 U998 ( .A(n895), .B(n894), .ZN(n918) );
  XNOR2_X1 U999 ( .A(n937), .B(G164), .ZN(n897) );
  XNOR2_X1 U1000 ( .A(n897), .B(n896), .ZN(n913) );
  XOR2_X1 U1001 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n911) );
  NAND2_X1 U1002 ( .A1(G139), .A2(n527), .ZN(n901) );
  NAND2_X1 U1003 ( .A1(G103), .A2(n899), .ZN(n900) );
  NAND2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(G115), .A2(n902), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(G127), .A2(n903), .ZN(n904) );
  NAND2_X1 U1007 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1008 ( .A(KEYINPUT120), .B(n906), .Z(n907) );
  XNOR2_X1 U1009 ( .A(KEYINPUT47), .B(n907), .ZN(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n932) );
  XNOR2_X1 U1011 ( .A(n932), .B(KEYINPUT121), .ZN(n910) );
  XNOR2_X1 U1012 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1013 ( .A(n913), .B(n912), .Z(n916) );
  XOR2_X1 U1014 ( .A(G160), .B(n914), .Z(n915) );
  XNOR2_X1 U1015 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(G162), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n920), .ZN(G395) );
  XNOR2_X1 U1019 ( .A(n987), .B(n921), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(G171), .B(n988), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1022 ( .A(G286), .B(n924), .Z(n925) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n925), .ZN(G397) );
  NAND2_X1 U1024 ( .A1(G319), .A2(n926), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(G227), .A2(G229), .ZN(n927) );
  XNOR2_X1 U1026 ( .A(KEYINPUT49), .B(n927), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(G395), .A2(G397), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(G225) );
  INV_X1 U1030 ( .A(G225), .ZN(G308) );
  INV_X1 U1031 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1032 ( .A(n932), .B(KEYINPUT123), .Z(n933) );
  XOR2_X1 U1033 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1036 ( .A(KEYINPUT50), .B(n936), .Z(n955) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n940) );
  XOR2_X1 U1038 ( .A(G160), .B(G2084), .Z(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n950) );
  INV_X1 U1040 ( .A(n941), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n948) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(n946), .B(KEYINPUT51), .ZN(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1048 ( .A(KEYINPUT122), .B(n953), .Z(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n956), .ZN(n957) );
  INV_X1 U1051 ( .A(KEYINPUT55), .ZN(n980) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n980), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G29), .ZN(n1038) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G26), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(G28), .A2(n961), .ZN(n964) );
  XOR2_X1 U1058 ( .A(n962), .B(G25), .Z(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(n965), .B(G32), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(G27), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(KEYINPUT53), .B(n971), .ZN(n978) );
  XOR2_X1 U1065 ( .A(KEYINPUT125), .B(G34), .Z(n973) );
  XNOR2_X1 U1066 ( .A(G2084), .B(KEYINPUT54), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(n973), .B(n972), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G35), .B(G2090), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(KEYINPUT124), .B(n974), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(n980), .B(n979), .ZN(n982) );
  INV_X1 U1073 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(G11), .A2(n983), .ZN(n1036) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1009) );
  XOR2_X1 U1077 ( .A(G168), .B(G1966), .Z(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n986), .Z(n1007) );
  XNOR2_X1 U1080 ( .A(n987), .B(G1341), .ZN(n1005) );
  XNOR2_X1 U1081 ( .A(G1348), .B(n988), .ZN(n1000) );
  XNOR2_X1 U1082 ( .A(n989), .B(G1956), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G171), .B(G1961), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1087 ( .A(G1971), .B(G166), .Z(n996) );
  XNOR2_X1 U1088 ( .A(KEYINPUT126), .B(n996), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(KEYINPUT127), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1034) );
  INV_X1 U1096 ( .A(G16), .ZN(n1032) );
  XNOR2_X1 U1097 ( .A(G20), .B(n1010), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1341), .B(G19), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G6), .B(G1981), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XOR2_X1 U1102 ( .A(KEYINPUT59), .B(G1348), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(G4), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1018), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G1966), .B(G21), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(G5), .B(G1961), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1029) );
  XNOR2_X1 U1110 ( .A(G1971), .B(G22), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(G23), .B(G1976), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XOR2_X1 U1113 ( .A(G1986), .B(G24), .Z(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT58), .B(n1027), .ZN(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1117 ( .A(KEYINPUT61), .B(n1030), .ZN(n1031) );
  NAND2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1119 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1120 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1121 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1039), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

