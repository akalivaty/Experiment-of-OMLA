//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT64), .Z(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT65), .ZN(new_n228));
  XOR2_X1   g0028(.A(G264), .B(G270), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n202), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n238), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(new_n206), .A2(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT68), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  AND2_X1   g0049(.A1(new_n249), .A2(new_n215), .ZN(new_n250));
  INV_X1    g0050(.A(G13), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n248), .A2(new_n254), .B1(G50), .B2(new_n253), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n203), .A2(G20), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n250), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT9), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n258), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n269), .B2(new_n270), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT67), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n267), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(G222), .A3(new_n275), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n271), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n266), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G41), .A2(G45), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G1), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n206), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  INV_X1    g0088(.A(new_n215), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n206), .A2(new_n296), .B1(new_n289), .B2(new_n290), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n293), .B1(G226), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n282), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G190), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(G200), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n265), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT72), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(KEYINPUT72), .A3(KEYINPUT10), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n265), .A2(new_n302), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT71), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .A4(new_n301), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT71), .B1(new_n303), .B2(KEYINPUT10), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n306), .A2(new_n307), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n264), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n300), .A2(G169), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  AOI211_X1 g0116(.A(new_n314), .B(new_n315), .C1(new_n316), .C2(new_n300), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT16), .ZN(new_n319));
  OR2_X1    g0119(.A1(KEYINPUT74), .A2(G33), .ZN(new_n320));
  NAND2_X1  g0120(.A1(KEYINPUT74), .A2(G33), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n268), .A3(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n270), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n270), .A2(new_n207), .ZN(new_n326));
  NOR2_X1   g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n240), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(G58), .A2(G68), .ZN(new_n330));
  OAI21_X1  g0130(.A(G20), .B1(new_n330), .B2(new_n201), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT75), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n260), .A2(G159), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT75), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n334), .B(G20), .C1(new_n330), .C2(new_n201), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n319), .B1(new_n329), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n249), .A2(new_n215), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT74), .B(G33), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n327), .B1(new_n339), .B2(KEYINPUT3), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n325), .B1(new_n340), .B2(new_n207), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT74), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT74), .A2(G33), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT3), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n344), .A2(new_n325), .A3(new_n207), .A4(new_n269), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G68), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n332), .A2(KEYINPUT16), .A3(new_n333), .A4(new_n335), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n337), .B(new_n338), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n256), .B1(new_n206), .B2(G20), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n251), .A2(new_n207), .A3(G1), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n338), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n350), .A2(new_n352), .B1(new_n351), .B2(new_n256), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n287), .A2(new_n291), .B1(new_n297), .B2(G232), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n344), .A2(new_n269), .ZN(new_n356));
  MUX2_X1   g0156(.A(G223), .B(G226), .S(G1698), .Z(new_n357));
  AOI22_X1  g0157(.A1(new_n356), .A2(new_n357), .B1(G33), .B2(G87), .ZN(new_n358));
  INV_X1    g0158(.A(new_n266), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G169), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n360), .B2(new_n316), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n354), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT18), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n353), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n344), .A2(new_n207), .A3(new_n269), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT7), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(G68), .A3(new_n345), .ZN(new_n369));
  INV_X1    g0169(.A(new_n348), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n250), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n371), .B2(new_n337), .ZN(new_n372));
  INV_X1    g0172(.A(G200), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n268), .B1(new_n320), .B2(new_n321), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n357), .B1(new_n374), .B2(new_n327), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G87), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n359), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n297), .A2(G232), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n292), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n373), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(G190), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n355), .B(new_n381), .C1(new_n358), .C2(new_n359), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT76), .B1(new_n372), .B2(new_n383), .ZN(new_n384));
  AND4_X1   g0184(.A1(KEYINPUT76), .A2(new_n383), .A3(new_n349), .A4(new_n353), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT17), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n349), .A3(new_n353), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n365), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  INV_X1    g0191(.A(new_n270), .ZN(new_n392));
  OAI211_X1 g0192(.A(G232), .B(G1698), .C1(new_n392), .C2(new_n327), .ZN(new_n393));
  OAI211_X1 g0193(.A(G226), .B(new_n275), .C1(new_n392), .C2(new_n327), .ZN(new_n394));
  INV_X1    g0194(.A(G97), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(new_n394), .C1(new_n258), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n266), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n287), .A2(new_n291), .B1(new_n297), .B2(G238), .ZN(new_n398));
  AOI211_X1 g0198(.A(KEYINPUT73), .B(new_n391), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n397), .A2(new_n391), .A3(new_n398), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(new_n316), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT73), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n397), .A2(new_n391), .A3(new_n398), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT14), .B1(new_n408), .B2(G169), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT14), .B(G169), .C1(new_n401), .C2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n406), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n351), .A2(new_n240), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT12), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n240), .ZN(new_n416));
  INV_X1    g0216(.A(new_n259), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n280), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .A3(new_n338), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n352), .A2(G68), .A3(new_n246), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n415), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT11), .B1(new_n418), .B2(new_n338), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n413), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(G200), .B1(new_n401), .B2(new_n410), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n400), .A2(new_n405), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n407), .A2(G190), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n423), .B(new_n426), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n260), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n256), .A2(new_n430), .B1(new_n207), .B2(new_n280), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n417), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n338), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT69), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n280), .B1(new_n206), .B2(G20), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n352), .A2(new_n437), .B1(new_n280), .B2(new_n351), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(G238), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n274), .B2(new_n277), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n271), .A2(G232), .A3(new_n275), .ZN(new_n443));
  INV_X1    g0243(.A(G107), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n271), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n266), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n293), .B1(G244), .B2(new_n297), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(G190), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n446), .A2(new_n447), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n440), .B(new_n448), .C1(new_n373), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT70), .B1(new_n449), .B2(G169), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n316), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT70), .A4(new_n316), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n439), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  AND4_X1   g0256(.A1(new_n425), .A2(new_n429), .A3(new_n450), .A4(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n318), .A2(new_n390), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT85), .ZN(new_n460));
  NAND2_X1  g0260(.A1(KEYINPUT22), .A2(G87), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n340), .A2(G20), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n339), .A2(new_n207), .A3(G116), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT23), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(new_n207), .B2(G107), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n444), .A2(KEYINPUT23), .A3(G20), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n207), .A2(G87), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n269), .B2(new_n270), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n463), .B(new_n467), .C1(KEYINPUT22), .C2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n460), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n356), .A2(KEYINPUT22), .A3(new_n207), .A4(G87), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n469), .A2(KEYINPUT22), .ZN(new_n473));
  INV_X1    g0273(.A(G116), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n320), .B2(new_n321), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n475), .A2(new_n207), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n472), .A2(KEYINPUT85), .A3(new_n473), .A4(new_n476), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n471), .A2(KEYINPUT24), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n338), .B1(new_n471), .B2(KEYINPUT24), .ZN(new_n479));
  OR2_X1    g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n254), .B1(new_n206), .B2(G33), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT25), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n253), .B2(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n351), .A2(KEYINPUT25), .A3(new_n444), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n481), .A2(G107), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G250), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n275), .ZN(new_n487));
  INV_X1    g0287(.A(G257), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G1698), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n344), .B2(new_n269), .ZN(new_n491));
  INV_X1    g0291(.A(G294), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n320), .B2(new_n321), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT86), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT86), .ZN(new_n495));
  INV_X1    g0295(.A(new_n493), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n340), .C2(new_n490), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n497), .A3(new_n266), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n295), .A2(G1), .ZN(new_n499));
  XNOR2_X1  g0299(.A(KEYINPUT5), .B(G41), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n266), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G264), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n500), .A2(new_n499), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n291), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n498), .A2(G190), .A3(new_n502), .A4(new_n504), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n480), .A2(new_n485), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n485), .B1(new_n478), .B2(new_n479), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n505), .A2(KEYINPUT87), .A3(G169), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n498), .A2(G179), .A3(new_n502), .A4(new_n504), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT87), .B1(new_n505), .B2(G169), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT21), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT82), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n517), .B1(new_n253), .B2(G116), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n351), .A2(KEYINPUT82), .A3(new_n474), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n481), .A2(G116), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n207), .C1(G33), .C2(new_n395), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n474), .A2(G20), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n338), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT83), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g0326(.A1(new_n338), .A2(new_n523), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT20), .A4(new_n522), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n525), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n520), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n501), .A2(G270), .B1(new_n503), .B2(new_n291), .ZN(new_n533));
  INV_X1    g0333(.A(G264), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G257), .B2(G1698), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(new_n269), .B2(new_n344), .ZN(new_n537));
  INV_X1    g0337(.A(G303), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n271), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n266), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G169), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n516), .B1(new_n532), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n520), .A2(new_n531), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n533), .A2(new_n540), .A3(G179), .ZN(new_n545));
  NAND2_X1  g0345(.A1(KEYINPUT21), .A2(G169), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n533), .B2(new_n540), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n541), .A2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n533), .A2(new_n540), .A3(G190), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n532), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n543), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT84), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n543), .A2(new_n551), .A3(KEYINPUT84), .A4(new_n548), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n475), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n441), .A2(new_n275), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G244), .B2(new_n275), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n340), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n266), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT79), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n499), .B(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n266), .A2(new_n486), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(new_n499), .B2(new_n291), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  AOI21_X1  g0367(.A(G20), .B1(new_n344), .B2(new_n269), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G68), .ZN(new_n569));
  NOR3_X1   g0369(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(G33), .B2(G97), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT19), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n259), .A2(new_n573), .A3(G97), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n576), .A2(new_n338), .B1(new_n351), .B2(new_n432), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n481), .A2(G87), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n561), .A2(G190), .A3(new_n565), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n567), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n432), .A2(new_n351), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n352), .B1(G1), .B2(new_n258), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n568), .A2(G68), .B1(new_n572), .B2(new_n574), .ZN(new_n583));
  OAI221_X1 g0383(.A(new_n581), .B1(new_n582), .B2(new_n432), .C1(new_n583), .C2(new_n250), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT81), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G169), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n566), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n576), .A2(new_n338), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n582), .A2(new_n432), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n589), .A2(KEYINPUT81), .A3(new_n581), .A4(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n586), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n561), .A2(new_n316), .A3(new_n565), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT80), .ZN(new_n594));
  XNOR2_X1  g0394(.A(new_n593), .B(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n580), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n395), .A2(new_n444), .ZN(new_n598));
  NOR2_X1   g0398(.A1(G97), .A2(G107), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(KEYINPUT6), .A2(G97), .ZN(new_n601));
  OR3_X1    g0401(.A1(new_n601), .A2(KEYINPUT77), .A3(G107), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT77), .B1(new_n601), .B2(G107), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G20), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n260), .A2(G77), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n324), .A2(new_n328), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n444), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n338), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT78), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n253), .B2(G97), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n351), .A2(KEYINPUT78), .A3(new_n395), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n582), .B2(new_n395), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n501), .A2(G257), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n504), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT4), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n275), .A2(G244), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n340), .B2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n275), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n276), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n618), .B1(new_n624), .B2(new_n266), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n316), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(new_n521), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n359), .B1(new_n629), .B2(new_n621), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n587), .B1(new_n630), .B2(new_n618), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n616), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n618), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n356), .A2(G244), .A3(new_n275), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n619), .B2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(G190), .B(new_n633), .C1(new_n635), .C2(new_n359), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n614), .B1(new_n608), .B2(new_n338), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(new_n373), .C2(new_n625), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n596), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n556), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n459), .A2(new_n515), .A3(new_n641), .ZN(G372));
  INV_X1    g0442(.A(new_n456), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n643), .A2(new_n429), .B1(new_n424), .B2(new_n413), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n386), .A2(new_n389), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n365), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n306), .A2(new_n307), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n311), .A2(new_n312), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n317), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n543), .A2(new_n548), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n514), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT88), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n514), .A2(KEYINPUT88), .A3(new_n651), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n485), .B(new_n507), .C1(new_n478), .C2(new_n479), .ZN(new_n656));
  INV_X1    g0456(.A(new_n506), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n586), .A2(new_n588), .A3(new_n591), .A4(new_n593), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n580), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n658), .A2(new_n660), .A3(new_n639), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n654), .A2(new_n655), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  INV_X1    g0463(.A(new_n580), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n588), .B1(new_n584), .B2(new_n585), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT81), .B1(new_n577), .B2(new_n590), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n593), .B(KEYINPUT80), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n616), .A2(new_n626), .A3(new_n631), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(new_n663), .A3(new_n580), .A4(new_n659), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n659), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n662), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n650), .B1(new_n459), .B2(new_n676), .ZN(G369));
  NAND2_X1  g0477(.A1(new_n252), .A2(new_n207), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G213), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(KEYINPUT27), .B2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n532), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n556), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n651), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n682), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n515), .B1(new_n509), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n514), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n651), .A2(new_n688), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n515), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n690), .B2(new_n682), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n210), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n570), .A2(new_n474), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n698), .A2(new_n699), .A3(new_n206), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n214), .B2(new_n698), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NOR2_X1   g0502(.A1(new_n658), .A2(new_n639), .ZN(new_n703));
  INV_X1    g0503(.A(new_n660), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(new_n652), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n667), .A2(new_n668), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n706), .A2(new_n663), .A3(new_n580), .A4(new_n670), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT26), .B1(new_n660), .B2(new_n632), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n659), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n682), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n688), .B1(new_n662), .B2(new_n674), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  MUX2_X1   g0512(.A(new_n710), .B(new_n711), .S(new_n712), .Z(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n561), .A2(new_n565), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n625), .A2(new_n715), .A3(new_n545), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n498), .A2(new_n502), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n566), .A2(new_n541), .A3(new_n316), .ZN(new_n719));
  INV_X1    g0519(.A(new_n717), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n719), .A2(KEYINPUT30), .A3(new_n720), .A4(new_n625), .ZN(new_n721));
  INV_X1    g0521(.A(new_n625), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n533), .B2(new_n540), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(new_n505), .A3(new_n566), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n718), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n726), .A2(KEYINPUT89), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(KEYINPUT89), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n725), .B2(new_n688), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n513), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n511), .A3(new_n510), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n658), .B1(new_n733), .B2(new_n509), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n556), .A3(new_n640), .A4(new_n682), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n713), .B1(G330), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n702), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n251), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n206), .B1(new_n740), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n698), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n686), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT90), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n207), .A2(new_n316), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n749), .B1(new_n751), .B2(new_n373), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n750), .A2(KEYINPUT90), .A3(G200), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(G190), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n381), .A2(G179), .A3(G200), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n207), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(G326), .B1(G294), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT93), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n751), .A2(new_n381), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n207), .A2(G179), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n762), .A2(G322), .B1(G329), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n271), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n750), .A2(new_n764), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n763), .A2(new_n381), .A3(G200), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n772), .A2(new_n773), .B1(new_n774), .B2(new_n538), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n761), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n752), .A2(new_n381), .A3(new_n753), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT92), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(G317), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n781), .A2(new_n783), .B1(new_n759), .B2(new_n760), .ZN(new_n784));
  INV_X1    g0584(.A(new_n774), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n766), .A2(G159), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT91), .B(KEYINPUT32), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n786), .B1(new_n395), .B2(new_n757), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n773), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n787), .A2(new_n788), .B1(G107), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n770), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n768), .B1(new_n792), .B2(G77), .ZN(new_n793));
  INV_X1    g0593(.A(G58), .ZN(new_n794));
  INV_X1    g0594(.A(new_n762), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n791), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n789), .B(new_n796), .C1(G50), .C2(new_n755), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n781), .A2(G68), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n776), .A2(new_n784), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n215), .B1(G20), .B2(new_n587), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n210), .A2(G116), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n244), .A2(new_n295), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n697), .A2(new_n356), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n805), .C1(new_n295), .C2(new_n214), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n697), .A2(new_n768), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n802), .B(new_n806), .C1(G355), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n746), .A2(new_n800), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n799), .A2(new_n801), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n743), .B1(new_n748), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G330), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n686), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n812), .B1(new_n814), .B2(new_n743), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT95), .Z(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n439), .A2(new_n688), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n453), .A2(new_n455), .B1(new_n450), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n453), .A2(new_n455), .A3(new_n682), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n711), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n737), .A2(G330), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n743), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n757), .A2(new_n395), .B1(new_n774), .B2(new_n444), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n768), .B1(new_n474), .B2(new_n770), .C1(new_n795), .C2(new_n492), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G303), .C2(new_n755), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n790), .A2(G87), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(new_n769), .B2(new_n765), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT96), .ZN(new_n831));
  INV_X1    g0631(.A(new_n781), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n828), .B(new_n831), .C1(new_n772), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n755), .A2(G137), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n762), .A2(G143), .B1(G159), .B2(new_n792), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n835), .C1(new_n832), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  NOR2_X1   g0638(.A1(new_n773), .A2(new_n240), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G58), .B2(new_n758), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n340), .B1(G132), .B2(new_n766), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(new_n202), .C2(new_n774), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n833), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n800), .ZN(new_n844));
  INV_X1    g0644(.A(new_n743), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n800), .A2(new_n744), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n280), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(new_n847), .C1(new_n745), .C2(new_n821), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n825), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  NOR2_X1   g0650(.A1(new_n365), .A2(new_n681), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT76), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n387), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT37), .B1(new_n354), .B2(new_n362), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n372), .A2(KEYINPUT76), .A3(new_n383), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n354), .A2(new_n681), .ZN(new_n857));
  AND4_X1   g0657(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n384), .A2(new_n385), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n338), .B1(new_n347), .B2(new_n348), .ZN(new_n860));
  INV_X1    g0660(.A(new_n336), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT16), .B1(new_n369), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n353), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT98), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT98), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n353), .C1(new_n860), .C2(new_n862), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n362), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n864), .A2(new_n681), .A3(new_n866), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n859), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n858), .B1(new_n869), .B2(KEYINPUT37), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT99), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n365), .A2(new_n386), .A3(new_n389), .ZN(new_n872));
  INV_X1    g0672(.A(new_n868), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n870), .A2(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n869), .A2(KEYINPUT37), .ZN(new_n875));
  INV_X1    g0675(.A(new_n858), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT99), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n874), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n874), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n423), .A2(new_n682), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(G169), .B1(new_n401), .B2(new_n410), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT14), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT73), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n410), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n399), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n886), .A2(new_n411), .B1(new_n889), .B2(new_n402), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n429), .B(new_n883), .C1(new_n890), .C2(new_n423), .ZN(new_n891));
  NOR3_X1   g0691(.A1(new_n888), .A2(new_n399), .A3(new_n428), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n426), .A2(new_n423), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n882), .B1(new_n413), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n891), .A2(new_n895), .A3(KEYINPUT97), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n890), .A2(new_n429), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT97), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n897), .A2(new_n898), .A3(new_n882), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n453), .A2(new_n455), .A3(new_n682), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n450), .A2(new_n818), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n902), .B1(new_n643), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n688), .B(new_n904), .C1(new_n662), .C2(new_n674), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n905), .B2(new_n820), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n852), .B1(new_n881), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n874), .A2(new_n878), .A3(KEYINPUT38), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n363), .A2(new_n387), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n910), .B2(new_n857), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n390), .B2(new_n857), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n858), .A2(KEYINPUT38), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT39), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT100), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT39), .B1(new_n879), .B2(new_n880), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n908), .A2(new_n914), .A3(KEYINPUT100), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n425), .A2(new_n688), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n907), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n713), .A2(new_n458), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n923), .A2(new_n650), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n688), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n729), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(new_n735), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n896), .A2(new_n821), .A3(new_n899), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n928), .A2(KEYINPUT101), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT101), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n896), .A2(new_n821), .A3(new_n899), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n927), .A2(new_n735), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT38), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n872), .A2(new_n873), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n877), .B2(KEYINPUT99), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n870), .A2(new_n871), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n908), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT40), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n912), .A2(new_n913), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n908), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n928), .A2(new_n945), .A3(new_n929), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n942), .A2(new_n948), .B1(new_n459), .B2(new_n928), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT101), .B1(new_n928), .B2(new_n929), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n932), .A2(new_n931), .A3(new_n933), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n945), .B1(new_n881), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n953), .A2(new_n458), .A3(new_n933), .A4(new_n947), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n949), .A2(new_n954), .A3(G330), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n925), .A2(new_n955), .B1(new_n206), .B2(new_n740), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT102), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n925), .A2(new_n955), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n604), .A2(KEYINPUT35), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n604), .A2(KEYINPUT35), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n962), .A2(G116), .A3(new_n216), .A4(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT36), .ZN(new_n965));
  OAI21_X1  g0765(.A(G77), .B1(new_n794), .B2(new_n240), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n239), .B1(new_n966), .B2(new_n213), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(G1), .A3(new_n251), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n961), .A2(new_n965), .A3(new_n968), .ZN(G367));
  NAND2_X1  g0769(.A1(new_n577), .A2(new_n578), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n688), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n704), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n659), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n632), .B(new_n638), .C1(new_n637), .C2(new_n682), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n670), .A2(new_n688), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n694), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT42), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n632), .B1(new_n976), .B2(new_n514), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n682), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT103), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n983), .A2(KEYINPUT103), .B1(KEYINPUT42), .B2(new_n979), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n975), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n692), .B1(new_n976), .B2(new_n977), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n698), .B(KEYINPUT41), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n694), .B1(new_n691), .B2(new_n693), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(new_n687), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n738), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(KEYINPUT104), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT104), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n738), .A2(new_n997), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n695), .A2(new_n978), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT45), .Z(new_n1004));
  NOR2_X1   g0804(.A1(new_n695), .A2(new_n978), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT44), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(new_n692), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n995), .B1(new_n1009), .B2(new_n738), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n994), .B1(new_n1010), .B2(new_n742), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(KEYINPUT105), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT105), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n994), .C1(new_n1010), .C2(new_n742), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n230), .A2(new_n804), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n809), .B1(new_n210), .B2(new_n432), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n743), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n758), .A2(G68), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n794), .B2(new_n774), .C1(new_n280), .C2(new_n773), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n271), .B1(new_n770), .B2(new_n202), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(KEYINPUT106), .B(G137), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n795), .A2(new_n836), .B1(new_n765), .B2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(G143), .ZN(new_n1025));
  INV_X1    g0825(.A(G159), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1024), .B1(new_n1025), .B2(new_n754), .C1(new_n832), .C2(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n762), .A2(G303), .B1(G283), .B2(new_n792), .ZN(new_n1028));
  INV_X1    g0828(.A(G317), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1029), .B2(new_n765), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n785), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT46), .B1(new_n785), .B2(G116), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n790), .A2(G97), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1034), .B(new_n340), .C1(new_n444), .C2(new_n757), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G311), .B2(new_n755), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1033), .B(new_n1036), .C1(new_n832), .C2(new_n492), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1027), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT47), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1018), .B1(new_n1039), .B2(new_n800), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n972), .A2(new_n746), .A3(new_n973), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1015), .A2(new_n1042), .ZN(G387));
  NAND2_X1  g0843(.A1(new_n999), .A2(new_n1001), .ZN(new_n1044));
  AOI21_X1  g0844(.A(KEYINPUT109), .B1(new_n1044), .B2(new_n698), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n698), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT109), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n738), .A2(new_n997), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT110), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n807), .A2(new_n699), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(G107), .B2(new_n210), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n234), .A2(G45), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n256), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n805), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1053), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n743), .B1(new_n1059), .B2(new_n810), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1034), .B1(new_n280), .B2(new_n774), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n340), .B(new_n1061), .C1(G150), .C2(new_n766), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT107), .Z(new_n1063));
  NOR2_X1   g0863(.A1(new_n757), .A2(new_n432), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n795), .A2(new_n202), .B1(new_n770), .B2(new_n240), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n755), .C2(G159), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1063), .B(new_n1066), .C1(new_n256), .C2(new_n832), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n356), .B1(G326), .B2(new_n766), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n757), .A2(new_n772), .B1(new_n774), .B2(new_n492), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n755), .A2(G322), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n762), .A2(G317), .B1(G303), .B2(new_n792), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n832), .C2(new_n769), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT49), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1068), .B1(new_n474), .B2(new_n773), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1067), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1060), .B1(new_n1079), .B2(new_n800), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n691), .A2(new_n746), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT108), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n997), .A2(new_n742), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1051), .A2(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n1008), .A2(new_n742), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n809), .B1(new_n395), .B2(new_n210), .C1(new_n805), .C2(new_n238), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n743), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n754), .A2(new_n836), .B1(new_n795), .B2(new_n1026), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n829), .B1(new_n240), .B2(new_n774), .C1(new_n280), .C2(new_n757), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n770), .A2(new_n256), .B1(new_n765), .B2(new_n1025), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1093), .A2(new_n340), .A3(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1092), .B(new_n1095), .C1(new_n202), .C2(new_n832), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n768), .B1(new_n770), .B2(new_n492), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n758), .A2(G116), .B1(new_n790), .B2(G107), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n772), .B2(new_n774), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(G322), .C2(new_n766), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n538), .B2(new_n832), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n754), .A2(new_n1029), .B1(new_n795), .B2(new_n769), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT52), .Z(new_n1103));
  OAI21_X1  g0903(.A(new_n1096), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1090), .B1(new_n1104), .B2(new_n800), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n978), .B2(new_n747), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1088), .A2(new_n1106), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n698), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1002), .B2(new_n1008), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G390));
  INV_X1    g0912(.A(KEYINPUT114), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n921), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n820), .B1(new_n711), .B2(new_n821), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n900), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n917), .A2(new_n918), .A3(new_n1116), .A4(new_n919), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n921), .B1(new_n908), .B2(new_n943), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n819), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n682), .B(new_n1119), .C1(new_n705), .C2(new_n709), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n902), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT111), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT111), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(new_n1123), .A3(new_n902), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n900), .B(KEYINPUT112), .Z(new_n1126));
  OAI21_X1  g0926(.A(new_n1118), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1117), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n928), .A2(new_n813), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n932), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT113), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n821), .C1(new_n731), .C2(new_n736), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1134), .A2(new_n900), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1117), .A2(new_n1127), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT113), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1128), .A2(new_n1137), .A3(new_n1131), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1113), .B1(new_n1139), .B2(new_n741), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1136), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1137), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1143), .A2(KEYINPUT114), .A3(new_n742), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n458), .A2(new_n1129), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n923), .A2(new_n1146), .A3(new_n650), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1126), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n928), .A2(new_n813), .A3(new_n904), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1135), .B(new_n1125), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1134), .A2(new_n900), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1131), .A2(new_n1151), .B1(new_n820), .B2(new_n905), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1147), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1133), .A2(new_n1136), .A3(new_n1138), .A4(new_n1153), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1155), .A2(new_n698), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n845), .B1(new_n256), .B2(new_n846), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT115), .Z(new_n1159));
  OAI22_X1  g0959(.A1(new_n795), .A2(new_n474), .B1(new_n770), .B2(new_n395), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n271), .B(new_n1160), .C1(G294), .C2(new_n766), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n786), .B1(new_n240), .B2(new_n773), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G77), .B2(new_n758), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(new_n772), .C2(new_n754), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G107), .B2(new_n781), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT116), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n832), .A2(new_n1022), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n762), .A2(G132), .ZN(new_n1168));
  INV_X1    g0968(.A(G125), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1168), .B1(new_n1169), .B2(new_n765), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT54), .B(G143), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n271), .B1(new_n770), .B2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n757), .A2(new_n1026), .B1(new_n773), .B2(new_n202), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n755), .A2(G128), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n774), .A2(new_n836), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT53), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1166), .B1(new_n1167), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(KEYINPUT116), .B2(new_n1165), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1159), .B1(new_n801), .B2(new_n1180), .C1(new_n920), .C2(new_n745), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1145), .A2(new_n1157), .A3(new_n1181), .ZN(G378));
  XNOR2_X1  g0982(.A(new_n1147), .B(KEYINPUT121), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1156), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT119), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n264), .A2(new_n681), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n313), .B2(new_n317), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n317), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n649), .A2(new_n1189), .A3(new_n1186), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1188), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n947), .A2(G330), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n942), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n813), .B1(new_n944), .B2(new_n946), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1195), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1192), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n953), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1198), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1185), .B1(new_n1204), .B2(new_n922), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT120), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n942), .A2(new_n1197), .A3(new_n1196), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1202), .B1(new_n953), .B2(new_n1199), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1206), .B(new_n922), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1206), .B1(new_n1204), .B2(new_n922), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1205), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n922), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT119), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n922), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT120), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1215), .A2(new_n1217), .A3(new_n1209), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1184), .A2(new_n1212), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT57), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1220), .B1(new_n1222), .B2(new_n1216), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1109), .B1(new_n1184), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1221), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1212), .A2(new_n1218), .A3(new_n742), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n766), .A2(G283), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n432), .B2(new_n770), .C1(new_n795), .C2(new_n444), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1019), .B1(new_n794), .B2(new_n773), .C1(new_n280), .C2(new_n774), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n340), .A2(new_n294), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n474), .B2(new_n754), .C1(new_n395), .C2(new_n832), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT58), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G50), .B1(new_n258), .B2(new_n294), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1234), .B(new_n1235), .C1(new_n1230), .C2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G33), .B(G41), .C1(new_n766), .C2(G124), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n1026), .B2(new_n773), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n762), .A2(G128), .B1(G137), .B2(new_n792), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n774), .B2(new_n1171), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n781), .B2(G132), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n754), .A2(new_n1169), .B1(new_n836), .B2(new_n757), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT117), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1239), .B1(new_n1245), .B2(KEYINPUT59), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(KEYINPUT59), .B2(new_n1245), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n801), .B1(new_n1237), .B2(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT118), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n845), .B1(new_n202), .B2(new_n846), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n1196), .C2(new_n745), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1226), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1225), .A2(new_n1252), .ZN(G375));
  XOR2_X1   g1053(.A(new_n995), .B(KEYINPUT122), .Z(new_n1254));
  NOR2_X1   g1054(.A1(new_n1153), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1147), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT123), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1064), .B1(G283), .B2(new_n762), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT124), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n768), .B1(new_n770), .B2(new_n444), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n280), .A2(new_n773), .B1(new_n774), .B2(new_n395), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(G303), .C2(new_n766), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1261), .B(new_n1264), .C1(new_n492), .C2(new_n754), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n832), .A2(new_n474), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n832), .A2(new_n1171), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G150), .A2(new_n792), .B1(new_n766), .B2(G128), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n795), .B2(new_n1022), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n755), .A2(G132), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n340), .B1(G58), .B2(new_n790), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n758), .A2(G50), .B1(new_n785), .B2(G159), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1273), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1265), .A2(new_n1266), .B1(new_n1267), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n800), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n845), .B1(new_n240), .B2(new_n846), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(new_n1148), .C2(new_n745), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1257), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(new_n741), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1259), .A2(new_n1281), .ZN(G381));
  NAND3_X1  g1082(.A1(new_n1051), .A2(new_n816), .A3(new_n1086), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1111), .A2(new_n849), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(G387), .A2(G381), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1145), .A2(new_n1157), .A3(new_n1181), .ZN(new_n1286));
  INV_X1    g1086(.A(G375), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(new_n1286), .A3(new_n1287), .ZN(G407));
  INV_X1    g1088(.A(G343), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(G213), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1286), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  NAND2_X1  g1093(.A1(G387), .A2(new_n1111), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G393), .A2(G396), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1295), .A2(new_n1283), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1015), .A2(new_n1042), .A3(G390), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1294), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1295), .A2(new_n1283), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G390), .B1(new_n1015), .B2(new_n1042), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1042), .ZN(new_n1301));
  AOI211_X1 g1101(.A(new_n1301), .B(new_n1111), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1299), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT63), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1225), .A2(G378), .A3(new_n1252), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1222), .A2(new_n1216), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n742), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1251), .B(new_n1308), .C1(new_n1219), .C2(new_n1254), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1286), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1306), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1279), .A2(KEYINPUT60), .A3(new_n1147), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(KEYINPUT125), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT60), .B1(new_n1279), .B2(new_n1147), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1314), .A2(new_n1109), .A3(new_n1153), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G384), .B1(new_n1316), .B2(new_n1281), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n849), .B(new_n1280), .C1(new_n1313), .C2(new_n1315), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1311), .A2(new_n1290), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1304), .B1(new_n1305), .B2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1291), .B1(new_n1306), .B2(new_n1310), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1311), .A2(new_n1290), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1317), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1318), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1291), .A2(G2897), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1325), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(G2897), .B(new_n1291), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1329));
  AND2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(KEYINPUT61), .B1(new_n1324), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1321), .A2(new_n1323), .A3(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT61), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1333), .B1(new_n1322), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1320), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1322), .A2(KEYINPUT62), .A3(new_n1319), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1335), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT126), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1304), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1338), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT62), .B1(new_n1322), .B2(new_n1319), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1340), .B(new_n1331), .C1(new_n1342), .C2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1332), .B1(new_n1341), .B2(new_n1345), .ZN(G405));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1286), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1306), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1319), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1347), .B(new_n1306), .C1(new_n1317), .C2(new_n1318), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1304), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1304), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT127), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1351), .B1(new_n1352), .B2(new_n1353), .ZN(new_n1354));
  AOI211_X1 g1154(.A(KEYINPUT127), .B(new_n1304), .C1(new_n1349), .C2(new_n1350), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1354), .A2(new_n1355), .ZN(G402));
endmodule


