//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n467), .B1(new_n464), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT68), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n466), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n463), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n473), .A2(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n475), .A2(G136), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n464), .A2(new_n466), .A3(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(new_n462), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n482), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR3_X1   g073(.A1(new_n498), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n497), .A2(new_n499), .B1(new_n501), .B2(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n500), .A2(new_n503), .A3(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n494), .B1(new_n502), .B2(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(KEYINPUT70), .A2(G651), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT70), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  OAI21_X1  g086(.A(G543), .B1(new_n511), .B2(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT5), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G62), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(new_n518), .B1(G75), .B2(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(KEYINPUT72), .A3(G62), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n510), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT6), .B1(new_n507), .B2(new_n508), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n522), .A2(G543), .A3(new_n525), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n521), .A2(new_n530), .ZN(G166));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n523), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n534), .B2(new_n506), .ZN(new_n535));
  NOR3_X1   g110(.A1(new_n535), .A2(new_n514), .A3(new_n524), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n536), .A2(G51), .B1(new_n516), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n526), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(KEYINPUT73), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(G168));
  NAND2_X1  g121(.A1(new_n512), .A2(new_n515), .ZN(new_n547));
  NOR3_X1   g122(.A1(new_n535), .A2(new_n547), .A3(new_n524), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G90), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G64), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(new_n509), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n536), .A2(G52), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n549), .A2(new_n553), .A3(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  AOI22_X1  g131(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n510), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT74), .B(G43), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n536), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n548), .A2(G81), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  AND3_X1   g139(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G36), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n565), .A2(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n547), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n523), .B1(new_n572), .B2(KEYINPUT75), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n573), .B1(KEYINPUT75), .B2(new_n572), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n522), .A2(G53), .A3(G543), .A4(new_n525), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n548), .A2(G91), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  INV_X1    g154(.A(G166), .ZN(G303));
  INV_X1    g155(.A(G74), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n523), .B1(new_n547), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n548), .A2(G87), .B1(new_n536), .B2(G49), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n547), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(new_n509), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n522), .A2(G48), .A3(G543), .A4(new_n525), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n516), .A2(new_n522), .A3(G86), .A4(new_n525), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT77), .ZN(G305));
  NAND2_X1  g169(.A1(new_n536), .A2(G47), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT78), .B(G85), .Z(new_n596));
  AOI22_X1  g171(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n595), .B1(new_n526), .B2(new_n596), .C1(new_n510), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n548), .A2(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n528), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n522), .A2(KEYINPUT79), .A3(G543), .A4(new_n525), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n604), .A2(G54), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n547), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n606), .A2(KEYINPUT80), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(KEYINPUT80), .B1(new_n606), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n602), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT81), .Z(new_n614));
  OAI21_X1  g189(.A(new_n599), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n599), .B1(new_n614), .B2(G868), .ZN(G321));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NAND2_X1  g192(.A1(G299), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G168), .B2(new_n617), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(G168), .B2(new_n617), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n614), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n614), .A2(new_n621), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n624), .A2(KEYINPUT82), .A3(new_n617), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT82), .B1(new_n624), .B2(new_n617), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n625), .B(new_n626), .C1(G868), .C2(new_n563), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n497), .A2(new_n477), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT13), .Z(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n475), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n483), .A2(G123), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n462), .A2(KEYINPUT83), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT83), .B1(new_n462), .B2(G111), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G2104), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT84), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT16), .B(G1341), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(G14), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n649), .B2(new_n655), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2067), .B(G2678), .Z(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(G2072), .A2(G2078), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n442), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(KEYINPUT17), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n661), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n664), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n668), .B1(KEYINPUT85), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(KEYINPUT85), .B2(new_n670), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT87), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1981), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n688), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n686), .A2(new_n689), .A3(new_n693), .ZN(new_n695));
  NAND4_X1  g270(.A1(new_n691), .A2(new_n692), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n683), .B(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G6), .B(G305), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G16), .A2(G23), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n582), .B(KEYINPUT76), .ZN(new_n703));
  INV_X1    g278(.A(G87), .ZN(new_n704));
  INV_X1    g279(.A(G49), .ZN(new_n705));
  OAI22_X1  g280(.A1(new_n526), .A2(new_n704), .B1(new_n528), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n702), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n584), .A2(KEYINPUT91), .A3(new_n585), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n701), .B1(new_n709), .B2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT92), .B(G1976), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT33), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n700), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G22), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G166), .B2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1971), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n698), .A2(new_n699), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n710), .A2(new_n712), .ZN(new_n720));
  NOR4_X1   g295(.A1(new_n714), .A2(new_n718), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT34), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n715), .A2(G24), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G290), .B2(G16), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  OAI21_X1  g302(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n728));
  INV_X1    g303(.A(G107), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(G2105), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT90), .ZN(new_n731));
  AOI22_X1  g306(.A1(G131), .A2(new_n475), .B1(new_n483), .B2(G119), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(KEYINPUT89), .A2(G29), .ZN(new_n734));
  NOR2_X1   g309(.A1(KEYINPUT89), .A2(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G25), .B(new_n733), .S(new_n736), .Z(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT35), .B(G1991), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n737), .B(new_n738), .Z(new_n739));
  NAND4_X1  g314(.A1(new_n722), .A2(new_n726), .A3(new_n727), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT36), .ZN(new_n741));
  NAND2_X1  g316(.A1(G168), .A2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT100), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G16), .B2(G21), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1966), .ZN(new_n745));
  NAND2_X1  g320(.A1(G171), .A2(G16), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G5), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n736), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n640), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G28), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n752), .A2(KEYINPUT30), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(KEYINPUT30), .ZN(new_n754));
  OR2_X1    g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n745), .A2(new_n749), .A3(new_n751), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT101), .ZN(new_n759));
  NOR2_X1   g334(.A1(G4), .A2(G16), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n614), .B2(G16), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n747), .A2(new_n748), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n750), .A2(G35), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G162), .B2(new_n750), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT102), .B(KEYINPUT29), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n769));
  AND3_X1   g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n477), .A2(G105), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI211_X1 g349(.A(new_n771), .B(new_n774), .C1(G141), .C2(new_n475), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n483), .A2(G129), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  AND2_X1   g352(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G29), .B2(G32), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n764), .B1(G2090), .B2(new_n768), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n475), .A2(G140), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n483), .A2(G128), .ZN(new_n784));
  OR2_X1    g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n783), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n787), .A2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT94), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n750), .A2(G26), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT28), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G2067), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n715), .A2(G19), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT93), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n562), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1341), .Z(new_n797));
  NOR3_X1   g372(.A1(new_n782), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n750), .A2(G27), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G164), .B2(new_n750), .ZN(new_n800));
  INV_X1    g375(.A(G2078), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G160), .A2(G29), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n750), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT96), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n798), .B(new_n802), .C1(G2084), .C2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G29), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G33), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n475), .A2(G139), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n477), .A2(G103), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT25), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(KEYINPUT25), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n497), .A2(G127), .ZN(new_n818));
  INV_X1    g393(.A(G115), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n463), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n820), .B2(G2105), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(new_n811), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2072), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n780), .B2(new_n781), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n809), .A2(G2084), .ZN(new_n825));
  AOI21_X1  g400(.A(KEYINPUT99), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n810), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT23), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n828), .A2(new_n715), .A3(G20), .ZN(new_n829));
  NAND2_X1  g404(.A1(G299), .A2(G16), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n828), .B1(new_n715), .B2(G20), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT103), .B(G1956), .Z(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n768), .A2(G2090), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n833), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT104), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n824), .A2(KEYINPUT99), .A3(new_n825), .ZN(new_n839));
  AND4_X1   g414(.A1(new_n763), .A2(new_n827), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n741), .A2(new_n759), .A3(new_n840), .ZN(G150));
  INV_X1    g416(.A(G150), .ZN(G311));
  NAND2_X1  g417(.A1(new_n614), .A2(G559), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n548), .A2(G93), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT105), .B(G55), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n536), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n510), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n563), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n851), .A2(new_n562), .A3(new_n853), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n845), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n858), .B2(new_n845), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n499), .B1(new_n468), .B2(new_n469), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n504), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n494), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n787), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n778), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n821), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n630), .B(new_n733), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n475), .A2(G142), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n483), .A2(G130), .ZN(new_n875));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n873), .B(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G160), .B(new_n640), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n879), .B(KEYINPUT107), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n880), .B(new_n883), .C1(new_n884), .C2(new_n872), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n884), .B(new_n872), .Z(new_n886));
  OAI211_X1 g461(.A(new_n864), .B(new_n885), .C1(new_n886), .C2(new_n883), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g463(.A1(new_n854), .A2(new_n617), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n623), .B(new_n858), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n613), .B(G299), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT108), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n893), .B1(new_n890), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n709), .B(G290), .ZN(new_n902));
  XNOR2_X1  g477(.A(G305), .B(G166), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n901), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n889), .B1(new_n906), .B2(new_n617), .ZN(G295));
  OAI21_X1  g482(.A(new_n889), .B1(new_n906), .B2(new_n617), .ZN(G331));
  INV_X1    g483(.A(KEYINPUT112), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  INV_X1    g485(.A(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(new_n896), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n898), .B1(new_n912), .B2(new_n894), .ZN(new_n913));
  INV_X1    g488(.A(new_n899), .ZN(new_n914));
  OR2_X1    g489(.A1(G301), .A2(KEYINPUT109), .ZN(new_n915));
  NAND2_X1  g490(.A1(G168), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT110), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(G301), .B2(KEYINPUT109), .ZN(new_n918));
  AND3_X1   g493(.A1(G301), .A2(KEYINPUT109), .A3(new_n917), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n918), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(G168), .A3(new_n915), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n857), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n920), .A2(new_n855), .A3(new_n922), .A4(new_n856), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n913), .A2(new_n914), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT111), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n927), .A3(new_n925), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n923), .A2(new_n857), .A3(KEYINPUT111), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n891), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n911), .B1(new_n926), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n925), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(new_n897), .B2(new_n899), .ZN(new_n933));
  INV_X1    g508(.A(new_n930), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(new_n934), .A3(new_n904), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n864), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(new_n929), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n912), .A2(new_n894), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n939), .A2(new_n940), .B1(new_n891), .B2(new_n932), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n941), .B2(new_n911), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .A3(new_n935), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n910), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n937), .A3(new_n935), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n910), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n909), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT44), .B1(new_n946), .B2(new_n947), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n944), .A2(new_n951), .A3(KEYINPUT112), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G8), .ZN(new_n954));
  INV_X1    g529(.A(G1971), .ZN(new_n955));
  INV_X1    g530(.A(G40), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n473), .A2(new_n956), .A3(new_n479), .ZN(new_n957));
  AOI21_X1  g532(.A(G1384), .B1(new_n867), .B2(new_n868), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n958), .B2(KEYINPUT45), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n960));
  AOI211_X1 g535(.A(new_n960), .B(G1384), .C1(new_n867), .C2(new_n868), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n955), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G2090), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n965), .A3(new_n966), .A4(new_n957), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n954), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT119), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(G166), .B2(new_n954), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT55), .B(G8), .C1(new_n521), .C2(new_n530), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n968), .A2(new_n969), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1976), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n707), .B2(new_n708), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n957), .A2(new_n958), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G8), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n703), .A2(new_n702), .A3(new_n706), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT91), .B1(new_n584), .B2(new_n585), .ZN(new_n981));
  OAI21_X1  g556(.A(G1976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(G288), .B2(new_n975), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n548), .A2(G86), .B1(new_n589), .B2(new_n509), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n591), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n590), .A2(new_n988), .A3(new_n591), .A4(new_n592), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT117), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n593), .B2(G1981), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n593), .A2(new_n993), .A3(G1981), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n992), .B(KEYINPUT49), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n984), .ZN(new_n998));
  INV_X1    g573(.A(new_n994), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n995), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT49), .B1(new_n1000), .B2(new_n992), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n979), .B(new_n985), .C1(new_n998), .C2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n974), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n962), .A2(new_n967), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(G8), .A3(new_n973), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n968), .A2(KEYINPUT116), .A3(new_n973), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n969), .B1(new_n968), .B2(new_n973), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n957), .B1(new_n958), .B2(new_n964), .ZN(new_n1011));
  NOR3_X1   g586(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n1011), .A2(new_n1012), .A3(G2084), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n476), .A2(new_n478), .ZN(new_n1014));
  INV_X1    g589(.A(new_n472), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n497), .B2(G125), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1014), .B(G40), .C1(new_n1016), .C2(new_n462), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n869), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1019), .B2(new_n960), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1966), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G8), .B1(new_n1013), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(G286), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1003), .A2(new_n1009), .A3(new_n1010), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT63), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NOR4_X1   g602(.A1(new_n1002), .A2(new_n1023), .A3(new_n1026), .A4(G286), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n1009), .C1(new_n973), .C2(new_n968), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G299), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n574), .A2(new_n576), .A3(new_n577), .A4(new_n1031), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1956), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n960), .B1(G164), .B2(G1384), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT56), .B(G2072), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1038), .A2(new_n1021), .A3(new_n957), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1035), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2067), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n957), .A2(new_n958), .A3(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT121), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n762), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n613), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1037), .A2(new_n1035), .A3(new_n1040), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1041), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT61), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1037), .A2(new_n1035), .A3(new_n1040), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n1041), .ZN(new_n1052));
  INV_X1    g627(.A(new_n613), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1046), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT60), .B(new_n1053), .C1(new_n1044), .C2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n613), .B(KEYINPUT60), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1045), .A2(new_n1056), .A3(new_n1046), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1035), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1017), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1956), .B1(new_n1060), .B2(new_n965), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1039), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n959), .A2(new_n961), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1059), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(KEYINPUT61), .A3(new_n1048), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n1066));
  INV_X1    g641(.A(G1996), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1020), .A2(new_n1067), .A3(new_n1021), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n977), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1066), .B1(new_n1071), .B2(new_n563), .ZN(new_n1072));
  AOI211_X1 g647(.A(KEYINPUT59), .B(new_n562), .C1(new_n1068), .C2(new_n1070), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1065), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1049), .B1(new_n1058), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1038), .A2(new_n1021), .A3(new_n801), .A4(new_n957), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1020), .A2(KEYINPUT53), .A3(new_n801), .A4(new_n1021), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n748), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1078), .A2(new_n1079), .A3(G301), .A4(new_n1080), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1084));
  AND3_X1   g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1082), .A2(new_n1083), .B1(new_n1086), .B2(KEYINPUT54), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1023), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  NAND3_X1  g666(.A1(G286), .A2(new_n1091), .A3(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT122), .B1(G168), .B2(new_n954), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1089), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1096));
  INV_X1    g671(.A(G2084), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1966), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n959), .B2(new_n961), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1098), .A2(new_n1100), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1094), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1023), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1095), .B1(new_n1103), .B2(new_n1089), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1002), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1004), .A2(G8), .ZN(new_n1106));
  INV_X1    g681(.A(new_n973), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(KEYINPUT119), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1108), .A3(new_n1010), .ZN(new_n1109));
  AND4_X1   g684(.A1(KEYINPUT116), .A2(new_n1004), .A3(G8), .A4(new_n973), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT116), .B1(new_n968), .B2(new_n973), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1075), .A2(new_n1088), .A3(new_n1104), .A4(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(G288), .A2(G1976), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n998), .B2(new_n1001), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n978), .B1(new_n1116), .B2(new_n992), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1112), .B2(new_n1105), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1030), .A2(new_n1114), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1082), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1113), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT125), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1109), .A2(new_n1112), .A3(new_n1082), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1126), .B(new_n1127), .C1(KEYINPUT62), .C2(new_n1104), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1030), .A2(new_n1114), .A3(KEYINPUT124), .A4(new_n1118), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1121), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n787), .B(new_n1042), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT113), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1038), .A2(new_n1017), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1136), .A2(KEYINPUT114), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n778), .B(new_n1067), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1137), .B(new_n1138), .C1(new_n1135), .C2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n733), .A2(new_n738), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n733), .A2(new_n738), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1135), .ZN(new_n1144));
  XNOR2_X1  g719(.A(G290), .B(new_n725), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1140), .B(new_n1143), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT115), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1132), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n778), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1134), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT46), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1135), .A2(new_n1067), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1150), .A2(new_n1135), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT47), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1144), .A2(G1986), .A3(G290), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT48), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1155), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n787), .A2(G2067), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1160), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1144), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1148), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1148), .A2(KEYINPUT127), .A3(new_n1165), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g745(.A1(new_n675), .A2(G319), .ZN(new_n1172));
  NOR3_X1   g746(.A1(new_n1172), .A2(G401), .A3(G229), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n887), .A3(new_n1173), .ZN(G225));
  INV_X1    g748(.A(G225), .ZN(G308));
endmodule


