

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730;

  XNOR2_X1 U367 ( .A(n346), .B(n345), .ZN(G51) );
  NOR2_X1 U368 ( .A1(n665), .A2(n703), .ZN(n666) );
  INV_X1 U369 ( .A(n678), .ZN(n345) );
  NOR2_X1 U370 ( .A1(n354), .A2(n620), .ZN(n621) );
  BUF_X1 U371 ( .A(G101), .Z(n353) );
  XNOR2_X1 U372 ( .A(n555), .B(KEYINPUT42), .ZN(n729) );
  INV_X1 U373 ( .A(n471), .ZN(n349) );
  XNOR2_X1 U374 ( .A(n348), .B(n347), .ZN(n594) );
  XNOR2_X1 U375 ( .A(n545), .B(n544), .ZN(n654) );
  NOR2_X2 U376 ( .A1(n569), .A2(n543), .ZN(n348) );
  INV_X1 U377 ( .A(KEYINPUT39), .ZN(n347) );
  XNOR2_X1 U378 ( .A(n475), .B(KEYINPUT94), .ZN(n510) );
  NOR2_X1 U379 ( .A1(n559), .A2(n558), .ZN(n690) );
  BUF_X1 U380 ( .A(n539), .Z(n591) );
  XNOR2_X1 U381 ( .A(n369), .B(G469), .ZN(n553) );
  XNOR2_X1 U382 ( .A(n351), .B(n350), .ZN(n557) );
  NOR2_X1 U383 ( .A1(n625), .A2(n476), .ZN(n623) );
  INV_X1 U384 ( .A(KEYINPUT19), .ZN(n350) );
  OR2_X1 U385 ( .A1(n675), .A2(n600), .ZN(n425) );
  XNOR2_X1 U386 ( .A(n371), .B(n389), .ZN(n715) );
  XNOR2_X1 U387 ( .A(n352), .B(n413), .ZN(n420) );
  XNOR2_X1 U388 ( .A(n414), .B(n412), .ZN(n352) );
  XNOR2_X1 U389 ( .A(n365), .B(G104), .ZN(n409) );
  XNOR2_X1 U390 ( .A(G110), .B(G107), .ZN(n365) );
  XNOR2_X1 U391 ( .A(G119), .B(G116), .ZN(n376) );
  INV_X1 U392 ( .A(G953), .ZN(n718) );
  NAND2_X1 U393 ( .A1(n677), .A2(n612), .ZN(n346) );
  NOR2_X1 U394 ( .A1(n729), .A2(n726), .ZN(n556) );
  XNOR2_X1 U395 ( .A(n661), .B(n349), .ZN(n489) );
  XNOR2_X2 U396 ( .A(n470), .B(n469), .ZN(n661) );
  NOR2_X2 U397 ( .A1(n539), .A2(n427), .ZN(n351) );
  NOR2_X1 U398 ( .A1(n510), .A2(n639), .ZN(n439) );
  NAND2_X1 U399 ( .A1(n602), .A2(n601), .ZN(n619) );
  NAND2_X1 U400 ( .A1(n599), .A2(n598), .ZN(n602) );
  AND2_X1 U401 ( .A1(n553), .A2(n623), .ZN(n508) );
  XNOR2_X1 U402 ( .A(n425), .B(n424), .ZN(n539) );
  BUF_X1 U403 ( .A(n486), .Z(n630) );
  XNOR2_X1 U404 ( .A(G134), .B(n414), .ZN(n460) );
  INV_X1 U405 ( .A(n717), .ZN(n598) );
  XNOR2_X1 U406 ( .A(n550), .B(n549), .ZN(n576) );
  XNOR2_X1 U407 ( .A(KEYINPUT20), .B(n398), .ZN(n402) );
  XNOR2_X1 U408 ( .A(n503), .B(KEYINPUT106), .ZN(n645) );
  XNOR2_X1 U409 ( .A(n460), .B(n362), .ZN(n371) );
  NAND2_X1 U410 ( .A1(n597), .A2(n596), .ZN(n717) );
  XNOR2_X1 U411 ( .A(n694), .B(n502), .ZN(n593) );
  INV_X1 U412 ( .A(KEYINPUT105), .ZN(n502) );
  AND2_X1 U413 ( .A1(n536), .A2(n547), .ZN(n537) );
  NAND2_X1 U414 ( .A1(n576), .A2(n630), .ZN(n552) );
  XNOR2_X1 U415 ( .A(n484), .B(KEYINPUT32), .ZN(n618) );
  XNOR2_X1 U416 ( .A(n611), .B(n360), .ZN(n613) );
  XNOR2_X1 U417 ( .A(n605), .B(n356), .ZN(n607) );
  XOR2_X1 U418 ( .A(KEYINPUT78), .B(n619), .Z(n354) );
  XOR2_X1 U419 ( .A(KEYINPUT103), .B(G122), .Z(n355) );
  XNOR2_X1 U420 ( .A(KEYINPUT124), .B(n604), .ZN(n356) );
  XOR2_X1 U421 ( .A(KEYINPUT104), .B(KEYINPUT102), .Z(n357) );
  XNOR2_X1 U422 ( .A(n438), .B(KEYINPUT34), .ZN(n358) );
  XOR2_X1 U423 ( .A(n675), .B(n674), .Z(n359) );
  XOR2_X1 U424 ( .A(n610), .B(n609), .Z(n360) );
  AND2_X1 U425 ( .A1(n618), .A2(n616), .ZN(n361) );
  INV_X1 U426 ( .A(KEYINPUT65), .ZN(n471) );
  AND2_X1 U427 ( .A1(n571), .A2(n570), .ZN(n580) );
  XNOR2_X1 U428 ( .A(G902), .B(KEYINPUT89), .ZN(n397) );
  XNOR2_X1 U429 ( .A(KEYINPUT4), .B(G131), .ZN(n362) );
  INV_X1 U430 ( .A(KEYINPUT68), .ZN(n549) );
  XNOR2_X1 U431 ( .A(KEYINPUT48), .B(KEYINPUT85), .ZN(n586) );
  BUF_X1 U432 ( .A(n672), .Z(n699) );
  INV_X1 U433 ( .A(n567), .ZN(n466) );
  OR2_X1 U434 ( .A1(n475), .A2(n479), .ZN(n482) );
  INV_X1 U435 ( .A(n703), .ZN(n612) );
  XNOR2_X2 U436 ( .A(G143), .B(G128), .ZN(n414) );
  XNOR2_X1 U437 ( .A(G137), .B(KEYINPUT66), .ZN(n389) );
  XOR2_X1 U438 ( .A(G140), .B(KEYINPUT73), .Z(n364) );
  NAND2_X1 U439 ( .A1(G227), .A2(n718), .ZN(n363) );
  XNOR2_X1 U440 ( .A(n364), .B(n363), .ZN(n366) );
  XNOR2_X1 U441 ( .A(n366), .B(n409), .ZN(n367) );
  XNOR2_X1 U442 ( .A(KEYINPUT64), .B(G101), .ZN(n413) );
  XNOR2_X1 U443 ( .A(n413), .B(G146), .ZN(n370) );
  XNOR2_X1 U444 ( .A(n367), .B(n370), .ZN(n368) );
  XNOR2_X1 U445 ( .A(n715), .B(n368), .ZN(n668) );
  INV_X1 U446 ( .A(G902), .ZN(n450) );
  NAND2_X1 U447 ( .A1(n668), .A2(n450), .ZN(n369) );
  XNOR2_X1 U448 ( .A(n553), .B(KEYINPUT1), .ZN(n485) );
  XOR2_X1 U449 ( .A(n371), .B(n370), .Z(n381) );
  XOR2_X1 U450 ( .A(KEYINPUT5), .B(KEYINPUT72), .Z(n373) );
  XNOR2_X1 U451 ( .A(G137), .B(KEYINPUT97), .ZN(n372) );
  XNOR2_X1 U452 ( .A(n373), .B(n372), .ZN(n375) );
  NOR2_X1 U453 ( .A1(G953), .A2(G237), .ZN(n446) );
  NAND2_X1 U454 ( .A1(n446), .A2(G210), .ZN(n374) );
  XNOR2_X1 U455 ( .A(n375), .B(n374), .ZN(n379) );
  XNOR2_X1 U456 ( .A(n376), .B(KEYINPUT3), .ZN(n378) );
  XNOR2_X1 U457 ( .A(G113), .B(KEYINPUT90), .ZN(n377) );
  XNOR2_X1 U458 ( .A(n378), .B(n377), .ZN(n411) );
  XNOR2_X1 U459 ( .A(n379), .B(n411), .ZN(n380) );
  XNOR2_X1 U460 ( .A(n381), .B(n380), .ZN(n610) );
  NAND2_X1 U461 ( .A1(n610), .A2(n450), .ZN(n382) );
  XNOR2_X1 U462 ( .A(n382), .B(G472), .ZN(n486) );
  XNOR2_X1 U463 ( .A(n486), .B(KEYINPUT6), .ZN(n573) );
  NAND2_X1 U464 ( .A1(n718), .A2(G234), .ZN(n384) );
  XNOR2_X1 U465 ( .A(KEYINPUT81), .B(KEYINPUT8), .ZN(n383) );
  XNOR2_X1 U466 ( .A(n384), .B(n383), .ZN(n459) );
  NAND2_X1 U467 ( .A1(G221), .A2(n459), .ZN(n388) );
  XOR2_X1 U468 ( .A(KEYINPUT24), .B(G110), .Z(n386) );
  XNOR2_X1 U469 ( .A(G119), .B(G128), .ZN(n385) );
  XNOR2_X1 U470 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U471 ( .A(n388), .B(n387), .Z(n395) );
  INV_X1 U472 ( .A(n389), .ZN(n390) );
  XOR2_X1 U473 ( .A(n390), .B(KEYINPUT23), .Z(n393) );
  XNOR2_X1 U474 ( .A(G125), .B(G146), .ZN(n418) );
  INV_X1 U475 ( .A(KEYINPUT10), .ZN(n391) );
  XNOR2_X1 U476 ( .A(n391), .B(G140), .ZN(n392) );
  XNOR2_X1 U477 ( .A(n418), .B(n392), .ZN(n716) );
  XNOR2_X1 U478 ( .A(n393), .B(n716), .ZN(n394) );
  XNOR2_X1 U479 ( .A(n395), .B(n394), .ZN(n604) );
  NAND2_X1 U480 ( .A1(n604), .A2(n450), .ZN(n401) );
  INV_X1 U481 ( .A(KEYINPUT15), .ZN(n396) );
  XNOR2_X1 U482 ( .A(n397), .B(n396), .ZN(n422) );
  NAND2_X1 U483 ( .A1(G234), .A2(n422), .ZN(n398) );
  NAND2_X1 U484 ( .A1(n402), .A2(G217), .ZN(n399) );
  XNOR2_X1 U485 ( .A(n399), .B(KEYINPUT25), .ZN(n400) );
  XNOR2_X2 U486 ( .A(n401), .B(n400), .ZN(n625) );
  NAND2_X1 U487 ( .A1(n402), .A2(G221), .ZN(n403) );
  XNOR2_X1 U488 ( .A(n403), .B(KEYINPUT21), .ZN(n626) );
  XOR2_X1 U489 ( .A(n626), .B(KEYINPUT95), .Z(n476) );
  INV_X1 U490 ( .A(n623), .ZN(n404) );
  NOR2_X1 U491 ( .A1(n573), .A2(n404), .ZN(n405) );
  NAND2_X1 U492 ( .A1(n485), .A2(n405), .ZN(n407) );
  INV_X1 U493 ( .A(KEYINPUT33), .ZN(n406) );
  XNOR2_X1 U494 ( .A(n407), .B(n406), .ZN(n639) );
  XNOR2_X1 U495 ( .A(KEYINPUT16), .B(G122), .ZN(n408) );
  XNOR2_X1 U496 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U497 ( .A(n411), .B(n410), .ZN(n704) );
  XNOR2_X1 U498 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n412) );
  NAND2_X1 U499 ( .A1(n718), .A2(G224), .ZN(n416) );
  XNOR2_X1 U500 ( .A(n416), .B(KEYINPUT4), .ZN(n417) );
  XNOR2_X1 U501 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U502 ( .A(n419), .B(n420), .ZN(n421) );
  XNOR2_X1 U503 ( .A(n704), .B(n421), .ZN(n675) );
  INV_X1 U504 ( .A(n422), .ZN(n600) );
  INV_X1 U505 ( .A(G237), .ZN(n423) );
  NAND2_X1 U506 ( .A1(n450), .A2(n423), .ZN(n426) );
  NAND2_X1 U507 ( .A1(n426), .A2(G210), .ZN(n424) );
  NAND2_X1 U508 ( .A1(n426), .A2(G214), .ZN(n640) );
  INV_X1 U509 ( .A(n640), .ZN(n427) );
  XOR2_X1 U510 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n430) );
  NAND2_X1 U511 ( .A1(G234), .A2(G237), .ZN(n429) );
  XNOR2_X1 U512 ( .A(n430), .B(n429), .ZN(n433) );
  NAND2_X1 U513 ( .A1(n433), .A2(G952), .ZN(n431) );
  XOR2_X1 U514 ( .A(KEYINPUT91), .B(n431), .Z(n652) );
  NOR2_X1 U515 ( .A1(n652), .A2(G953), .ZN(n534) );
  INV_X1 U516 ( .A(n534), .ZN(n435) );
  XOR2_X1 U517 ( .A(G898), .B(KEYINPUT92), .Z(n710) );
  NAND2_X1 U518 ( .A1(n710), .A2(G953), .ZN(n432) );
  XOR2_X1 U519 ( .A(KEYINPUT93), .B(n432), .Z(n705) );
  NAND2_X1 U520 ( .A1(G902), .A2(n433), .ZN(n530) );
  OR2_X1 U521 ( .A1(n705), .A2(n530), .ZN(n434) );
  NAND2_X1 U522 ( .A1(n435), .A2(n434), .ZN(n436) );
  NAND2_X1 U523 ( .A1(n557), .A2(n436), .ZN(n437) );
  XNOR2_X2 U524 ( .A(n437), .B(KEYINPUT0), .ZN(n475) );
  INV_X1 U525 ( .A(KEYINPUT75), .ZN(n438) );
  XNOR2_X1 U526 ( .A(n439), .B(n358), .ZN(n467) );
  XOR2_X1 U527 ( .A(G104), .B(G122), .Z(n441) );
  XNOR2_X1 U528 ( .A(G113), .B(G143), .ZN(n440) );
  XNOR2_X1 U529 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U530 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n443) );
  XNOR2_X1 U531 ( .A(G131), .B(KEYINPUT11), .ZN(n442) );
  XNOR2_X1 U532 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U533 ( .A(n445), .B(n444), .Z(n449) );
  AND2_X1 U534 ( .A1(G214), .A2(n446), .ZN(n447) );
  XNOR2_X1 U535 ( .A(n716), .B(n447), .ZN(n448) );
  XNOR2_X1 U536 ( .A(n449), .B(n448), .ZN(n662) );
  NAND2_X1 U537 ( .A1(n662), .A2(n450), .ZN(n454) );
  XOR2_X1 U538 ( .A(KEYINPUT13), .B(KEYINPUT101), .Z(n452) );
  XNOR2_X1 U539 ( .A(KEYINPUT100), .B(G475), .ZN(n451) );
  XNOR2_X1 U540 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U541 ( .A(n454), .B(n453), .ZN(n499) );
  XNOR2_X1 U542 ( .A(G116), .B(G107), .ZN(n455) );
  XNOR2_X1 U543 ( .A(n355), .B(n455), .ZN(n458) );
  XNOR2_X1 U544 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n456) );
  XNOR2_X1 U545 ( .A(n357), .B(n456), .ZN(n457) );
  XOR2_X1 U546 ( .A(n458), .B(n457), .Z(n463) );
  NAND2_X1 U547 ( .A1(G217), .A2(n459), .ZN(n461) );
  XNOR2_X1 U548 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U549 ( .A(n463), .B(n462), .ZN(n701) );
  INV_X1 U550 ( .A(n701), .ZN(n464) );
  NAND2_X1 U551 ( .A1(n464), .A2(n450), .ZN(n465) );
  XNOR2_X1 U552 ( .A(G478), .B(n465), .ZN(n498) );
  INV_X1 U553 ( .A(n498), .ZN(n500) );
  OR2_X1 U554 ( .A1(n499), .A2(n500), .ZN(n567) );
  NAND2_X1 U555 ( .A1(n467), .A2(n466), .ZN(n470) );
  XNOR2_X1 U556 ( .A(KEYINPUT84), .B(KEYINPUT35), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n468), .B(KEYINPUT74), .ZN(n469) );
  XNOR2_X1 U558 ( .A(KEYINPUT88), .B(n485), .ZN(n578) );
  NAND2_X1 U559 ( .A1(n578), .A2(n573), .ZN(n473) );
  INV_X1 U560 ( .A(n625), .ZN(n546) );
  NOR2_X1 U561 ( .A1(n473), .A2(n546), .ZN(n474) );
  XNOR2_X1 U562 ( .A(n474), .B(KEYINPUT76), .ZN(n483) );
  NAND2_X1 U563 ( .A1(n499), .A2(n500), .ZN(n643) );
  NOR2_X1 U564 ( .A1(n476), .A2(n643), .ZN(n478) );
  INV_X1 U565 ( .A(KEYINPUT108), .ZN(n477) );
  XNOR2_X1 U566 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U567 ( .A(KEYINPUT70), .B(KEYINPUT22), .ZN(n480) );
  XNOR2_X1 U568 ( .A(n480), .B(KEYINPUT69), .ZN(n481) );
  XNOR2_X1 U569 ( .A(n482), .B(n481), .ZN(n517) );
  NAND2_X1 U570 ( .A1(n483), .A2(n517), .ZN(n484) );
  INV_X1 U571 ( .A(n485), .ZN(n505) );
  INV_X1 U572 ( .A(n505), .ZN(n622) );
  OR2_X1 U573 ( .A1(n630), .A2(n546), .ZN(n487) );
  NOR2_X1 U574 ( .A1(n622), .A2(n487), .ZN(n488) );
  NAND2_X1 U575 ( .A1(n517), .A2(n488), .ZN(n616) );
  NAND2_X1 U576 ( .A1(n489), .A2(n361), .ZN(n491) );
  INV_X1 U577 ( .A(KEYINPUT44), .ZN(n490) );
  NAND2_X1 U578 ( .A1(n491), .A2(n490), .ZN(n497) );
  NAND2_X1 U579 ( .A1(n661), .A2(KEYINPUT86), .ZN(n495) );
  AND2_X1 U580 ( .A1(n471), .A2(KEYINPUT44), .ZN(n492) );
  AND2_X1 U581 ( .A1(n616), .A2(n492), .ZN(n493) );
  AND2_X1 U582 ( .A1(n618), .A2(n493), .ZN(n494) );
  NAND2_X1 U583 ( .A1(n495), .A2(n494), .ZN(n496) );
  NAND2_X1 U584 ( .A1(n497), .A2(n496), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n498), .A2(n499), .ZN(n572) );
  INV_X1 U586 ( .A(n499), .ZN(n501) );
  NOR2_X4 U587 ( .A1(n501), .A2(n500), .ZN(n694) );
  NOR2_X1 U588 ( .A1(n572), .A2(n593), .ZN(n503) );
  XNOR2_X1 U589 ( .A(KEYINPUT80), .B(n645), .ZN(n565) );
  NAND2_X1 U590 ( .A1(n630), .A2(n623), .ZN(n504) );
  NOR2_X1 U591 ( .A1(n505), .A2(n504), .ZN(n635) );
  INV_X1 U592 ( .A(n475), .ZN(n506) );
  NAND2_X1 U593 ( .A1(n635), .A2(n506), .ZN(n507) );
  XNOR2_X1 U594 ( .A(n507), .B(KEYINPUT31), .ZN(n695) );
  XNOR2_X1 U595 ( .A(KEYINPUT96), .B(n508), .ZN(n536) );
  INV_X1 U596 ( .A(n630), .ZN(n509) );
  NAND2_X1 U597 ( .A1(n536), .A2(n509), .ZN(n511) );
  NOR2_X1 U598 ( .A1(n511), .A2(n510), .ZN(n512) );
  XNOR2_X1 U599 ( .A(n512), .B(KEYINPUT98), .ZN(n683) );
  NOR2_X1 U600 ( .A1(n695), .A2(n683), .ZN(n513) );
  NOR2_X1 U601 ( .A1(n565), .A2(n513), .ZN(n514) );
  XNOR2_X1 U602 ( .A(n514), .B(KEYINPUT107), .ZN(n519) );
  NAND2_X1 U603 ( .A1(n573), .A2(n546), .ZN(n515) );
  NOR2_X1 U604 ( .A1(n622), .A2(n515), .ZN(n516) );
  AND2_X1 U605 ( .A1(n517), .A2(n516), .ZN(n680) );
  INV_X1 U606 ( .A(n680), .ZN(n518) );
  NAND2_X1 U607 ( .A1(n519), .A2(n518), .ZN(n523) );
  NAND2_X1 U608 ( .A1(n661), .A2(KEYINPUT44), .ZN(n521) );
  INV_X1 U609 ( .A(KEYINPUT86), .ZN(n520) );
  AND2_X1 U610 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U611 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U612 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U613 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n526) );
  XNOR2_X1 U614 ( .A(n527), .B(n526), .ZN(n707) );
  INV_X1 U615 ( .A(n707), .ZN(n599) );
  NAND2_X1 U616 ( .A1(n630), .A2(n640), .ZN(n529) );
  XOR2_X1 U617 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n528) );
  XNOR2_X1 U618 ( .A(n529), .B(n528), .ZN(n538) );
  OR2_X1 U619 ( .A1(n718), .A2(n530), .ZN(n531) );
  XNOR2_X1 U620 ( .A(KEYINPUT110), .B(n531), .ZN(n532) );
  NOR2_X1 U621 ( .A1(G900), .A2(n532), .ZN(n533) );
  NOR2_X1 U622 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U623 ( .A(KEYINPUT77), .B(n535), .ZN(n547) );
  NAND2_X1 U624 ( .A1(n538), .A2(n537), .ZN(n569) );
  XOR2_X1 U625 ( .A(KEYINPUT38), .B(n591), .Z(n543) );
  NAND2_X1 U626 ( .A1(n572), .A2(n594), .ZN(n542) );
  XOR2_X1 U627 ( .A(KEYINPUT114), .B(KEYINPUT40), .Z(n541) );
  XNOR2_X1 U628 ( .A(n542), .B(n541), .ZN(n726) );
  INV_X1 U629 ( .A(n543), .ZN(n641) );
  NAND2_X1 U630 ( .A1(n641), .A2(n640), .ZN(n644) );
  NOR2_X1 U631 ( .A1(n644), .A2(n643), .ZN(n545) );
  XOR2_X1 U632 ( .A(KEYINPUT41), .B(KEYINPUT115), .Z(n544) );
  NOR2_X1 U633 ( .A1(n626), .A2(n546), .ZN(n548) );
  NAND2_X1 U634 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U635 ( .A(KEYINPUT28), .B(KEYINPUT113), .ZN(n551) );
  XNOR2_X1 U636 ( .A(n552), .B(n551), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n554), .A2(n553), .ZN(n559) );
  NOR2_X1 U638 ( .A1(n654), .A2(n559), .ZN(n555) );
  XNOR2_X1 U639 ( .A(KEYINPUT46), .B(n556), .ZN(n585) );
  INV_X1 U640 ( .A(n557), .ZN(n558) );
  INV_X1 U641 ( .A(n690), .ZN(n560) );
  NAND2_X1 U642 ( .A1(n560), .A2(KEYINPUT47), .ZN(n561) );
  XNOR2_X1 U643 ( .A(n561), .B(KEYINPUT79), .ZN(n562) );
  INV_X1 U644 ( .A(n562), .ZN(n564) );
  NAND2_X1 U645 ( .A1(n645), .A2(KEYINPUT47), .ZN(n563) );
  NAND2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n565), .A2(KEYINPUT47), .ZN(n566) );
  NAND2_X1 U648 ( .A1(n566), .A2(n690), .ZN(n571) );
  OR2_X1 U649 ( .A1(n567), .A2(n591), .ZN(n568) );
  NOR2_X1 U650 ( .A1(n569), .A2(n568), .ZN(n615) );
  INV_X1 U651 ( .A(n615), .ZN(n570) );
  XNOR2_X1 U652 ( .A(n572), .B(KEYINPUT109), .ZN(n681) );
  NOR2_X1 U653 ( .A1(n573), .A2(n681), .ZN(n574) );
  AND2_X1 U654 ( .A1(n574), .A2(n640), .ZN(n575) );
  NAND2_X1 U655 ( .A1(n576), .A2(n575), .ZN(n588) );
  NOR2_X1 U656 ( .A1(n588), .A2(n591), .ZN(n577) );
  XNOR2_X1 U657 ( .A(n577), .B(KEYINPUT36), .ZN(n579) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n698) );
  NAND2_X1 U659 ( .A1(n580), .A2(n698), .ZN(n581) );
  OR2_X2 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U661 ( .A(KEYINPUT67), .B(n583), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U663 ( .A(n587), .B(n586), .ZN(n597) );
  XOR2_X1 U664 ( .A(KEYINPUT111), .B(n588), .Z(n589) );
  NOR2_X1 U665 ( .A1(n622), .A2(n589), .ZN(n590) );
  XOR2_X1 U666 ( .A(n590), .B(KEYINPUT43), .Z(n592) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n617) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U669 ( .A(n595), .B(KEYINPUT116), .ZN(n727) );
  AND2_X1 U670 ( .A1(n617), .A2(n727), .ZN(n596) );
  INV_X1 U671 ( .A(KEYINPUT2), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n619), .A2(n600), .ZN(n603) );
  NOR2_X2 U673 ( .A1(n602), .A2(n601), .ZN(n620) );
  NOR2_X4 U674 ( .A1(n603), .A2(n620), .ZN(n672) );
  NAND2_X1 U675 ( .A1(n672), .A2(G217), .ZN(n605) );
  INV_X1 U676 ( .A(G952), .ZN(n606) );
  AND2_X1 U677 ( .A1(n606), .A2(G953), .ZN(n703) );
  NAND2_X1 U678 ( .A1(n607), .A2(n612), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U680 ( .A1(n672), .A2(G472), .ZN(n611) );
  XNOR2_X1 U681 ( .A(KEYINPUT117), .B(KEYINPUT62), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U683 ( .A(n614), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U684 ( .A(G143), .B(n615), .Z(G45) );
  XNOR2_X1 U685 ( .A(n616), .B(G110), .ZN(G12) );
  XNOR2_X1 U686 ( .A(n617), .B(G140), .ZN(G42) );
  XNOR2_X1 U687 ( .A(n618), .B(G119), .ZN(G21) );
  XNOR2_X1 U688 ( .A(n621), .B(KEYINPUT82), .ZN(n659) );
  NOR2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U690 ( .A(KEYINPUT50), .B(n624), .ZN(n633) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U692 ( .A(n627), .B(KEYINPUT49), .ZN(n628) );
  XNOR2_X1 U693 ( .A(n628), .B(KEYINPUT120), .ZN(n629) );
  NOR2_X1 U694 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U695 ( .A(KEYINPUT121), .B(n631), .ZN(n632) );
  NOR2_X1 U696 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U697 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U698 ( .A(KEYINPUT51), .B(n636), .Z(n637) );
  NOR2_X1 U699 ( .A1(n654), .A2(n637), .ZN(n638) );
  XNOR2_X1 U700 ( .A(n638), .B(KEYINPUT122), .ZN(n650) );
  NOR2_X1 U701 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U702 ( .A1(n643), .A2(n642), .ZN(n647) );
  NOR2_X1 U703 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U704 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U705 ( .A1(n639), .A2(n648), .ZN(n649) );
  NOR2_X1 U706 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U707 ( .A(n651), .B(KEYINPUT52), .ZN(n653) );
  OR2_X1 U708 ( .A1(n653), .A2(n652), .ZN(n657) );
  NOR2_X1 U709 ( .A1(n654), .A2(n639), .ZN(n655) );
  NOR2_X1 U710 ( .A1(n655), .A2(G953), .ZN(n656) );
  NAND2_X1 U711 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U712 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U713 ( .A(n660), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U714 ( .A(n661), .B(G122), .Z(G24) );
  NAND2_X1 U715 ( .A1(n672), .A2(G475), .ZN(n664) );
  XNOR2_X1 U716 ( .A(n662), .B(KEYINPUT59), .ZN(n663) );
  XNOR2_X1 U717 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U718 ( .A(n666), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U719 ( .A1(n699), .A2(G469), .ZN(n670) );
  XNOR2_X1 U720 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n667) );
  XNOR2_X1 U721 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U722 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U723 ( .A1(n671), .A2(n703), .ZN(G54) );
  NAND2_X1 U724 ( .A1(n672), .A2(G210), .ZN(n676) );
  XNOR2_X1 U725 ( .A(KEYINPUT87), .B(KEYINPUT54), .ZN(n673) );
  XNOR2_X1 U726 ( .A(n673), .B(KEYINPUT55), .ZN(n674) );
  XNOR2_X1 U727 ( .A(n676), .B(n359), .ZN(n677) );
  XOR2_X1 U728 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n678) );
  XOR2_X1 U729 ( .A(n353), .B(n680), .Z(G3) );
  INV_X1 U730 ( .A(n681), .ZN(n692) );
  NAND2_X1 U731 ( .A1(n683), .A2(n692), .ZN(n682) );
  XNOR2_X1 U732 ( .A(n682), .B(G104), .ZN(G6) );
  NAND2_X1 U733 ( .A1(n683), .A2(n694), .ZN(n684) );
  XNOR2_X1 U734 ( .A(n684), .B(KEYINPUT118), .ZN(n685) );
  XOR2_X1 U735 ( .A(n685), .B(KEYINPUT27), .Z(n687) );
  XNOR2_X1 U736 ( .A(G107), .B(KEYINPUT26), .ZN(n686) );
  XNOR2_X1 U737 ( .A(n687), .B(n686), .ZN(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n689) );
  NAND2_X1 U739 ( .A1(n690), .A2(n694), .ZN(n688) );
  XNOR2_X1 U740 ( .A(n689), .B(n688), .ZN(G30) );
  NAND2_X1 U741 ( .A1(n690), .A2(n692), .ZN(n691) );
  XNOR2_X1 U742 ( .A(n691), .B(G146), .ZN(G48) );
  NAND2_X1 U743 ( .A1(n695), .A2(n692), .ZN(n693) );
  XNOR2_X1 U744 ( .A(n693), .B(G113), .ZN(G15) );
  NAND2_X1 U745 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U746 ( .A(n696), .B(G116), .ZN(G18) );
  XOR2_X1 U747 ( .A(G125), .B(KEYINPUT37), .Z(n697) );
  XNOR2_X1 U748 ( .A(n698), .B(n697), .ZN(G27) );
  NAND2_X1 U749 ( .A1(n699), .A2(G478), .ZN(n700) );
  XNOR2_X1 U750 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U751 ( .A1(n703), .A2(n702), .ZN(G63) );
  XOR2_X1 U752 ( .A(n704), .B(n353), .Z(n706) );
  NAND2_X1 U753 ( .A1(n706), .A2(n705), .ZN(n714) );
  NOR2_X1 U754 ( .A1(n707), .A2(G953), .ZN(n712) );
  NAND2_X1 U755 ( .A1(G953), .A2(G224), .ZN(n708) );
  XOR2_X1 U756 ( .A(KEYINPUT61), .B(n708), .Z(n709) );
  NOR2_X1 U757 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U758 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U759 ( .A(n714), .B(n713), .ZN(G69) );
  XNOR2_X1 U760 ( .A(n716), .B(n715), .ZN(n720) );
  XNOR2_X1 U761 ( .A(n720), .B(n717), .ZN(n719) );
  NAND2_X1 U762 ( .A1(n719), .A2(n718), .ZN(n725) );
  XNOR2_X1 U763 ( .A(G227), .B(n720), .ZN(n721) );
  NAND2_X1 U764 ( .A1(n721), .A2(G900), .ZN(n722) );
  XNOR2_X1 U765 ( .A(KEYINPUT126), .B(n722), .ZN(n723) );
  NAND2_X1 U766 ( .A1(n723), .A2(G953), .ZN(n724) );
  NAND2_X1 U767 ( .A1(n725), .A2(n724), .ZN(G72) );
  XOR2_X1 U768 ( .A(n726), .B(G131), .Z(G33) );
  XOR2_X1 U769 ( .A(G134), .B(n727), .Z(n728) );
  XNOR2_X1 U770 ( .A(KEYINPUT119), .B(n728), .ZN(G36) );
  XNOR2_X1 U771 ( .A(G137), .B(KEYINPUT127), .ZN(n730) );
  XNOR2_X1 U772 ( .A(n730), .B(n729), .ZN(G39) );
endmodule

