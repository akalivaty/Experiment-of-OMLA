//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n201), .A2(new_n203), .A3(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n200), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n200), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n203), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n208), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT69), .B1(new_n199), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n196), .A2(new_n198), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n220));
  AOI21_X1  g034(.A(G143), .B1(new_n201), .B2(new_n203), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n215), .B1(new_n221), .B2(new_n210), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .A4(new_n208), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G116), .B(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT2), .A2(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT2), .A3(G113), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT2), .A2(G113), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n225), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(new_n231), .A3(new_n225), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT71), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n230), .A2(new_n231), .A3(new_n225), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n237), .B2(new_n232), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n192), .A2(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n194), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT66), .B1(new_n242), .B2(G131), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  AOI211_X1 g058(.A(new_n244), .B(new_n197), .C1(new_n241), .C2(new_n194), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n198), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT70), .B(new_n198), .C1(new_n243), .C2(new_n245), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n204), .A2(new_n206), .A3(new_n251), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT67), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT67), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n255), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n256), .B2(new_n213), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n248), .A2(new_n249), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n224), .A2(new_n240), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(G237), .A2(G953), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G210), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT27), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT72), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n237), .A2(new_n232), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n224), .B2(new_n258), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n222), .A2(new_n272), .A3(new_n208), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n219), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n257), .B(new_n198), .C1(new_n243), .C2(new_n245), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n274), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n268), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n259), .A2(new_n278), .A3(new_n264), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n266), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT31), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n266), .A2(new_n277), .A3(KEYINPUT31), .A4(new_n279), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n219), .A2(new_n222), .A3(new_n208), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n285), .A2(new_n235), .A3(new_n238), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT28), .B1(new_n286), .B2(new_n258), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n222), .A2(new_n272), .A3(new_n208), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n272), .B1(new_n222), .B2(new_n208), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n288), .A2(new_n289), .A3(new_n199), .ZN(new_n290));
  INV_X1    g104(.A(new_n257), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n246), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n268), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n259), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n287), .B1(new_n294), .B2(KEYINPUT28), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n295), .A2(new_n264), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G472), .A2(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n188), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  INV_X1    g115(.A(new_n264), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n277), .A2(new_n301), .A3(new_n259), .A4(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT75), .B(G902), .Z(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n285), .A2(new_n235), .A3(new_n238), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT64), .B(G146), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(G143), .ZN(new_n309));
  OAI22_X1  g123(.A1(new_n309), .A2(new_n255), .B1(new_n210), .B2(new_n221), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n246), .A2(new_n247), .B1(new_n310), .B2(new_n252), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n306), .B1(new_n249), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT74), .B1(new_n312), .B2(KEYINPUT28), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT74), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n287), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n224), .A2(new_n258), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n239), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n319), .B2(new_n259), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT29), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n302), .B1(new_n295), .B2(new_n301), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n305), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G472), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n296), .B1(new_n282), .B2(new_n283), .ZN(new_n325));
  INV_X1    g139(.A(new_n299), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT32), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n187), .B1(new_n300), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n329), .B1(new_n284), .B2(new_n297), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n322), .A2(new_n321), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n303), .A2(new_n304), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n324), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n188), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n325), .B2(new_n326), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(KEYINPUT76), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G217), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n304), .B2(G234), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(G902), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT23), .B1(new_n250), .B2(G119), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n250), .A2(G119), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OR2_X1    g160(.A1(KEYINPUT67), .A2(G128), .ZN(new_n347));
  NAND2_X1  g161(.A1(KEYINPUT67), .A2(G128), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n347), .A2(KEYINPUT23), .A3(G119), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT79), .B1(new_n350), .B2(G110), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n352));
  INV_X1    g166(.A(G110), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n346), .A2(new_n349), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT24), .B(G110), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(KEYINPUT77), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G119), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n253), .A2(new_n254), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n345), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n351), .B(new_n354), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT16), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G125), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(G125), .ZN(new_n367));
  INV_X1    g181(.A(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G140), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(G146), .B(new_n366), .C1(new_n370), .C2(new_n364), .ZN(new_n371));
  XNOR2_X1  g185(.A(G125), .B(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n308), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n363), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n366), .B1(new_n370), .B2(new_n364), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n200), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n371), .ZN(new_n377));
  INV_X1    g191(.A(new_n358), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(new_n362), .A3(new_n356), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n350), .B2(G110), .ZN(new_n381));
  AOI211_X1 g195(.A(KEYINPUT78), .B(new_n353), .C1(new_n346), .C2(new_n349), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n377), .B(new_n379), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G137), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(G221), .A3(G234), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n384), .B(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n374), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n374), .B2(new_n383), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT81), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n374), .A2(new_n383), .ZN(new_n393));
  INV_X1    g207(.A(new_n387), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n395), .A2(KEYINPUT81), .A3(new_n388), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n343), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT82), .ZN(new_n398));
  OR2_X1    g212(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n391), .B2(new_n304), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n304), .A3(new_n388), .A4(new_n399), .ZN(new_n401));
  NAND2_X1  g215(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n342), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(new_n343), .C1(new_n392), .C2(new_n396), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n398), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT85), .Z(new_n410));
  OAI21_X1  g224(.A(G210), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n360), .A2(G116), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n413), .B1(new_n414), .B2(KEYINPUT5), .ZN(new_n415));
  INV_X1    g229(.A(G116), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G119), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n417), .A3(KEYINPUT5), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(new_n360), .A3(KEYINPUT86), .A4(G116), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n415), .A2(new_n418), .A3(G113), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n234), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT89), .ZN(new_n425));
  INV_X1    g239(.A(G104), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT3), .B1(new_n426), .B2(G107), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT3), .ZN(new_n428));
  INV_X1    g242(.A(G107), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(G104), .ZN(new_n430));
  INV_X1    g244(.A(G101), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n426), .A2(G107), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n427), .A2(new_n430), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n426), .A2(G107), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n429), .A2(G104), .ZN(new_n435));
  OAI21_X1  g249(.A(G101), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n421), .A2(new_n234), .A3(KEYINPUT88), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n424), .A2(new_n425), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT8), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n421), .A2(new_n234), .A3(KEYINPUT88), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT88), .B1(new_n421), .B2(new_n234), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n443), .A2(new_n444), .A3(new_n437), .ZN(new_n445));
  INV_X1    g259(.A(new_n422), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT89), .B1(new_n446), .B2(new_n438), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n440), .B(new_n442), .C1(new_n445), .C2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n438), .A2(new_n234), .A3(new_n421), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n427), .A2(new_n430), .A3(new_n432), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G101), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT4), .A3(new_n433), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n453), .A3(G101), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n441), .B(new_n449), .C1(new_n455), .C2(new_n267), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n310), .A2(new_n368), .A3(new_n252), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n217), .A2(G125), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n385), .A2(G224), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT87), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n457), .A2(new_n458), .A3(new_n463), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n448), .A2(new_n456), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n468));
  INV_X1    g282(.A(G902), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n459), .B(new_n461), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n449), .B1(new_n455), .B2(new_n267), .ZN(new_n472));
  INV_X1    g286(.A(new_n441), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n476), .A3(new_n473), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n468), .B1(new_n467), .B2(new_n469), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n412), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n467), .A2(new_n469), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT90), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(new_n411), .A3(new_n478), .A4(new_n470), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n410), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT9), .B(G234), .ZN(new_n486));
  OAI21_X1  g300(.A(G221), .B1(new_n486), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n304), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT10), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n205), .B1(new_n308), .B2(G143), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n250), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n252), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n492), .A2(new_n493), .A3(new_n438), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n492), .B2(new_n438), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n489), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n452), .A2(new_n222), .A3(new_n208), .A4(new_n454), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n437), .A2(new_n489), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n257), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n500), .A3(new_n199), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n496), .A2(new_n500), .A3(KEYINPUT84), .A4(new_n199), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n497), .A2(new_n499), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n492), .A2(new_n438), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT83), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n492), .A2(new_n438), .A3(new_n493), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n506), .B1(new_n510), .B2(new_n489), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n511), .A2(new_n199), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G110), .B(G140), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n385), .A2(G227), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n514), .B(new_n515), .Z(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n503), .B2(new_n504), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT12), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n508), .A2(new_n509), .B1(new_n291), .B2(new_n437), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(new_n199), .ZN(new_n521));
  OAI22_X1  g335(.A1(new_n494), .A2(new_n495), .B1(new_n257), .B2(new_n438), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(KEYINPUT12), .A3(new_n219), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  AOI211_X1 g339(.A(G469), .B(new_n488), .C1(new_n517), .C2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n516), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n505), .A2(new_n512), .A3(new_n527), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n503), .A2(new_n504), .B1(new_n521), .B2(new_n523), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n528), .B(G469), .C1(new_n527), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G469), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n469), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n485), .B(new_n487), .C1(new_n526), .C2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G475), .A2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n260), .A2(G143), .A3(G214), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G143), .B1(new_n260), .B2(G214), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT17), .B(G131), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n376), .A2(new_n541), .A3(new_n371), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT92), .ZN(new_n545));
  OAI21_X1  g359(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n546));
  INV_X1    g360(.A(new_n540), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(new_n197), .A3(new_n538), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n545), .B1(new_n549), .B2(KEYINPUT17), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n376), .A2(new_n541), .A3(KEYINPUT91), .A4(new_n371), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n546), .A2(new_n548), .A3(KEYINPUT92), .A4(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n544), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G113), .B(G122), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(new_n426), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n373), .B1(new_n200), .B2(new_n372), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT18), .B(G131), .C1(new_n539), .C2(new_n540), .ZN(new_n558));
  NAND2_X1  g372(.A1(KEYINPUT18), .A2(G131), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n547), .A2(new_n538), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n372), .B(KEYINPUT19), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n371), .B(new_n549), .C1(new_n564), .C2(new_n211), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n561), .ZN(new_n566));
  INV_X1    g380(.A(new_n556), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n537), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT20), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT94), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n562), .A2(new_n568), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n536), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT20), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT93), .B1(new_n569), .B2(new_n570), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n578), .A3(new_n570), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n572), .A2(new_n576), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n554), .A2(new_n561), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n567), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n582), .B2(new_n562), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G475), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G952), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G953), .ZN(new_n588));
  INV_X1    g402(.A(G234), .ZN(new_n589));
  INV_X1    g403(.A(G237), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI211_X1 g406(.A(new_n385), .B(new_n304), .C1(G234), .C2(G237), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT21), .B(G898), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n347), .A2(G143), .A3(new_n348), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n212), .A2(G128), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n190), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT13), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n596), .B(new_n597), .C1(new_n599), .C2(new_n190), .ZN(new_n602));
  INV_X1    g416(.A(G122), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT95), .B1(new_n603), .B2(G116), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n416), .A3(G122), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(G116), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n429), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n607), .A2(new_n429), .A3(new_n608), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n601), .B(new_n602), .C1(new_n609), .C2(new_n611), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n607), .A2(KEYINPUT14), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n607), .A2(KEYINPUT14), .B1(G116), .B2(new_n603), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n429), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n596), .A2(new_n190), .A3(new_n597), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n610), .B1(new_n617), .B2(new_n598), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n612), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n486), .A2(new_n341), .A3(G953), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT96), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n612), .B(new_n621), .C1(new_n615), .C2(new_n618), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n304), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT98), .A4(new_n304), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(G478), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT15), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(KEYINPUT97), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(KEYINPUT97), .B2(new_n631), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT99), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n625), .B2(new_n626), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n635), .A2(new_n636), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n633), .B1(new_n627), .B2(new_n628), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT99), .B1(new_n640), .B2(new_n637), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n595), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n586), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n535), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n340), .A2(new_n408), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G101), .ZN(G3));
  INV_X1    g460(.A(new_n487), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n511), .A2(new_n199), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n503), .B2(new_n504), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n525), .B1(new_n649), .B2(new_n527), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n531), .A3(new_n304), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT84), .B1(new_n511), .B2(new_n199), .ZN(new_n652));
  INV_X1    g466(.A(new_n504), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n524), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n654), .A2(new_n516), .B1(new_n518), .B2(new_n512), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n532), .B1(new_n655), .B2(G469), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n647), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n408), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n298), .A2(new_n299), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n325), .B2(new_n488), .ZN(new_n660));
  INV_X1    g474(.A(new_n595), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n485), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n488), .A2(new_n630), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n623), .A2(new_n624), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT33), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT33), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n625), .A2(new_n630), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(KEYINPUT100), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n674));
  INV_X1    g488(.A(new_n672), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n674), .B1(new_n670), .B2(new_n675), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n580), .A2(new_n585), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n663), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT34), .B(G104), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  NAND3_X1  g497(.A1(new_n584), .A2(KEYINPUT101), .A3(G475), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  INV_X1    g499(.A(G475), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n685), .B1(new_n583), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n576), .A2(new_n577), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(new_n571), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n639), .A2(new_n641), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n663), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT35), .B(G107), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NOR2_X1   g510(.A1(new_n394), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n393), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n343), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n404), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n586), .A2(new_n642), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n659), .A2(new_n660), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n535), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT37), .B(G110), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G12));
  NAND2_X1  g522(.A1(new_n657), .A2(new_n701), .ZN(new_n709));
  INV_X1    g523(.A(new_n593), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n591), .B1(new_n710), .B2(G900), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n711), .B(KEYINPUT103), .Z(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n690), .A2(new_n485), .A3(new_n691), .A4(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n340), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G128), .ZN(G30));
  XOR2_X1   g531(.A(new_n712), .B(KEYINPUT39), .Z(new_n718));
  NAND2_X1  g532(.A1(new_n657), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(KEYINPUT40), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n481), .A2(new_n484), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT38), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n319), .A2(new_n259), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n302), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n280), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(G472), .B1(new_n725), .B2(G902), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n338), .B(new_n726), .C1(new_n325), .C2(new_n329), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n691), .A2(new_n678), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n728), .A2(new_n410), .A3(new_n701), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n720), .A2(new_n722), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G143), .ZN(G45));
  NAND4_X1  g545(.A1(new_n677), .A2(new_n678), .A3(new_n701), .A4(new_n713), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n535), .A2(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n300), .A2(new_n330), .A3(new_n187), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT76), .B1(new_n336), .B2(new_n338), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT104), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n340), .A2(new_n738), .A3(new_n733), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  AOI21_X1  g555(.A(new_n407), .B1(new_n331), .B2(new_n339), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n680), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n488), .B1(new_n517), .B2(new_n525), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n647), .B1(new_n744), .B2(new_n531), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n744), .A2(new_n746), .A3(new_n531), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n505), .A2(new_n527), .A3(new_n524), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n527), .B1(new_n505), .B2(new_n512), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n304), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT105), .B1(new_n750), .B2(G469), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n745), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n753));
  INV_X1    g567(.A(new_n485), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n595), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n746), .B1(new_n744), .B2(new_n531), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n750), .A2(KEYINPUT105), .A3(G469), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(new_n745), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n753), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n743), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT41), .B(G113), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NOR2_X1   g578(.A1(new_n752), .A2(KEYINPUT106), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n759), .B1(new_n758), .B2(new_n745), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n742), .A3(new_n755), .A4(new_n693), .ZN(new_n768));
  XOR2_X1   g582(.A(KEYINPUT107), .B(G116), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n768), .B(new_n769), .ZN(G18));
  AOI21_X1  g584(.A(new_n702), .B1(new_n331), .B2(new_n339), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n485), .A3(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT108), .B(G119), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G21));
  OAI21_X1  g588(.A(new_n302), .B1(new_n316), .B2(new_n320), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n284), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n299), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n660), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(new_n407), .A3(new_n728), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n767), .A2(new_n755), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n660), .A3(new_n701), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n782), .A2(new_n679), .A3(new_n712), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n753), .A3(new_n485), .A4(new_n760), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  XNOR2_X1  g599(.A(new_n332), .B(KEYINPUT111), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n335), .B1(new_n659), .B2(new_n327), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n407), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n679), .A2(new_n712), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n530), .A2(KEYINPUT109), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n655), .A2(new_n791), .A3(G469), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n651), .A2(new_n790), .A3(new_n792), .A4(new_n533), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n721), .A2(new_n410), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n793), .A2(new_n487), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n788), .A2(KEYINPUT42), .A3(new_n789), .A4(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n340), .A2(new_n408), .A3(new_n789), .A4(new_n795), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT42), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n797), .A2(KEYINPUT110), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT110), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  NAND4_X1  g616(.A1(new_n742), .A2(new_n693), .A3(new_n713), .A4(new_n795), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G134), .ZN(G36));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n805));
  OAI211_X1 g619(.A(KEYINPUT112), .B(G469), .C1(new_n655), .C2(KEYINPUT45), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n655), .A2(KEYINPUT45), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n528), .B1(new_n527), .B2(new_n529), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT112), .B1(new_n811), .B2(G469), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n805), .B1(new_n808), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(G469), .B1(new_n655), .B2(KEYINPUT45), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT113), .A3(new_n807), .A4(new_n806), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n813), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n533), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT46), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n532), .A2(new_n820), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n822), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n823), .ZN(new_n825));
  AOI211_X1 g639(.A(KEYINPUT114), .B(new_n825), .C1(new_n813), .C2(new_n817), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n821), .B(new_n651), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT43), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n586), .A2(new_n828), .A3(new_n677), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n673), .A2(new_n676), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT43), .B1(new_n678), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n829), .A2(new_n703), .A3(new_n701), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT44), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n794), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n832), .A2(new_n836), .A3(new_n833), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n836), .B1(new_n832), .B2(new_n833), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n718), .A2(new_n487), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n827), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G137), .ZN(G39));
  INV_X1    g656(.A(new_n340), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n407), .A3(new_n789), .A4(new_n794), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT116), .Z(new_n845));
  INV_X1    g659(.A(KEYINPUT47), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n827), .A2(new_n846), .A3(new_n487), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n532), .B1(new_n813), .B2(new_n817), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n651), .B1(new_n848), .B2(KEYINPUT46), .ZN(new_n849));
  INV_X1    g663(.A(new_n824), .ZN(new_n850));
  INV_X1    g664(.A(new_n826), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT47), .B1(new_n852), .B2(new_n647), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n845), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(G140), .ZN(G42));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n728), .A2(new_n754), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n727), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n404), .A2(new_n700), .A3(new_n713), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT120), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n793), .A2(new_n487), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n340), .A2(new_n738), .A3(new_n733), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n738), .B1(new_n340), .B2(new_n733), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n784), .A2(new_n716), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n737), .B2(new_n739), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n784), .A2(new_n716), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT121), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n856), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(KEYINPUT121), .A3(new_n871), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(KEYINPUT52), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n768), .A2(new_n772), .A3(new_n780), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n678), .B1(new_n635), .B2(new_n638), .ZN(new_n879));
  AOI22_X1  g693(.A1(new_n663), .A2(new_n879), .B1(new_n704), .B2(new_n705), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n743), .B2(new_n761), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(new_n645), .B2(new_n681), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n645), .A2(new_n882), .A3(new_n681), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n640), .A2(new_n637), .A3(new_n712), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n794), .A2(new_n690), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n709), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n888), .A2(new_n340), .B1(new_n783), .B2(new_n795), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n878), .A2(new_n884), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n801), .A2(new_n803), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n867), .A2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n784), .A2(new_n895), .A3(new_n716), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(KEYINPUT52), .A3(new_n870), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n873), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT53), .B1(new_n899), .B2(new_n892), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT54), .B1(new_n893), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n892), .ZN(new_n902));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT54), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n891), .B(new_n890), .C1(new_n873), .C2(new_n876), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n902), .B(new_n903), .C1(new_n904), .C2(KEYINPUT53), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n753), .A2(new_n760), .ZN(new_n906));
  INV_X1    g720(.A(new_n794), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n829), .A2(new_n592), .A3(new_n831), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n788), .A3(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT48), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n727), .A2(new_n407), .A3(new_n591), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n680), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n777), .A2(new_n660), .A3(new_n408), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n767), .A2(new_n485), .A3(new_n914), .A4(new_n909), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n911), .A2(new_n588), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n908), .A2(new_n909), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n908), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n586), .A2(new_n830), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n782), .A2(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n909), .A2(new_n914), .ZN(new_n921));
  INV_X1    g735(.A(new_n410), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n921), .A2(new_n906), .A3(new_n922), .A4(new_n722), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n923), .A2(KEYINPUT50), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(KEYINPUT50), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n758), .A2(new_n651), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n487), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n853), .B2(new_n847), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n921), .A2(new_n907), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT123), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n926), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT51), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT51), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n934), .B(new_n926), .C1(new_n929), .C2(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n916), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n901), .A2(new_n905), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT124), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n901), .A2(new_n905), .A3(new_n936), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n587), .A2(new_n385), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n408), .A2(new_n487), .A3(new_n922), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n943), .A2(new_n678), .A3(new_n830), .ZN(new_n944));
  INV_X1    g758(.A(new_n927), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT49), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT117), .ZN(new_n948));
  AOI211_X1 g762(.A(new_n722), .B(new_n727), .C1(new_n945), .C2(new_n946), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n942), .A2(new_n950), .ZN(G75));
  NAND2_X1  g765(.A1(new_n877), .A2(new_n892), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT53), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n902), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n488), .A3(new_n412), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT56), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n475), .A2(new_n477), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n471), .ZN(new_n959));
  XNOR2_X1  g773(.A(KEYINPUT125), .B(KEYINPUT55), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n956), .A2(new_n957), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n956), .B2(new_n957), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n385), .A2(G952), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(G51));
  XNOR2_X1  g779(.A(new_n532), .B(KEYINPUT57), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n954), .A2(new_n903), .A3(new_n902), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n903), .B1(new_n954), .B2(new_n902), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n650), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n955), .A2(new_n488), .A3(new_n813), .A4(new_n817), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(G54));
  AND2_X1   g786(.A1(KEYINPUT58), .A2(G475), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n955), .A2(new_n488), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n562), .A3(new_n568), .ZN(new_n975));
  INV_X1    g789(.A(new_n964), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n955), .A2(new_n488), .A3(new_n573), .A4(new_n973), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(G60));
  NAND2_X1  g792(.A1(new_n668), .A2(new_n669), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT59), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n979), .B(new_n981), .C1(new_n967), .C2(new_n968), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n976), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n901), .A2(new_n905), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n979), .B1(new_n984), .B2(new_n981), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(G63));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT60), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n892), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT53), .B1(new_n877), .B2(new_n892), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n699), .B(new_n989), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n988), .B1(new_n954), .B2(new_n902), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n392), .A2(new_n396), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n992), .B(new_n976), .C1(new_n993), .C2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G66));
  NAND3_X1  g812(.A1(new_n878), .A2(new_n884), .A3(new_n885), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n385), .ZN(new_n1000));
  INV_X1    g814(.A(G224), .ZN(new_n1001));
  OAI21_X1  g815(.A(G953), .B1(new_n594), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n958), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(G898), .B2(new_n385), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1003), .B(new_n1005), .ZN(G69));
  AOI22_X1  g820(.A1(new_n894), .A2(new_n896), .B1(new_n739), .B2(new_n737), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n730), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1009));
  INV_X1    g823(.A(new_n841), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n794), .B1(new_n680), .B2(new_n879), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(new_n719), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1010), .B1(new_n742), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1009), .A2(new_n854), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n385), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n270), .A2(new_n276), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(new_n564), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n385), .B1(G227), .B2(G900), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1018), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n385), .A2(G900), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n827), .A2(new_n788), .A3(new_n840), .A4(new_n857), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n1023), .A2(new_n801), .A3(new_n803), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT126), .ZN(new_n1025));
  AND3_X1   g839(.A1(new_n1007), .A2(new_n1025), .A3(new_n841), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1025), .B1(new_n1007), .B2(new_n841), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1024), .B(new_n854), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1022), .B1(new_n1028), .B2(new_n385), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1021), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1023), .A2(new_n801), .A3(new_n803), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n852), .A2(KEYINPUT47), .A3(new_n647), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n846), .B1(new_n827), .B2(new_n487), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1032), .B1(new_n1035), .B2(new_n845), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1007), .A2(new_n841), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT126), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1007), .A2(new_n841), .A3(new_n1025), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(G953), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1041), .A2(KEYINPUT127), .A3(new_n1022), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1019), .B(new_n1020), .C1(new_n1031), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g857(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(KEYINPUT127), .B1(new_n1041), .B2(new_n1022), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1028), .A2(new_n385), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1022), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1046), .A2(new_n1030), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1045), .A2(new_n1021), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1020), .B1(new_n1049), .B2(new_n1019), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1044), .A2(new_n1050), .ZN(G72));
  NAND2_X1  g865(.A1(G472), .A2(G902), .ZN(new_n1052));
  XOR2_X1   g866(.A(new_n1052), .B(KEYINPUT63), .Z(new_n1053));
  OAI21_X1  g867(.A(new_n1053), .B1(new_n1015), .B2(new_n999), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n277), .A2(new_n259), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1054), .A2(new_n264), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1053), .B1(new_n1028), .B2(new_n999), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n1057), .A2(new_n259), .A3(new_n302), .A4(new_n277), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1055), .A2(new_n302), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1059), .A2(new_n280), .ZN(new_n1060));
  OAI211_X1 g874(.A(new_n1053), .B(new_n1060), .C1(new_n893), .C2(new_n900), .ZN(new_n1061));
  AND4_X1   g875(.A1(new_n976), .A2(new_n1056), .A3(new_n1058), .A4(new_n1061), .ZN(G57));
endmodule


