

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XNOR2_X1 U324 ( .A(KEYINPUT38), .B(n454), .ZN(n508) );
  XOR2_X1 U325 ( .A(n378), .B(n391), .Z(n526) );
  XNOR2_X1 U326 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U327 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n292) );
  INV_X1 U328 ( .A(KEYINPUT25), .ZN(n397) );
  XNOR2_X1 U329 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U330 ( .A(G176GAT), .B(G92GAT), .ZN(n365) );
  XNOR2_X1 U331 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U332 ( .A(n365), .B(G64GAT), .ZN(n440) );
  XNOR2_X1 U333 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U334 ( .A(n369), .B(n292), .ZN(n370) );
  XNOR2_X1 U335 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U336 ( .A1(n571), .A2(n414), .ZN(n416) );
  INV_X1 U337 ( .A(KEYINPUT106), .ZN(n455) );
  XNOR2_X1 U338 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n484) );
  XNOR2_X1 U339 ( .A(n455), .B(G36GAT), .ZN(n456) );
  XNOR2_X1 U340 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n457), .B(n456), .ZN(G1329GAT) );
  XOR2_X1 U342 ( .A(G64GAT), .B(G155GAT), .Z(n294) );
  XNOR2_X1 U343 ( .A(G127GAT), .B(G71GAT), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U345 ( .A(G57GAT), .B(KEYINPUT13), .Z(n443) );
  XOR2_X1 U346 ( .A(n295), .B(n443), .Z(n297) );
  XNOR2_X1 U347 ( .A(G183GAT), .B(G211GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n302) );
  XOR2_X1 U349 ( .A(G8GAT), .B(KEYINPUT79), .Z(n369) );
  XNOR2_X1 U350 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n298), .B(G15GAT), .ZN(n429) );
  XOR2_X1 U352 ( .A(n369), .B(n429), .Z(n300) );
  NAND2_X1 U353 ( .A1(G231GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U355 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n304) );
  XNOR2_X1 U357 ( .A(G22GAT), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U359 ( .A(KEYINPUT12), .B(KEYINPUT82), .Z(n306) );
  XNOR2_X1 U360 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n571) );
  XOR2_X1 U364 ( .A(G99GAT), .B(G85GAT), .Z(n444) );
  XOR2_X1 U365 ( .A(KEYINPUT10), .B(n444), .Z(n312) );
  XOR2_X1 U366 ( .A(G36GAT), .B(G190GAT), .Z(n366) );
  XNOR2_X1 U367 ( .A(G218GAT), .B(n366), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U369 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n314) );
  NAND2_X1 U370 ( .A1(G232GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U372 ( .A(n316), .B(n315), .Z(n318) );
  XOR2_X1 U373 ( .A(G134GAT), .B(KEYINPUT78), .Z(n337) );
  XNOR2_X1 U374 ( .A(n337), .B(G92GAT), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT68), .B(G106GAT), .Z(n320) );
  XNOR2_X1 U377 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n319) );
  XNOR2_X1 U378 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U379 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U380 ( .A(G29GAT), .B(G43GAT), .Z(n324) );
  XNOR2_X1 U381 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n323) );
  XNOR2_X1 U382 ( .A(n324), .B(n323), .ZN(n430) );
  XNOR2_X1 U383 ( .A(G50GAT), .B(G162GAT), .ZN(n325) );
  XNOR2_X1 U384 ( .A(n325), .B(KEYINPUT77), .ZN(n386) );
  XNOR2_X1 U385 ( .A(n430), .B(n386), .ZN(n326) );
  XNOR2_X1 U386 ( .A(n327), .B(n326), .ZN(n466) );
  XNOR2_X1 U387 ( .A(n466), .B(KEYINPUT36), .ZN(n590) );
  XOR2_X1 U388 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n329) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n347) );
  XOR2_X1 U391 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n331) );
  XNOR2_X1 U392 ( .A(G57GAT), .B(KEYINPUT5), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U394 ( .A(G148GAT), .B(G162GAT), .Z(n333) );
  XNOR2_X1 U395 ( .A(G29GAT), .B(G85GAT), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n345) );
  XNOR2_X1 U398 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n336) );
  XNOR2_X1 U399 ( .A(n336), .B(G127GAT), .ZN(n352) );
  XOR2_X1 U400 ( .A(n337), .B(n352), .Z(n339) );
  NAND2_X1 U401 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n341) );
  XNOR2_X1 U403 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n340), .B(KEYINPUT2), .ZN(n393) );
  XOR2_X1 U405 ( .A(n341), .B(n393), .Z(n343) );
  XNOR2_X1 U406 ( .A(G141GAT), .B(G120GAT), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n524) );
  INV_X1 U410 ( .A(n524), .ZN(n406) );
  XNOR2_X1 U411 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n348), .B(KEYINPUT18), .ZN(n349) );
  XOR2_X1 U413 ( .A(n349), .B(KEYINPUT17), .Z(n351) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n373) );
  XOR2_X1 U416 ( .A(G120GAT), .B(G71GAT), .Z(n447) );
  XOR2_X1 U417 ( .A(n447), .B(n352), .Z(n354) );
  XNOR2_X1 U418 ( .A(G99GAT), .B(G190GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U420 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n356) );
  NAND2_X1 U421 ( .A1(G227GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U423 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U424 ( .A(G176GAT), .B(G134GAT), .Z(n360) );
  XNOR2_X1 U425 ( .A(G43GAT), .B(G15GAT), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n361), .B(KEYINPUT84), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n373), .B(n364), .ZN(n538) );
  XOR2_X1 U430 ( .A(n366), .B(n440), .Z(n368) );
  NAND2_X1 U431 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U432 ( .A(n368), .B(n367), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U434 ( .A(KEYINPUT87), .B(G204GAT), .Z(n375) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(G211GAT), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U437 ( .A(G218GAT), .B(KEYINPUT21), .Z(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n391) );
  INV_X1 U439 ( .A(n526), .ZN(n473) );
  NAND2_X1 U440 ( .A1(n538), .A2(n473), .ZN(n379) );
  XOR2_X1 U441 ( .A(KEYINPUT99), .B(n379), .Z(n396) );
  XOR2_X1 U442 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XOR2_X1 U443 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT22), .B(KEYINPUT88), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U446 ( .A(n420), .B(n382), .Z(n384) );
  NAND2_X1 U447 ( .A1(G228GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U448 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U449 ( .A(n385), .B(KEYINPUT90), .Z(n388) );
  XNOR2_X1 U450 ( .A(n386), .B(KEYINPUT24), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n390) );
  XNOR2_X1 U452 ( .A(G148GAT), .B(G106GAT), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n389), .B(G78GAT), .ZN(n442) );
  XOR2_X1 U454 ( .A(n390), .B(n442), .Z(n395) );
  INV_X1 U455 ( .A(n391), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n479) );
  AND2_X1 U458 ( .A1(n396), .A2(n479), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n404) );
  XNOR2_X1 U460 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n399) );
  XNOR2_X1 U461 ( .A(n399), .B(n473), .ZN(n408) );
  NOR2_X1 U462 ( .A1(n479), .A2(n538), .ZN(n401) );
  XNOR2_X1 U463 ( .A(KEYINPUT98), .B(KEYINPUT26), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n575) );
  INV_X1 U465 ( .A(n575), .ZN(n402) );
  NOR2_X1 U466 ( .A1(n408), .A2(n402), .ZN(n403) );
  NOR2_X1 U467 ( .A1(n404), .A2(n403), .ZN(n405) );
  NOR2_X1 U468 ( .A1(n406), .A2(n405), .ZN(n407) );
  XOR2_X1 U469 ( .A(KEYINPUT100), .B(n407), .Z(n413) );
  NOR2_X1 U470 ( .A1(n524), .A2(n408), .ZN(n535) );
  XNOR2_X1 U471 ( .A(n479), .B(KEYINPUT28), .ZN(n540) );
  NAND2_X1 U472 ( .A1(n535), .A2(n540), .ZN(n409) );
  XNOR2_X1 U473 ( .A(KEYINPUT96), .B(n409), .ZN(n410) );
  NOR2_X1 U474 ( .A1(n538), .A2(n410), .ZN(n411) );
  XNOR2_X1 U475 ( .A(KEYINPUT97), .B(n411), .ZN(n412) );
  NAND2_X1 U476 ( .A1(n413), .A2(n412), .ZN(n490) );
  NAND2_X1 U477 ( .A1(n590), .A2(n490), .ZN(n414) );
  XNOR2_X1 U478 ( .A(KEYINPUT105), .B(KEYINPUT37), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n523) );
  XOR2_X1 U480 ( .A(G113GAT), .B(G50GAT), .Z(n418) );
  XNOR2_X1 U481 ( .A(G169GAT), .B(G36GAT), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U483 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U484 ( .A1(G229GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n434) );
  XOR2_X1 U486 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n424) );
  XNOR2_X1 U487 ( .A(KEYINPUT69), .B(KEYINPUT30), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U489 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n426) );
  XNOR2_X1 U490 ( .A(G197GAT), .B(G8GAT), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U492 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U495 ( .A(n434), .B(n433), .Z(n563) );
  INV_X1 U496 ( .A(n563), .ZN(n576) );
  XOR2_X1 U497 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n436) );
  XNOR2_X1 U498 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n453) );
  NAND2_X1 U500 ( .A1(G230GAT), .A2(G233GAT), .ZN(n438) );
  INV_X1 U501 ( .A(KEYINPUT76), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n445) );
  XNOR2_X1 U504 ( .A(n446), .B(n445), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n447), .B(G204GAT), .ZN(n449) );
  INV_X1 U506 ( .A(KEYINPUT74), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n463) );
  NOR2_X1 U508 ( .A1(n576), .A2(n463), .ZN(n491) );
  NAND2_X1 U509 ( .A1(n523), .A2(n491), .ZN(n454) );
  NOR2_X1 U510 ( .A1(n508), .A2(n526), .ZN(n457) );
  INV_X1 U511 ( .A(KEYINPUT64), .ZN(n478) );
  XNOR2_X1 U512 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n459) );
  NAND2_X1 U513 ( .A1(n571), .A2(n590), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U515 ( .A1(n463), .A2(n460), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n461), .A2(n576), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(KEYINPUT114), .ZN(n471) );
  INV_X1 U518 ( .A(KEYINPUT41), .ZN(n464) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n568) );
  NAND2_X1 U520 ( .A1(n568), .A2(n563), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT46), .ZN(n468) );
  INV_X1 U522 ( .A(n466), .ZN(n561) );
  INV_X1 U523 ( .A(n561), .ZN(n486) );
  NOR2_X1 U524 ( .A1(n486), .A2(n571), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U526 ( .A(n469), .B(KEYINPUT47), .Z(n470) );
  NAND2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT48), .ZN(n536) );
  NAND2_X1 U529 ( .A1(n536), .A2(n473), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n474) );
  XNOR2_X1 U531 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n476), .A2(n524), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n478), .B(n477), .ZN(n574) );
  NAND2_X1 U534 ( .A1(n574), .A2(n479), .ZN(n481) );
  XOR2_X1 U535 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n480) );
  XNOR2_X1 U536 ( .A(n481), .B(n480), .ZN(n482) );
  NAND2_X1 U537 ( .A1(n538), .A2(n482), .ZN(n483) );
  XOR2_X1 U538 ( .A(KEYINPUT122), .B(n483), .Z(n572) );
  NAND2_X1 U539 ( .A1(n572), .A2(n486), .ZN(n485) );
  INV_X1 U540 ( .A(n571), .ZN(n586) );
  NOR2_X1 U541 ( .A1(n586), .A2(n486), .ZN(n487) );
  XNOR2_X1 U542 ( .A(n487), .B(KEYINPUT16), .ZN(n488) );
  XOR2_X1 U543 ( .A(KEYINPUT83), .B(n488), .Z(n489) );
  AND2_X1 U544 ( .A1(n490), .A2(n489), .ZN(n510) );
  NAND2_X1 U545 ( .A1(n491), .A2(n510), .ZN(n492) );
  XOR2_X1 U546 ( .A(KEYINPUT101), .B(n492), .Z(n500) );
  NOR2_X1 U547 ( .A1(n524), .A2(n500), .ZN(n494) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U549 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n495), .Z(G1324GAT) );
  NOR2_X1 U551 ( .A1(n526), .A2(n500), .ZN(n496) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  INV_X1 U553 ( .A(n538), .ZN(n529) );
  NOR2_X1 U554 ( .A1(n529), .A2(n500), .ZN(n498) );
  XNOR2_X1 U555 ( .A(KEYINPUT35), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U557 ( .A(G15GAT), .B(n499), .Z(G1326GAT) );
  NOR2_X1 U558 ( .A1(n540), .A2(n500), .ZN(n501) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(n501), .Z(n502) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(n502), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n508), .A2(n524), .ZN(n503) );
  XNOR2_X1 U562 ( .A(n503), .B(KEYINPUT39), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(n504), .ZN(G1328GAT) );
  XNOR2_X1 U564 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n506) );
  NOR2_X1 U565 ( .A1(n529), .A2(n508), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U567 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NOR2_X1 U568 ( .A1(n508), .A2(n540), .ZN(n509) );
  XOR2_X1 U569 ( .A(G50GAT), .B(n509), .Z(G1331GAT) );
  INV_X1 U570 ( .A(n568), .ZN(n554) );
  NOR2_X1 U571 ( .A1(n563), .A2(n554), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n510), .A2(n522), .ZN(n517) );
  NOR2_X1 U573 ( .A1(n524), .A2(n517), .ZN(n511) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U575 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U576 ( .A1(n526), .A2(n517), .ZN(n514) );
  XNOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n529), .A2(n517), .ZN(n516) );
  XOR2_X1 U581 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U582 ( .A1(n517), .A2(n540), .ZN(n521) );
  XOR2_X1 U583 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n519) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(KEYINPUT111), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n522), .ZN(n532) );
  NOR2_X1 U588 ( .A1(n524), .A2(n532), .ZN(n525) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n526), .A2(n532), .ZN(n527) );
  XOR2_X1 U591 ( .A(KEYINPUT112), .B(n527), .Z(n528) );
  XNOR2_X1 U592 ( .A(G92GAT), .B(n528), .ZN(G1337GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n532), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1338GAT) );
  NOR2_X1 U596 ( .A1(n540), .A2(n532), .ZN(n533) );
  XOR2_X1 U597 ( .A(KEYINPUT44), .B(n533), .Z(n534) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U600 ( .A(KEYINPUT115), .B(n537), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n551), .A2(n538), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(n539), .Z(n541) );
  NAND2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n576), .A2(n548), .ZN(n543) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(KEYINPUT117), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  NOR2_X1 U607 ( .A1(n554), .A2(n548), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U610 ( .A1(n586), .A2(n548), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  NOR2_X1 U613 ( .A1(n561), .A2(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n551), .A2(n575), .ZN(n560) );
  NOR2_X1 U617 ( .A1(n576), .A2(n560), .ZN(n552) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n552), .Z(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT118), .B(n553), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n560), .A2(n554), .ZN(n558) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n586), .A2(n560), .ZN(n559) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n572), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n566) );
  XNOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT123), .B(n567), .Z(n570) );
  NAND2_X1 U635 ( .A1(n572), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n588) );
  NOR2_X1 U640 ( .A1(n576), .A2(n588), .ZN(n581) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(KEYINPUT59), .B(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  INV_X1 U646 ( .A(n463), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n582), .A2(n588), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n585), .Z(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n588), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  INV_X1 U653 ( .A(n588), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

