

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U551 ( .A(KEYINPUT66), .B(n535), .Z(n797) );
  XOR2_X1 U552 ( .A(G543), .B(KEYINPUT0), .Z(n575) );
  XNOR2_X1 U553 ( .A(n558), .B(KEYINPUT5), .ZN(n562) );
  NOR2_X1 U554 ( .A1(G651), .A2(n575), .ZN(n790) );
  NOR2_X1 U555 ( .A1(n527), .A2(n526), .ZN(G160) );
  XOR2_X1 U556 ( .A(KEYINPUT6), .B(n561), .Z(n516) );
  XNOR2_X1 U557 ( .A(KEYINPUT88), .B(KEYINPUT27), .ZN(n595) );
  XNOR2_X1 U558 ( .A(n596), .B(n595), .ZN(n598) );
  INV_X1 U559 ( .A(n656), .ZN(n638) );
  NOR2_X1 U560 ( .A1(n654), .A2(n653), .ZN(n667) );
  XNOR2_X1 U561 ( .A(KEYINPUT92), .B(KEYINPUT32), .ZN(n664) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n796) );
  AND2_X1 U563 ( .A1(n562), .A2(n516), .ZN(n563) );
  XNOR2_X1 U564 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X1 U566 ( .A(KEYINPUT17), .B(n517), .Z(n528) );
  NAND2_X1 U567 ( .A1(G137), .A2(n528), .ZN(n519) );
  AND2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U569 ( .A1(G113), .A2(n891), .ZN(n518) );
  NAND2_X1 U570 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U571 ( .A(n520), .B(KEYINPUT65), .ZN(n522) );
  INV_X1 U572 ( .A(G2105), .ZN(n523) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n523), .ZN(n890) );
  NAND2_X1 U574 ( .A1(G125), .A2(n890), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X1 U576 ( .A1(G2104), .A2(n523), .ZN(n524) );
  XNOR2_X2 U577 ( .A(n524), .B(KEYINPUT64), .ZN(n887) );
  NAND2_X1 U578 ( .A1(G101), .A2(n887), .ZN(n525) );
  XNOR2_X1 U579 ( .A(KEYINPUT23), .B(n525), .ZN(n526) );
  BUF_X1 U580 ( .A(n528), .Z(n886) );
  NAND2_X1 U581 ( .A1(G138), .A2(n886), .ZN(n530) );
  NAND2_X1 U582 ( .A1(G102), .A2(n887), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G126), .A2(n890), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G114), .A2(n891), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U587 ( .A1(n534), .A2(n533), .ZN(G164) );
  INV_X1 U588 ( .A(G651), .ZN(n537) );
  OR2_X1 U589 ( .A1(n537), .A2(n575), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n797), .A2(G78), .ZN(n536) );
  XOR2_X1 U591 ( .A(KEYINPUT68), .B(n536), .Z(n543) );
  NOR2_X1 U592 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n538), .Z(n792) );
  NAND2_X1 U594 ( .A1(G65), .A2(n792), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G53), .A2(n790), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U597 ( .A(KEYINPUT69), .B(n541), .Z(n542) );
  NOR2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n796), .A2(G91), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(G299) );
  NAND2_X1 U601 ( .A1(G64), .A2(n792), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G52), .A2(n790), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U604 ( .A1(n796), .A2(G90), .ZN(n548) );
  XOR2_X1 U605 ( .A(KEYINPUT67), .B(n548), .Z(n550) );
  NAND2_X1 U606 ( .A1(G77), .A2(n797), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n551), .Z(n552) );
  NOR2_X1 U609 ( .A1(n553), .A2(n552), .ZN(G171) );
  INV_X1 U610 ( .A(G171), .ZN(G301) );
  NAND2_X1 U611 ( .A1(n796), .A2(G89), .ZN(n554) );
  XNOR2_X1 U612 ( .A(KEYINPUT4), .B(n554), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G76), .A2(n797), .ZN(n555) );
  XOR2_X1 U614 ( .A(KEYINPUT73), .B(n555), .Z(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G63), .A2(n792), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G51), .A2(n790), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U619 ( .A(KEYINPUT74), .B(n563), .Z(n564) );
  XOR2_X1 U620 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U621 ( .A1(n796), .A2(G88), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G62), .A2(n792), .ZN(n565) );
  XOR2_X1 U623 ( .A(KEYINPUT81), .B(n565), .Z(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n790), .A2(G50), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G75), .A2(n797), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U628 ( .A1(n571), .A2(n570), .ZN(G166) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  NAND2_X1 U630 ( .A1(G49), .A2(n790), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G74), .A2(G651), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U633 ( .A1(n792), .A2(n574), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n575), .A2(G87), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n577), .A2(n576), .ZN(G288) );
  NAND2_X1 U636 ( .A1(n790), .A2(G48), .ZN(n578) );
  XNOR2_X1 U637 ( .A(KEYINPUT80), .B(n578), .ZN(n587) );
  NAND2_X1 U638 ( .A1(n792), .A2(G61), .ZN(n579) );
  XNOR2_X1 U639 ( .A(n579), .B(KEYINPUT78), .ZN(n581) );
  NAND2_X1 U640 ( .A1(G86), .A2(n796), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n797), .A2(G73), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n582), .Z(n583) );
  NOR2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT79), .B(n585), .Z(n586) );
  NAND2_X1 U646 ( .A1(n587), .A2(n586), .ZN(G305) );
  AND2_X1 U647 ( .A1(n796), .A2(G85), .ZN(n591) );
  NAND2_X1 U648 ( .A1(G60), .A2(n792), .ZN(n589) );
  NAND2_X1 U649 ( .A1(G47), .A2(n790), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U651 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U652 ( .A1(G72), .A2(n797), .ZN(n592) );
  NAND2_X1 U653 ( .A1(n593), .A2(n592), .ZN(G290) );
  NAND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n678) );
  INV_X1 U655 ( .A(n678), .ZN(n594) );
  NOR2_X1 U656 ( .A1(G164), .A2(G1384), .ZN(n679) );
  NAND2_X1 U657 ( .A1(n594), .A2(n679), .ZN(n656) );
  NAND2_X1 U658 ( .A1(G2072), .A2(n638), .ZN(n596) );
  INV_X1 U659 ( .A(G1956), .ZN(n859) );
  NOR2_X1 U660 ( .A1(n638), .A2(n859), .ZN(n597) );
  NOR2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n601) );
  INV_X1 U662 ( .A(G299), .ZN(n962) );
  NOR2_X1 U663 ( .A1(n601), .A2(n962), .ZN(n600) );
  XNOR2_X1 U664 ( .A(KEYINPUT89), .B(KEYINPUT28), .ZN(n599) );
  XNOR2_X1 U665 ( .A(n600), .B(n599), .ZN(n633) );
  NAND2_X1 U666 ( .A1(n601), .A2(n962), .ZN(n631) );
  NAND2_X1 U667 ( .A1(G56), .A2(n792), .ZN(n602) );
  XOR2_X1 U668 ( .A(KEYINPUT14), .B(n602), .Z(n608) );
  NAND2_X1 U669 ( .A1(n796), .A2(G81), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U671 ( .A1(G68), .A2(n797), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U673 ( .A(KEYINPUT13), .B(n606), .Z(n607) );
  NOR2_X1 U674 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U675 ( .A1(n790), .A2(G43), .ZN(n609) );
  NAND2_X1 U676 ( .A1(n610), .A2(n609), .ZN(n965) );
  INV_X1 U677 ( .A(G1996), .ZN(n915) );
  NOR2_X1 U678 ( .A1(n656), .A2(n915), .ZN(n611) );
  XOR2_X1 U679 ( .A(n611), .B(KEYINPUT26), .Z(n613) );
  NAND2_X1 U680 ( .A1(n656), .A2(G1341), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U682 ( .A1(n965), .A2(n614), .ZN(n623) );
  NAND2_X1 U683 ( .A1(n790), .A2(G54), .ZN(n616) );
  NAND2_X1 U684 ( .A1(G79), .A2(n797), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U686 ( .A(KEYINPUT72), .B(n617), .ZN(n621) );
  NAND2_X1 U687 ( .A1(G66), .A2(n792), .ZN(n619) );
  NAND2_X1 U688 ( .A1(G92), .A2(n796), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U690 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U691 ( .A(KEYINPUT15), .B(n622), .Z(n982) );
  OR2_X1 U692 ( .A1(n623), .A2(n982), .ZN(n629) );
  NAND2_X1 U693 ( .A1(n623), .A2(n982), .ZN(n627) );
  NAND2_X1 U694 ( .A1(G1348), .A2(n656), .ZN(n625) );
  NAND2_X1 U695 ( .A1(G2067), .A2(n638), .ZN(n624) );
  NAND2_X1 U696 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U698 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n635) );
  XNOR2_X1 U701 ( .A(KEYINPUT90), .B(KEYINPUT29), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n635), .B(n634), .ZN(n642) );
  XNOR2_X1 U703 ( .A(G2078), .B(KEYINPUT25), .ZN(n636) );
  XNOR2_X1 U704 ( .A(n636), .B(KEYINPUT86), .ZN(n917) );
  NAND2_X1 U705 ( .A1(n638), .A2(n917), .ZN(n637) );
  XNOR2_X1 U706 ( .A(n637), .B(KEYINPUT87), .ZN(n640) );
  NOR2_X1 U707 ( .A1(n638), .A2(G1961), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n643) );
  NOR2_X1 U709 ( .A1(n643), .A2(G301), .ZN(n641) );
  NOR2_X1 U710 ( .A1(n642), .A2(n641), .ZN(n654) );
  AND2_X1 U711 ( .A1(G301), .A2(n643), .ZN(n651) );
  NAND2_X1 U712 ( .A1(G8), .A2(n656), .ZN(n728) );
  NOR2_X1 U713 ( .A1(G1966), .A2(n728), .ZN(n668) );
  NOR2_X1 U714 ( .A1(G2084), .A2(n656), .ZN(n644) );
  XOR2_X1 U715 ( .A(KEYINPUT85), .B(n644), .Z(n666) );
  INV_X1 U716 ( .A(n666), .ZN(n645) );
  NAND2_X1 U717 ( .A1(G8), .A2(n645), .ZN(n646) );
  NOR2_X1 U718 ( .A1(n668), .A2(n646), .ZN(n648) );
  XNOR2_X1 U719 ( .A(KEYINPUT91), .B(KEYINPUT30), .ZN(n647) );
  XNOR2_X1 U720 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U721 ( .A1(n649), .A2(G168), .ZN(n650) );
  NOR2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n652), .B(KEYINPUT31), .ZN(n653) );
  INV_X1 U724 ( .A(n667), .ZN(n655) );
  NAND2_X1 U725 ( .A1(n655), .A2(G286), .ZN(n663) );
  INV_X1 U726 ( .A(G8), .ZN(n661) );
  NOR2_X1 U727 ( .A1(G1971), .A2(n728), .ZN(n658) );
  NOR2_X1 U728 ( .A1(G2090), .A2(n656), .ZN(n657) );
  NOR2_X1 U729 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n659), .A2(G303), .ZN(n660) );
  OR2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  AND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(n664), .ZN(n718) );
  NAND2_X1 U734 ( .A1(n666), .A2(G8), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n716) );
  NAND2_X1 U737 ( .A1(G288), .A2(G1976), .ZN(n671) );
  XOR2_X1 U738 ( .A(KEYINPUT93), .B(n671), .Z(n968) );
  AND2_X1 U739 ( .A1(n716), .A2(n968), .ZN(n672) );
  NAND2_X1 U740 ( .A1(n718), .A2(n672), .ZN(n676) );
  INV_X1 U741 ( .A(n968), .ZN(n674) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n706) );
  NOR2_X1 U743 ( .A1(G1971), .A2(G303), .ZN(n673) );
  NOR2_X1 U744 ( .A1(n706), .A2(n673), .ZN(n981) );
  OR2_X1 U745 ( .A1(n674), .A2(n981), .ZN(n675) );
  AND2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U747 ( .A(n677), .B(KEYINPUT94), .ZN(n711) );
  XOR2_X1 U748 ( .A(G1981), .B(G305), .Z(n970) );
  NOR2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n748) );
  NAND2_X1 U750 ( .A1(G140), .A2(n886), .ZN(n681) );
  NAND2_X1 U751 ( .A1(G104), .A2(n887), .ZN(n680) );
  NAND2_X1 U752 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U753 ( .A(KEYINPUT34), .B(n682), .ZN(n688) );
  NAND2_X1 U754 ( .A1(n890), .A2(G128), .ZN(n683) );
  XOR2_X1 U755 ( .A(KEYINPUT83), .B(n683), .Z(n685) );
  NAND2_X1 U756 ( .A1(n891), .A2(G116), .ZN(n684) );
  NAND2_X1 U757 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U758 ( .A(KEYINPUT35), .B(n686), .Z(n687) );
  NOR2_X1 U759 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U760 ( .A(KEYINPUT36), .B(n689), .ZN(n872) );
  XNOR2_X1 U761 ( .A(G2067), .B(KEYINPUT37), .ZN(n738) );
  NOR2_X1 U762 ( .A1(n872), .A2(n738), .ZN(n1007) );
  NAND2_X1 U763 ( .A1(n748), .A2(n1007), .ZN(n745) );
  NAND2_X1 U764 ( .A1(G131), .A2(n886), .ZN(n691) );
  NAND2_X1 U765 ( .A1(G95), .A2(n887), .ZN(n690) );
  NAND2_X1 U766 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U767 ( .A(KEYINPUT84), .B(n692), .Z(n696) );
  NAND2_X1 U768 ( .A1(G119), .A2(n890), .ZN(n694) );
  NAND2_X1 U769 ( .A1(G107), .A2(n891), .ZN(n693) );
  AND2_X1 U770 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U771 ( .A1(n696), .A2(n695), .ZN(n898) );
  NAND2_X1 U772 ( .A1(G1991), .A2(n898), .ZN(n705) );
  NAND2_X1 U773 ( .A1(G129), .A2(n890), .ZN(n698) );
  NAND2_X1 U774 ( .A1(G117), .A2(n891), .ZN(n697) );
  NAND2_X1 U775 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U776 ( .A1(n887), .A2(G105), .ZN(n699) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n699), .Z(n700) );
  NOR2_X1 U778 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U779 ( .A1(n886), .A2(G141), .ZN(n702) );
  NAND2_X1 U780 ( .A1(n703), .A2(n702), .ZN(n870) );
  NAND2_X1 U781 ( .A1(G1996), .A2(n870), .ZN(n704) );
  NAND2_X1 U782 ( .A1(n705), .A2(n704), .ZN(n1006) );
  NAND2_X1 U783 ( .A1(n748), .A2(n1006), .ZN(n741) );
  AND2_X1 U784 ( .A1(n745), .A2(n741), .ZN(n732) );
  NAND2_X1 U785 ( .A1(n970), .A2(n732), .ZN(n709) );
  NAND2_X1 U786 ( .A1(n706), .A2(KEYINPUT33), .ZN(n707) );
  NOR2_X1 U787 ( .A1(n728), .A2(n707), .ZN(n708) );
  OR2_X1 U788 ( .A1(n709), .A2(n708), .ZN(n712) );
  OR2_X1 U789 ( .A1(n728), .A2(n712), .ZN(n710) );
  NOR2_X1 U790 ( .A1(n711), .A2(n710), .ZN(n715) );
  INV_X1 U791 ( .A(n712), .ZN(n713) );
  AND2_X1 U792 ( .A1(n713), .A2(KEYINPUT33), .ZN(n714) );
  NOR2_X1 U793 ( .A1(n715), .A2(n714), .ZN(n734) );
  AND2_X1 U794 ( .A1(n716), .A2(n728), .ZN(n717) );
  NAND2_X1 U795 ( .A1(n718), .A2(n717), .ZN(n723) );
  INV_X1 U796 ( .A(n728), .ZN(n721) );
  NOR2_X1 U797 ( .A1(G2090), .A2(G303), .ZN(n719) );
  NAND2_X1 U798 ( .A1(G8), .A2(n719), .ZN(n720) );
  OR2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n722) );
  AND2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n725) );
  INV_X1 U801 ( .A(KEYINPUT95), .ZN(n724) );
  XNOR2_X1 U802 ( .A(n725), .B(n724), .ZN(n730) );
  NOR2_X1 U803 ( .A1(G1981), .A2(G305), .ZN(n726) );
  XOR2_X1 U804 ( .A(n726), .B(KEYINPUT24), .Z(n727) );
  OR2_X1 U805 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U806 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U807 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U808 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U809 ( .A(n735), .B(KEYINPUT96), .ZN(n737) );
  XNOR2_X1 U810 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U811 ( .A1(n979), .A2(n748), .ZN(n736) );
  NAND2_X1 U812 ( .A1(n737), .A2(n736), .ZN(n751) );
  NAND2_X1 U813 ( .A1(n872), .A2(n738), .ZN(n1003) );
  NOR2_X1 U814 ( .A1(G1991), .A2(n898), .ZN(n1002) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n739) );
  NOR2_X1 U816 ( .A1(n1002), .A2(n739), .ZN(n740) );
  XNOR2_X1 U817 ( .A(n740), .B(KEYINPUT97), .ZN(n742) );
  NAND2_X1 U818 ( .A1(n742), .A2(n741), .ZN(n743) );
  OR2_X1 U819 ( .A1(n870), .A2(G1996), .ZN(n998) );
  NAND2_X1 U820 ( .A1(n743), .A2(n998), .ZN(n744) );
  XOR2_X1 U821 ( .A(KEYINPUT39), .B(n744), .Z(n746) );
  NAND2_X1 U822 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U823 ( .A1(n1003), .A2(n747), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U825 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U826 ( .A(n752), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U827 ( .A(G2454), .B(KEYINPUT100), .Z(n754) );
  XNOR2_X1 U828 ( .A(G2443), .B(G2451), .ZN(n753) );
  XNOR2_X1 U829 ( .A(n754), .B(n753), .ZN(n758) );
  XOR2_X1 U830 ( .A(KEYINPUT102), .B(G2435), .Z(n756) );
  XNOR2_X1 U831 ( .A(G2438), .B(KEYINPUT98), .ZN(n755) );
  XNOR2_X1 U832 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n758), .B(n757), .ZN(n765) );
  XOR2_X1 U834 ( .A(G2430), .B(G2427), .Z(n760) );
  XNOR2_X1 U835 ( .A(KEYINPUT101), .B(G2446), .ZN(n759) );
  XNOR2_X1 U836 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U837 ( .A(n761), .B(KEYINPUT99), .Z(n763) );
  XNOR2_X1 U838 ( .A(G1348), .B(G1341), .ZN(n762) );
  XNOR2_X1 U839 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U840 ( .A(n765), .B(n764), .ZN(n766) );
  AND2_X1 U841 ( .A1(n766), .A2(G14), .ZN(G401) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U843 ( .A(G57), .ZN(G237) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  NAND2_X1 U846 ( .A1(G7), .A2(G661), .ZN(n767) );
  XNOR2_X1 U847 ( .A(n767), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U848 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n769) );
  INV_X1 U849 ( .A(G223), .ZN(n830) );
  NAND2_X1 U850 ( .A1(G567), .A2(n830), .ZN(n768) );
  XNOR2_X1 U851 ( .A(n769), .B(n768), .ZN(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n775) );
  OR2_X1 U853 ( .A1(n965), .A2(n775), .ZN(G153) );
  INV_X1 U854 ( .A(G868), .ZN(n813) );
  NOR2_X1 U855 ( .A1(G171), .A2(n813), .ZN(n770) );
  XNOR2_X1 U856 ( .A(n770), .B(KEYINPUT71), .ZN(n772) );
  OR2_X1 U857 ( .A1(G868), .A2(n982), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(G284) );
  NAND2_X1 U859 ( .A1(G868), .A2(G286), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G299), .A2(n813), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n775), .A2(G559), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n776), .A2(n982), .ZN(n777) );
  XNOR2_X1 U864 ( .A(n777), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(G868), .A2(n965), .ZN(n780) );
  NAND2_X1 U866 ( .A1(G868), .A2(n982), .ZN(n778) );
  NOR2_X1 U867 ( .A1(G559), .A2(n778), .ZN(n779) );
  NOR2_X1 U868 ( .A1(n780), .A2(n779), .ZN(G282) );
  NAND2_X1 U869 ( .A1(n890), .A2(G123), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G111), .A2(n891), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U873 ( .A1(G135), .A2(n886), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G99), .A2(n887), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n1001) );
  XNOR2_X1 U877 ( .A(n1001), .B(G2096), .ZN(n789) );
  INV_X1 U878 ( .A(G2100), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(G156) );
  NAND2_X1 U880 ( .A1(n790), .A2(G55), .ZN(n791) );
  XNOR2_X1 U881 ( .A(n791), .B(KEYINPUT76), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G67), .A2(n792), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U884 ( .A(KEYINPUT77), .B(n795), .ZN(n802) );
  NAND2_X1 U885 ( .A1(G93), .A2(n796), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G80), .A2(n797), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT75), .B(n800), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n814) );
  NAND2_X1 U890 ( .A1(n982), .A2(G559), .ZN(n811) );
  XNOR2_X1 U891 ( .A(n965), .B(n811), .ZN(n803) );
  NOR2_X1 U892 ( .A1(G860), .A2(n803), .ZN(n804) );
  XOR2_X1 U893 ( .A(n814), .B(n804), .Z(G145) );
  XNOR2_X1 U894 ( .A(G166), .B(G290), .ZN(n805) );
  XNOR2_X1 U895 ( .A(n805), .B(n965), .ZN(n806) );
  XNOR2_X1 U896 ( .A(KEYINPUT19), .B(n806), .ZN(n808) );
  XNOR2_X1 U897 ( .A(G288), .B(n962), .ZN(n807) );
  XNOR2_X1 U898 ( .A(n808), .B(n807), .ZN(n809) );
  XNOR2_X1 U899 ( .A(n809), .B(G305), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n810), .B(n814), .ZN(n836) );
  XOR2_X1 U901 ( .A(n836), .B(n811), .Z(n812) );
  NOR2_X1 U902 ( .A1(n813), .A2(n812), .ZN(n816) );
  NOR2_X1 U903 ( .A1(G868), .A2(n814), .ZN(n815) );
  NOR2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U905 ( .A(KEYINPUT82), .B(n817), .ZN(G295) );
  NAND2_X1 U906 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XOR2_X1 U907 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U908 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U909 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U910 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n822) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n822), .Z(n823) );
  NOR2_X1 U914 ( .A1(G218), .A2(n823), .ZN(n824) );
  NAND2_X1 U915 ( .A1(G96), .A2(n824), .ZN(n834) );
  NAND2_X1 U916 ( .A1(n834), .A2(G2106), .ZN(n828) );
  NAND2_X1 U917 ( .A1(G120), .A2(G108), .ZN(n825) );
  NOR2_X1 U918 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U919 ( .A1(G69), .A2(n826), .ZN(n835) );
  NAND2_X1 U920 ( .A1(n835), .A2(G567), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n912) );
  NAND2_X1 U922 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U923 ( .A1(n912), .A2(n829), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U927 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(G188) );
  XNOR2_X1 U930 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U936 ( .A(n982), .B(n836), .ZN(n838) );
  XNOR2_X1 U937 ( .A(G286), .B(G171), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  NOR2_X1 U939 ( .A1(G37), .A2(n839), .ZN(G397) );
  XOR2_X1 U940 ( .A(G2678), .B(KEYINPUT103), .Z(n841) );
  XNOR2_X1 U941 ( .A(KEYINPUT43), .B(KEYINPUT104), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n845) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2072), .Z(n843) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(n845), .B(n844), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2096), .B(G2100), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n849) );
  XOR2_X1 U949 ( .A(G2078), .B(G2084), .Z(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1961), .B(G1976), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1981), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U954 ( .A(G1966), .B(G1971), .Z(n853) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U957 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U958 ( .A(KEYINPUT105), .B(KEYINPUT41), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U960 ( .A(G2474), .B(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U962 ( .A1(n890), .A2(G124), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G136), .A2(n886), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n864) );
  XOR2_X1 U966 ( .A(KEYINPUT106), .B(n864), .Z(n866) );
  NAND2_X1 U967 ( .A1(G100), .A2(n887), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G112), .A2(n891), .ZN(n867) );
  XNOR2_X1 U970 ( .A(KEYINPUT107), .B(n867), .ZN(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U972 ( .A(G164), .B(n870), .Z(n871) );
  XNOR2_X1 U973 ( .A(n871), .B(G162), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n903) );
  NAND2_X1 U975 ( .A1(G130), .A2(n890), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G118), .A2(n891), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n886), .A2(G142), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n876), .B(KEYINPUT108), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G106), .A2(n887), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n885) );
  XOR2_X1 U984 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n883) );
  XNOR2_X1 U985 ( .A(n1001), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n901) );
  NAND2_X1 U988 ( .A1(G139), .A2(n886), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G103), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U991 ( .A1(G127), .A2(n890), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G115), .A2(n891), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U995 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(KEYINPUT109), .B(n897), .Z(n993) );
  XNOR2_X1 U997 ( .A(G160), .B(n993), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n904), .ZN(G395) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n912), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT49), .B(n905), .Z(n906) );
  XNOR2_X1 U1005 ( .A(n906), .B(KEYINPUT111), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n907), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(n910), .A2(G395), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(KEYINPUT112), .ZN(G308) );
  INV_X1 U1010 ( .A(G308), .ZN(G225) );
  INV_X1 U1011 ( .A(n912), .ZN(G319) );
  INV_X1 U1012 ( .A(G69), .ZN(G235) );
  INV_X1 U1013 ( .A(KEYINPUT55), .ZN(n1017) );
  XNOR2_X1 U1014 ( .A(G2067), .B(G26), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(G33), .B(G2072), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(G32), .B(n915), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n916), .A2(G28), .ZN(n921) );
  XOR2_X1 U1019 ( .A(G1991), .B(G25), .Z(n919) );
  XNOR2_X1 U1020 ( .A(G27), .B(n917), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT53), .B(n924), .ZN(n931) );
  XOR2_X1 U1025 ( .A(G34), .B(KEYINPUT117), .Z(n926) );
  XNOR2_X1 U1026 ( .A(G2084), .B(KEYINPUT54), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n926), .B(n925), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT116), .B(G2090), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(G35), .B(n927), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(n1017), .B(n932), .ZN(n934) );
  INV_X1 U1033 ( .A(G29), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(G11), .A2(n935), .ZN(n992) );
  XNOR2_X1 U1036 ( .A(G1981), .B(G6), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(n936), .B(KEYINPUT122), .ZN(n939) );
  XOR2_X1 U1038 ( .A(G1341), .B(G19), .Z(n937) );
  XNOR2_X1 U1039 ( .A(KEYINPUT121), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1041 ( .A(KEYINPUT123), .B(n940), .Z(n944) );
  XNOR2_X1 U1042 ( .A(KEYINPUT59), .B(G4), .ZN(n941) );
  XNOR2_X1 U1043 ( .A(n941), .B(KEYINPUT124), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(G1348), .B(n942), .ZN(n943) );
  NAND2_X1 U1045 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(G20), .B(G1956), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(KEYINPUT60), .B(n947), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(G1961), .B(G5), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(G21), .B(G1966), .ZN(n948) );
  NOR2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1052 ( .A1(n951), .A2(n950), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G1976), .B(G23), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n952) );
  NOR2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n955) );
  XOR2_X1 U1056 ( .A(G1986), .B(G24), .Z(n954) );
  NAND2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1058 ( .A(KEYINPUT58), .B(n956), .ZN(n957) );
  NOR2_X1 U1059 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1060 ( .A(KEYINPUT61), .B(n959), .Z(n960) );
  NOR2_X1 U1061 ( .A1(G16), .A2(n960), .ZN(n961) );
  XNOR2_X1 U1062 ( .A(KEYINPUT125), .B(n961), .ZN(n990) );
  XNOR2_X1 U1063 ( .A(KEYINPUT56), .B(G16), .ZN(n988) );
  XNOR2_X1 U1064 ( .A(G1956), .B(n962), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(G1971), .A2(G303), .ZN(n963) );
  NAND2_X1 U1066 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1067 ( .A(G1341), .B(n965), .ZN(n966) );
  NOR2_X1 U1068 ( .A1(n967), .A2(n966), .ZN(n969) );
  NAND2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G168), .B(G1966), .ZN(n971) );
  NAND2_X1 U1071 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1072 ( .A(n972), .B(KEYINPUT119), .ZN(n974) );
  XNOR2_X1 U1073 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n973) );
  XNOR2_X1 U1074 ( .A(n974), .B(n973), .ZN(n975) );
  NOR2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(G1961), .B(KEYINPUT120), .ZN(n977) );
  XNOR2_X1 U1077 ( .A(n977), .B(G301), .ZN(n978) );
  NOR2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1079 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1080 ( .A(G1348), .B(n982), .Z(n983) );
  NOR2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1082 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n1021) );
  XNOR2_X1 U1086 ( .A(G2072), .B(n993), .ZN(n996) );
  XOR2_X1 U1087 ( .A(G164), .B(G2078), .Z(n994) );
  XNOR2_X1 U1088 ( .A(KEYINPUT115), .B(n994), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n997), .B(KEYINPUT50), .ZN(n1015) );
  XNOR2_X1 U1091 ( .A(G2090), .B(G162), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n1000), .B(KEYINPUT51), .ZN(n1013) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(G160), .B(G2084), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1005), .B(KEYINPUT114), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT52), .B(n1016), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(G29), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT62), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(KEYINPUT126), .B(n1023), .ZN(G150) );
  INV_X1 U1109 ( .A(G150), .ZN(G311) );
endmodule

