//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(KEYINPUT69), .B1(new_n460), .B2(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n460), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n463), .A2(G137), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n465), .A2(G101), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(new_n467), .B2(new_n468), .ZN(new_n473));
  AND2_X1   g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n478));
  AND2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n467), .A2(KEYINPUT70), .A3(new_n468), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n463), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G112), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  NOR3_X1   g062(.A1(new_n479), .A2(new_n480), .A3(new_n478), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT70), .B1(new_n467), .B2(new_n468), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n463), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n481), .A2(new_n482), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(new_n493), .A3(new_n463), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  AOI211_X1 g070(.A(new_n484), .B(new_n487), .C1(new_n495), .C2(G136), .ZN(G162));
  OAI21_X1  g071(.A(G2105), .B1(KEYINPUT72), .B2(G114), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT72), .A2(G114), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n479), .A2(new_n480), .ZN(new_n501));
  NAND2_X1  g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n463), .A2(G138), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n469), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n469), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n503), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT73), .A3(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(G543), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n520), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n515), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n518), .A2(new_n528), .ZN(G166));
  NAND3_X1  g104(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n522), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n526), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n530), .B(new_n531), .C1(new_n535), .C2(KEYINPUT74), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n515), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT75), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n544), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(G651), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n526), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G90), .B1(G52), .B2(new_n522), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  AOI22_X1  g125(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n517), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n522), .A2(G43), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n526), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  AOI22_X1  g136(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n562), .A2(new_n563), .A3(new_n517), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n562), .B2(new_n517), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(KEYINPUT76), .B2(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n522), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n569), .B1(KEYINPUT76), .B2(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g145(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n522), .A2(new_n571), .A3(new_n568), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n570), .A2(new_n572), .B1(G91), .B2(new_n547), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n566), .A2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND2_X1  g151(.A1(new_n547), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n522), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n517), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n522), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n526), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n517), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n522), .A2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n526), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n522), .A2(G54), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT78), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n515), .B2(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n596), .B1(new_n599), .B2(new_n517), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g177(.A(KEYINPUT79), .B(new_n596), .C1(new_n599), .C2(new_n517), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n526), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n547), .A2(KEYINPUT10), .A3(G92), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n602), .A2(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n595), .B1(G868), .B2(new_n608), .ZN(G284));
  OAI21_X1  g184(.A(new_n595), .B1(G868), .B2(new_n608), .ZN(G321));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(G286), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(G299), .B(KEYINPUT80), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(G297));
  AOI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n608), .B1(new_n616), .B2(G860), .ZN(G148));
  OAI21_X1  g192(.A(KEYINPUT81), .B1(new_n556), .B2(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n602), .A2(new_n603), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n607), .A2(new_n606), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n621), .A2(G559), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n622), .A2(new_n611), .ZN(new_n623));
  MUX2_X1   g198(.A(new_n618), .B(KEYINPUT81), .S(new_n623), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n465), .A2(new_n469), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n493), .B1(new_n492), .B2(new_n463), .ZN(new_n630));
  AOI211_X1 g205(.A(KEYINPUT71), .B(G2105), .C1(new_n481), .C2(new_n482), .ZN(new_n631));
  OAI21_X1  g206(.A(G135), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n633), .A2(new_n634), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  AOI22_X1  g212(.A1(new_n483), .A2(G123), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n629), .A2(new_n640), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT84), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2451), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  XNOR2_X1  g222(.A(G2427), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2430), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT15), .B(G2435), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n652), .A3(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n647), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2454), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(G14), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n675), .A2(new_n676), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n674), .A2(new_n677), .A3(new_n680), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT86), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(KEYINPUT24), .B2(G34), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(KEYINPUT24), .B2(G34), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n476), .B2(G29), .ZN(new_n695));
  INV_X1    g270(.A(G2084), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  NOR2_X1   g273(.A1(G164), .A2(new_n692), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G27), .B2(new_n692), .ZN(new_n700));
  INV_X1    g275(.A(G2078), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n697), .B(new_n698), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G28), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT30), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n704), .B2(KEYINPUT30), .ZN(new_n706));
  OR2_X1    g281(.A1(KEYINPUT31), .A2(G11), .ZN(new_n707));
  NAND2_X1  g282(.A1(KEYINPUT31), .A2(G11), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n705), .A2(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n703), .B(new_n709), .C1(new_n639), .C2(new_n692), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n495), .A2(G139), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT91), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT25), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n463), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(new_n692), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n692), .B2(G33), .ZN(new_n719));
  INV_X1    g294(.A(G2072), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n702), .B(new_n710), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G5), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G171), .B2(new_n722), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(G1961), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(G1961), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n721), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(G286), .A2(G16), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT92), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n722), .A2(G21), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n719), .A2(new_n720), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n692), .A2(G32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n495), .A2(G141), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT26), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n465), .A2(G105), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n740), .B(new_n741), .C1(G129), .C2(new_n483), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(new_n692), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT27), .B(G1996), .Z(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n736), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n727), .A2(KEYINPUT93), .A3(new_n735), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n608), .A2(new_n722), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G4), .B2(new_n722), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n722), .A2(G19), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n556), .B2(new_n722), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G1341), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n692), .A2(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n692), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2090), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n761), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n752), .A2(new_n753), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n722), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1956), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n754), .A2(new_n764), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n692), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G140), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n491), .B2(new_n494), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n463), .A2(G116), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n483), .B2(G128), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(KEYINPUT89), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(G140), .B1(new_n630), .B2(new_n631), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n782), .A2(new_n783), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n773), .B1(new_n785), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n770), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n750), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n727), .A2(new_n749), .A3(new_n735), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n722), .A2(G23), .ZN(new_n795));
  INV_X1    g370(.A(G288), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n722), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n797), .B(new_n798), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n722), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n722), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT88), .Z(new_n802));
  AOI21_X1  g377(.A(new_n799), .B1(G1971), .B2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(G1971), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  NOR2_X1   g381(.A1(G6), .A2(G16), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n586), .B2(G16), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT32), .ZN(new_n809));
  INV_X1    g384(.A(G1981), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n805), .A2(new_n806), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G25), .A2(G29), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n495), .A2(G131), .ZN(new_n814));
  OAI21_X1  g389(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n815));
  INV_X1    g390(.A(G107), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G2105), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n483), .B2(G119), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(G29), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n822), .ZN(new_n824));
  INV_X1    g399(.A(G24), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n825), .A2(KEYINPUT87), .A3(G16), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT87), .B1(new_n825), .B2(G16), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n826), .B(new_n827), .C1(new_n593), .C2(new_n722), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G1986), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n823), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n812), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n806), .B1(new_n805), .B2(new_n811), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT36), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT36), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n834), .A2(new_n835), .A3(new_n812), .A4(new_n830), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n794), .B1(new_n833), .B2(new_n836), .ZN(G311));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n836), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n838), .A2(new_n793), .A3(new_n790), .ZN(G150));
  NAND2_X1  g414(.A1(new_n608), .A2(G559), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT38), .Z(new_n841));
  NAND3_X1  g416(.A1(new_n515), .A2(G93), .A3(new_n525), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n522), .A2(G55), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT95), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(new_n517), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n556), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n848), .A2(new_n556), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n841), .B(new_n855), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n857), .A2(new_n858), .A3(G860), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n851), .A2(G860), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT37), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n859), .A2(new_n861), .ZN(G145));
  INV_X1    g437(.A(new_n819), .ZN(new_n863));
  OAI21_X1  g438(.A(G142), .B1(new_n630), .B2(new_n631), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  INV_X1    g441(.A(G118), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(G2105), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n483), .B2(G130), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n627), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n865), .B1(new_n864), .B2(new_n869), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n864), .A2(new_n869), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT97), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n627), .B1(new_n876), .B2(new_n870), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n863), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n872), .B1(new_n871), .B2(new_n873), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n627), .A3(new_n870), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n819), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n781), .A2(G164), .A3(new_n784), .ZN(new_n883));
  AOI21_X1  g458(.A(G164), .B1(new_n781), .B2(new_n784), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n717), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n506), .A2(new_n508), .ZN(new_n886));
  INV_X1    g461(.A(new_n503), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n782), .A2(new_n783), .A3(new_n779), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n783), .B1(new_n782), .B2(new_n779), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n711), .A2(new_n716), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n781), .A2(G164), .A3(new_n784), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n885), .A2(new_n744), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n744), .B1(new_n885), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n882), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n892), .B1(new_n891), .B2(new_n893), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n743), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n878), .A2(new_n881), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n885), .A2(new_n744), .A3(new_n894), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n639), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT96), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(KEYINPUT96), .ZN(new_n908));
  OAI21_X1  g483(.A(G160), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n905), .A2(KEYINPUT96), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n476), .A3(new_n906), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n909), .A2(new_n911), .A3(G162), .ZN(new_n912));
  AOI21_X1  g487(.A(G162), .B1(new_n909), .B2(new_n911), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n904), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n903), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT98), .A4(new_n902), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n912), .A2(new_n913), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n917), .A2(new_n918), .A3(new_n897), .A4(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n915), .A2(KEYINPUT99), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT99), .B1(new_n915), .B2(new_n920), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n914), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  INV_X1    g503(.A(new_n917), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n897), .A2(new_n918), .A3(new_n919), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n927), .B(new_n928), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n915), .A2(KEYINPUT99), .A3(new_n920), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT40), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n924), .A2(new_n935), .ZN(G395));
  XOR2_X1   g511(.A(new_n586), .B(new_n593), .Z(new_n937));
  XNOR2_X1  g512(.A(G166), .B(G288), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT42), .B1(new_n939), .B2(KEYINPUT101), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(KEYINPUT101), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n622), .B(new_n855), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT100), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n566), .A2(new_n945), .A3(new_n573), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n608), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n566), .B2(new_n573), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(KEYINPUT100), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n950), .A2(new_n608), .A3(new_n946), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n951), .A3(KEYINPUT41), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n947), .A2(new_n948), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n621), .A2(KEYINPUT100), .A3(G299), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n944), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n949), .A2(new_n951), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n944), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n943), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n942), .A2(new_n961), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n851), .A2(new_n611), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n954), .A2(new_n955), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n853), .A2(G301), .A3(new_n854), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G301), .B1(new_n853), .B2(new_n854), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n973), .A2(new_n974), .A3(G286), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n855), .A2(G171), .ZN(new_n976));
  AOI21_X1  g551(.A(G168), .B1(new_n976), .B2(new_n972), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n971), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G286), .B1(new_n973), .B2(new_n974), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(G168), .A3(new_n972), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n956), .A2(new_n979), .A3(new_n980), .A4(new_n952), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n939), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n981), .A3(new_n939), .ZN(new_n985));
  AND4_X1   g560(.A1(new_n970), .A2(new_n984), .A3(new_n928), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n982), .B2(new_n983), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n970), .B1(new_n987), .B2(new_n985), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n989), .B1(new_n986), .B2(new_n988), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(G397));
  XNOR2_X1  g567(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n471), .A2(new_n475), .A3(new_n995), .A4(G40), .ZN(new_n996));
  INV_X1    g571(.A(G40), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT104), .B1(new_n476), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n994), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n889), .A2(new_n890), .A3(G2067), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n787), .B1(new_n781), .B2(new_n784), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n785), .A2(G2067), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n787), .A3(new_n784), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(KEYINPUT105), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1000), .B1(new_n1008), .B2(new_n744), .ZN(new_n1009));
  INV_X1    g584(.A(G1996), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n744), .A2(new_n999), .A3(new_n1010), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(KEYINPUT106), .A3(new_n1013), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n863), .A2(new_n822), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1000), .B1(new_n1019), .B2(new_n1006), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n819), .A2(new_n821), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n999), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G290), .A2(G1986), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n999), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n1024), .B(KEYINPUT48), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1016), .A2(new_n1017), .A3(new_n1022), .A4(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT46), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT126), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT126), .B(KEYINPUT46), .Z(new_n1029));
  NAND2_X1  g604(.A1(new_n999), .A2(new_n1010), .ZN(new_n1030));
  MUX2_X1   g605(.A(new_n1028), .B(new_n1029), .S(new_n1030), .Z(new_n1031));
  NOR2_X1   g606(.A1(new_n1009), .A2(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n1032), .B(KEYINPUT47), .Z(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1020), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT61), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1037));
  XNOR2_X1  g612(.A(G299), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1956), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n998), .A2(new_n996), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n888), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1039), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n1045), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1040), .A2(new_n994), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT56), .B(G2072), .Z(new_n1052));
  OR2_X1    g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1038), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1038), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1036), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT60), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1040), .A2(new_n1041), .A3(new_n1046), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n753), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n888), .A2(new_n1045), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n996), .B2(new_n998), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n787), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n608), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(new_n1062), .A3(new_n621), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1057), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(KEYINPUT120), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1040), .A2(new_n994), .A3(new_n1010), .A4(new_n1050), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(KEYINPUT58), .B(G1341), .Z(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1060), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n1040), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n556), .B(new_n1068), .C1(new_n1070), .C2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1059), .A2(new_n1062), .A3(new_n1057), .A4(new_n608), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1074), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n852), .B1(new_n1077), .B2(new_n1069), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1079));
  OAI211_X1 g654(.A(new_n1075), .B(new_n1076), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1066), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1038), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1038), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(KEYINPUT61), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1056), .A2(new_n1081), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1064), .B(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1089), .B2(new_n1055), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1050), .A2(KEYINPUT53), .A3(new_n701), .ZN(new_n1092));
  INV_X1    g667(.A(new_n994), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n471), .A2(KEYINPUT124), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n471), .A2(KEYINPUT124), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1094), .A2(G40), .A3(new_n475), .A4(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n1097));
  OR3_X1    g672(.A1(new_n1093), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1092), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G301), .B(KEYINPUT54), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT123), .B(new_n1103), .C1(new_n1051), .C2(G2078), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1040), .A2(new_n1041), .A3(new_n1046), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(G1961), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1103), .B1(new_n1051), .B2(G2078), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT45), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1060), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1112), .B(new_n1040), .C1(new_n1060), .C2(new_n993), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n701), .A2(KEYINPUT53), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(new_n1109), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1101), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1110), .A2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT109), .B(G8), .ZN(new_n1119));
  NOR2_X1   g694(.A1(G168), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n734), .A2(new_n1113), .B1(new_n1105), .B2(new_n696), .ZN(new_n1122));
  INV_X1    g697(.A(G8), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT121), .B(KEYINPUT51), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1113), .A2(new_n734), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1105), .A2(new_n696), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1119), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1120), .A2(KEYINPUT51), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT122), .B1(new_n1122), .B2(new_n1119), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1126), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1122), .A2(new_n1121), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1118), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT113), .B1(new_n586), .B2(new_n810), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT113), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1142), .B(G1981), .C1(new_n582), .C2(new_n585), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT112), .B(G1981), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n586), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT114), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT49), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT49), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1061), .A2(new_n1119), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n796), .A2(G1976), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1073), .A2(new_n1040), .ZN(new_n1155));
  INV_X1    g730(.A(G1976), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT52), .B1(G288), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1154), .A2(new_n1155), .A3(new_n1131), .A4(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT111), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1154), .A2(new_n1155), .A3(new_n1131), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT110), .B1(new_n1160), .B2(KEYINPUT52), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1160), .A2(KEYINPUT52), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT110), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1153), .B(new_n1159), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT108), .B(G2090), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1105), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(KEYINPUT107), .B(G1971), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1051), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1123), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(G166), .A2(new_n1123), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT55), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1048), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(new_n1046), .A3(new_n1043), .A4(new_n1166), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1119), .B1(new_n1175), .B2(new_n1169), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1173), .B1(new_n1176), .B2(new_n1172), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1165), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1091), .A2(new_n1140), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1133), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1119), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1180), .B1(new_n1181), .B2(new_n1130), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1182), .A2(new_n1135), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT62), .B1(new_n1183), .B2(new_n1138), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1137), .A2(new_n1185), .A3(new_n1139), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1116), .A2(G171), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1165), .A2(new_n1177), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1184), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1181), .A2(G168), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1165), .A2(new_n1177), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT117), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1172), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1193), .B(new_n1170), .ZN(new_n1194));
  NAND4_X1  g769(.A1(new_n1194), .A2(KEYINPUT63), .A3(G168), .A4(new_n1181), .ZN(new_n1195));
  OAI22_X1  g770(.A1(new_n1191), .A2(KEYINPUT63), .B1(new_n1195), .B2(new_n1165), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1165), .A2(new_n1173), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1153), .A2(new_n1156), .A3(new_n796), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1145), .B(KEYINPUT115), .Z(new_n1199));
  NAND2_X1  g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1152), .B2(new_n1200), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1179), .A2(new_n1189), .A3(new_n1196), .A4(new_n1201), .ZN(new_n1202));
  AND2_X1   g777(.A1(G290), .A2(G1986), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n999), .B1(new_n1203), .B2(new_n1023), .ZN(new_n1204));
  AND4_X1   g779(.A1(new_n1204), .A2(new_n1016), .A3(new_n1017), .A4(new_n1022), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1035), .A2(new_n1206), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g782(.A1(G401), .A2(new_n458), .A3(G227), .A4(G229), .ZN(new_n1209));
  OAI21_X1  g783(.A(new_n1209), .B1(new_n986), .B2(new_n988), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n933), .B2(new_n934), .ZN(G308));
  OAI221_X1 g785(.A(new_n1209), .B1(new_n986), .B2(new_n988), .C1(new_n921), .C2(new_n922), .ZN(G225));
endmodule


