//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1208, new_n1209,
    new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G125), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g038(.A(KEYINPUT66), .B(G125), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  XNOR2_X1  g041(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n470), .C1(new_n459), .C2(new_n460), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n459), .A2(new_n460), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n470), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n479), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(G2105), .B1(KEYINPUT68), .B2(G114), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT68), .A2(G114), .ZN(new_n491));
  OAI211_X1 g066(.A(G2104), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n459), .B2(new_n460), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n481), .A2(new_n482), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(new_n496), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n494), .B1(new_n498), .B2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n510), .A2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n511), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n509), .B1(new_n531), .B2(KEYINPUT69), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n532), .B1(KEYINPUT69), .B2(new_n531), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n507), .A2(new_n511), .ZN(new_n534));
  OR2_X1    g109(.A1(KEYINPUT6), .A2(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(KEYINPUT6), .A2(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n504), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n534), .A2(G90), .B1(G52), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n533), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n509), .ZN(new_n541));
  INV_X1    g116(.A(G81), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n512), .A2(new_n542), .B1(new_n514), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT70), .Z(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT71), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(new_n534), .A2(G91), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  AND3_X1   g129(.A1(new_n537), .A2(new_n554), .A3(G53), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n554), .B1(new_n537), .B2(G53), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n553), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  NOR3_X1   g134(.A1(new_n522), .A2(new_n523), .A3(KEYINPUT72), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT72), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n505), .B2(new_n506), .ZN(new_n562));
  OAI21_X1  g137(.A(G65), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n559), .B1(new_n566), .B2(G651), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT72), .B1(new_n522), .B2(new_n523), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n505), .A2(new_n561), .A3(new_n506), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n559), .B(G651), .C1(new_n571), .C2(new_n564), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n558), .B1(new_n567), .B2(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n533), .A2(new_n538), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n505), .A2(new_n578), .A3(new_n506), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n537), .A2(G49), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n507), .A2(new_n511), .A3(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(G288));
  INV_X1    g157(.A(KEYINPUT74), .ZN(new_n583));
  INV_X1    g158(.A(G73), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n504), .ZN(new_n585));
  NAND3_X1  g160(.A1(KEYINPUT74), .A2(G73), .A3(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n524), .C2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G48), .B2(new_n537), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n534), .A2(G86), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n592), .A2(KEYINPUT75), .A3(new_n509), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT75), .B1(new_n592), .B2(new_n509), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n534), .A2(G85), .B1(G47), .B2(new_n537), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT77), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n569), .A2(new_n570), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G66), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT78), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n509), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(new_n601), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n512), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G54), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n609), .B1(new_n514), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n537), .A2(KEYINPUT76), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n605), .A2(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n597), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n597), .B1(new_n614), .B2(G868), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n564), .B1(new_n600), .B2(G65), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT73), .B1(new_n618), .B2(new_n509), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n557), .B1(new_n619), .B2(new_n572), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G860), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT79), .Z(G148));
  NAND2_X1  g200(.A1(new_n614), .A2(new_n623), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n499), .A2(new_n473), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n478), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n483), .A2(G123), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n635), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT81), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT14), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT82), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n649), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n645), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n652), .A2(new_n653), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n650), .A2(KEYINPUT82), .A3(new_n651), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n659), .A2(new_n644), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n643), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n655), .A3(new_n645), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n644), .ZN(new_n663));
  INV_X1    g238(.A(new_n643), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2451), .B(G2454), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT16), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n661), .A2(new_n668), .A3(new_n665), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n677), .B2(KEYINPUT18), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT83), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n633), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT18), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(KEYINPUT17), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n675), .A2(new_n676), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n680), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(KEYINPUT84), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT19), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(KEYINPUT84), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT87), .Z(new_n698));
  AND2_X1   g273(.A1(new_n687), .A2(new_n688), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n691), .B(KEYINPUT19), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n689), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(KEYINPUT86), .B2(new_n692), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT86), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n703), .C1(new_n699), .C2(new_n689), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n696), .A2(new_n698), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1991), .B(G1996), .Z(new_n708));
  AOI21_X1  g283(.A(new_n698), .B1(new_n696), .B2(new_n705), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n712), .ZN(new_n715));
  INV_X1    g290(.A(new_n708), .ZN(new_n716));
  INV_X1    g291(.A(new_n709), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n706), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n715), .B1(new_n718), .B2(new_n710), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n714), .A2(new_n719), .ZN(G229));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G26), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n478), .A2(G140), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT92), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n726));
  INV_X1    g301(.A(G116), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G2105), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G128), .B2(new_n483), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n730), .A2(KEYINPUT93), .A3(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(KEYINPUT93), .B1(new_n730), .B2(G29), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n723), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G2067), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G35), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G162), .B2(G29), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT29), .Z(new_n737));
  INV_X1    g312(.A(G2090), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NOR2_X1   g315(.A1(G171), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G5), .B2(new_n740), .ZN(new_n742));
  INV_X1    g317(.A(G1961), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n721), .B1(KEYINPUT24), .B2(G34), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(KEYINPUT24), .B2(G34), .ZN(new_n747));
  INV_X1    g322(.A(G160), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2084), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n737), .A2(new_n738), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n734), .A2(new_n745), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G4), .A2(G16), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n614), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT89), .B(G16), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G20), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT100), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n740), .B2(new_n620), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n640), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n765), .A2(KEYINPUT98), .A3(G29), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n640), .B2(new_n721), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT97), .ZN(new_n770));
  INV_X1    g345(.A(G28), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(KEYINPUT30), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n771), .B2(KEYINPUT30), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n766), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT99), .Z(new_n776));
  NOR2_X1   g351(.A1(G286), .A2(new_n740), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT96), .B1(G16), .B2(G21), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1966), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT25), .ZN(new_n785));
  NAND2_X1  g360(.A1(G115), .A2(G2104), .ZN(new_n786));
  INV_X1    g361(.A(G127), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n477), .B2(new_n787), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n788), .A2(G2105), .B1(new_n478), .B2(G139), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  NAND2_X1  g366(.A1(new_n791), .A2(G2072), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n721), .A2(G27), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G164), .B2(new_n721), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n776), .A2(new_n782), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n781), .A2(G1966), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n791), .A2(G2072), .ZN(new_n799));
  INV_X1    g374(.A(new_n758), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G19), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n545), .B2(new_n800), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(G1341), .Z(new_n803));
  NAND2_X1  g378(.A1(new_n721), .A2(G32), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n473), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n483), .A2(G129), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT26), .Z(new_n808));
  NAND3_X1  g383(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n804), .B1(new_n810), .B2(new_n721), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT27), .B(G1996), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n798), .A2(new_n799), .A3(new_n803), .A4(new_n814), .ZN(new_n815));
  OAI22_X1  g390(.A1(new_n742), .A2(new_n743), .B1(new_n750), .B2(new_n749), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n797), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n753), .A2(new_n757), .A3(new_n764), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n478), .A2(G131), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n483), .A2(G119), .ZN(new_n820));
  OR2_X1    g395(.A1(G95), .A2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  MUX2_X1   g398(.A(G25), .B(new_n823), .S(G29), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT88), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G1991), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(G290), .A2(KEYINPUT90), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n758), .B1(G290), .B2(KEYINPUT90), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n829), .A2(new_n830), .B1(G24), .B2(new_n758), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n828), .B1(G1986), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n832), .A2(G1986), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n800), .A2(G22), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G166), .B2(new_n800), .ZN(new_n836));
  INV_X1    g411(.A(G1971), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n740), .A2(G23), .ZN(new_n839));
  INV_X1    g414(.A(G288), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n740), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT33), .B(G1976), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n740), .A2(G6), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G305), .B2(G16), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT32), .B(G1981), .Z(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n838), .A2(new_n843), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n833), .A2(new_n834), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT91), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(new_n852), .A3(KEYINPUT34), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n849), .B2(KEYINPUT34), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n851), .A2(KEYINPUT36), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT36), .B1(new_n851), .B2(new_n856), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n818), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(G311));
  INV_X1    g436(.A(new_n859), .ZN(G150));
  NAND2_X1  g437(.A1(new_n604), .A2(new_n613), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n623), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT38), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(new_n509), .ZN(new_n867));
  INV_X1    g442(.A(G93), .ZN(new_n868));
  INV_X1    g443(.A(G55), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n512), .A2(new_n868), .B1(new_n514), .B2(new_n869), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n867), .A2(new_n870), .A3(KEYINPUT102), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT102), .B1(new_n867), .B2(new_n870), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT103), .B1(new_n873), .B2(new_n545), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n545), .B1(new_n867), .B2(new_n870), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n876));
  INV_X1    g451(.A(new_n545), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n871), .A2(new_n876), .A3(new_n877), .A4(new_n872), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n865), .B(new_n879), .Z(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(KEYINPUT39), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(KEYINPUT104), .Z(new_n882));
  AOI21_X1  g457(.A(G860), .B1(new_n880), .B2(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n873), .A2(G860), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT37), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(G145));
  XOR2_X1   g462(.A(KEYINPUT107), .B(G37), .Z(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G160), .B(KEYINPUT105), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n487), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n765), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n890), .B(G162), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n640), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n730), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(G164), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n498), .A2(new_n501), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT68), .ZN(new_n899));
  INV_X1    g474(.A(G114), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(KEYINPUT68), .A2(G114), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(G2105), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(G126), .A2(new_n483), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n898), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n730), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n483), .A2(G130), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT106), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  INV_X1    g487(.A(G118), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(G2105), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n478), .A2(G142), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR3_X1   g491(.A1(new_n911), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n909), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n917), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n897), .A2(new_n908), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n790), .B(new_n810), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n631), .B(new_n823), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n790), .B(new_n809), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n922), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n918), .A2(new_n920), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n918), .A2(new_n920), .B1(new_n924), .B2(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n895), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n927), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n892), .B(new_n894), .C1(new_n931), .C2(new_n928), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n889), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g509(.A(new_n626), .B(KEYINPUT108), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(new_n879), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n863), .B(new_n620), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT41), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n614), .A2(new_n620), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n863), .A2(G299), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n936), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n937), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n936), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(G290), .B(G305), .ZN(new_n948));
  XNOR2_X1  g523(.A(G166), .B(G288), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n948), .B(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n945), .A2(new_n947), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n945), .B2(new_n947), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n873), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n958), .B1(G868), .B2(new_n959), .ZN(G295));
  OAI21_X1  g535(.A(new_n958), .B1(G868), .B2(new_n959), .ZN(G331));
  OAI21_X1  g536(.A(KEYINPUT110), .B1(G171), .B2(G286), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n963));
  NAND3_X1  g538(.A1(G301), .A2(new_n963), .A3(G168), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(G301), .B2(G168), .ZN(new_n966));
  NAND4_X1  g541(.A1(G286), .A2(new_n533), .A3(KEYINPUT111), .A4(new_n538), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n962), .A2(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n878), .A2(new_n875), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n874), .A3(new_n969), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n962), .A2(new_n964), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n966), .A2(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n879), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n970), .A2(new_n973), .B1(new_n938), .B2(new_n942), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n973), .A2(new_n970), .A3(new_n946), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n950), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n970), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n943), .ZN(new_n978));
  INV_X1    g553(.A(new_n950), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n973), .A2(new_n970), .A3(new_n946), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(G37), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n889), .C1(new_n976), .C2(new_n981), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT44), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n974), .A2(new_n975), .A3(new_n950), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n984), .B(new_n888), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n984), .B2(new_n982), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n986), .B1(new_n991), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n469), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n999), .A2(G1996), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n1000), .A2(new_n809), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n730), .B(G2067), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G2067), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n730), .B(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n810), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1008), .B(new_n998), .C1(new_n1009), .C2(G1996), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n823), .A2(new_n827), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n823), .A2(new_n827), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n998), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OR3_X1    g588(.A1(new_n999), .A2(G1986), .A3(G290), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n998), .A2(G1986), .A3(G290), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT112), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n1001), .A2(new_n1010), .A3(new_n1013), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n907), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n995), .B1(new_n468), .B2(G2105), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n907), .A2(new_n1023), .A3(new_n1019), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1021), .A2(new_n750), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n907), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n994), .A2(new_n1026), .A3(new_n1022), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(G1966), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(G8), .A3(G286), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1025), .B(G168), .C1(new_n1027), .C2(G1966), .ZN(new_n1030));
  AND2_X1   g605(.A1(KEYINPUT124), .A2(G8), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1030), .A2(KEYINPUT51), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1029), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT62), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT62), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1036), .B(new_n1029), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT49), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT117), .B(G86), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n534), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n589), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n585), .A2(new_n586), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n587), .B1(new_n505), .B2(new_n506), .ZN(new_n1044));
  OAI21_X1  g619(.A(G651), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n537), .A2(G48), .ZN(new_n1046));
  AND4_X1   g621(.A1(new_n1039), .A2(new_n590), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1038), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1041), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G1981), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n589), .A2(new_n1039), .A3(new_n590), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1051), .A3(KEYINPUT49), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1384), .B1(new_n898), .B2(new_n906), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1022), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1048), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n580), .A2(G1976), .A3(new_n581), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT114), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n580), .A2(new_n1059), .A3(G1976), .A4(new_n581), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT115), .B(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n580), .B2(new_n581), .ZN(new_n1065));
  OR3_X1    g640(.A1(new_n1065), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT116), .B1(new_n1065), .B2(KEYINPUT52), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1055), .A3(new_n1061), .A4(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1056), .A2(new_n1063), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G303), .A2(G8), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n994), .A2(new_n1026), .A3(new_n1022), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n837), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1021), .A2(new_n738), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1053), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1070), .B(KEYINPUT55), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1022), .B1(new_n1054), .B2(new_n1023), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1024), .A2(KEYINPUT118), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1054), .A2(new_n1081), .A3(new_n1023), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1083), .A2(new_n738), .B1(new_n837), .B2(new_n1073), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1078), .B1(new_n1084), .B2(new_n1053), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n997), .B1(new_n993), .B2(new_n1020), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1086), .A2(KEYINPUT53), .A3(new_n795), .A4(new_n1026), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n994), .A2(new_n795), .A3(new_n1026), .A4(new_n1022), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1024), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n743), .B1(new_n1091), .B2(new_n1079), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1077), .A2(new_n1085), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1035), .A2(new_n1037), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1076), .A2(new_n1072), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n1069), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1056), .ZN(new_n1099));
  OR2_X1    g674(.A1(G288), .A2(G1976), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1051), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1055), .B2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n994), .A2(new_n1026), .A3(new_n1022), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1083), .B2(G1956), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n1106));
  NAND3_X1  g681(.A1(G299), .A2(new_n1106), .A3(KEYINPUT57), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n620), .B2(KEYINPUT120), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1105), .A2(new_n1110), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n756), .B1(new_n1091), .B2(new_n1079), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1022), .A2(new_n1054), .A3(new_n1005), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n614), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1111), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  NOR4_X1   g692(.A1(G164), .A2(KEYINPUT118), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1081), .B1(new_n1054), .B2(new_n1023), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n763), .B1(new_n1120), .B2(new_n1079), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1121), .A2(new_n1104), .B1(new_n1109), .B2(new_n1107), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT61), .B1(new_n1122), .B2(new_n1112), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n1109), .A3(new_n1107), .A4(new_n1104), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n1111), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1123), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1113), .A2(new_n1114), .A3(KEYINPUT60), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n863), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT121), .B(G1996), .Z(new_n1131));
  NAND4_X1  g706(.A1(new_n994), .A2(new_n1026), .A3(new_n1022), .A4(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  OAI21_X1  g708(.A(new_n1133), .B1(new_n997), .B2(new_n1020), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n545), .A4(new_n1138), .ZN(new_n1139));
  AOI211_X1 g714(.A(KEYINPUT123), .B(new_n877), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1140), .B2(KEYINPUT59), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1113), .A2(new_n863), .A3(KEYINPUT60), .A4(new_n1114), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n877), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1130), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1117), .B1(new_n1127), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1092), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT125), .B(new_n743), .C1(new_n1091), .C2(new_n1079), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1087), .A3(new_n1090), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(G171), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1152), .B2(new_n1094), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1069), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1085), .A2(new_n1097), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(G171), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1087), .A2(new_n1090), .A3(G301), .A4(new_n1092), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(KEYINPUT54), .A3(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1153), .A2(new_n1155), .A3(new_n1034), .A4(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1096), .B(new_n1102), .C1(new_n1146), .C2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1028), .A2(G8), .A3(G168), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1085), .A2(new_n1161), .A3(new_n1097), .A4(new_n1154), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT119), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1163), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1161), .B(KEYINPUT63), .C1(new_n1072), .C2(new_n1076), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1077), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1166), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1018), .B1(new_n1160), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1010), .A2(new_n1001), .A3(new_n1013), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT47), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1008), .A2(new_n998), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1000), .B(KEYINPUT46), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1006), .A2(KEYINPUT113), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n809), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1177), .B(new_n1175), .C1(new_n1181), .C2(new_n999), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1174), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1010), .A2(new_n1001), .A3(new_n1011), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n896), .A2(new_n1005), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n999), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1172), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(KEYINPUT126), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1172), .A2(new_n1191), .A3(new_n1188), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g768(.A(G319), .ZN(new_n1195));
  OR2_X1    g769(.A1(G227), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n714), .B2(new_n719), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n672), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g772(.A1(new_n1198), .A2(new_n933), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n976), .A2(new_n981), .ZN(new_n1200));
  INV_X1    g774(.A(G37), .ZN(new_n1201));
  AOI21_X1  g775(.A(new_n984), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g776(.A(KEYINPUT43), .B(new_n889), .C1(new_n976), .C2(new_n981), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n1199), .B(KEYINPUT127), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  INV_X1    g778(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g779(.A(KEYINPUT127), .B1(new_n990), .B2(new_n1199), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1205), .A2(new_n1206), .ZN(G308));
  NAND2_X1  g781(.A1(new_n990), .A2(new_n1199), .ZN(new_n1208));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1210), .A2(new_n1204), .ZN(G225));
endmodule


