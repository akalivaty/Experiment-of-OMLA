

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724;

  INV_X2 U367 ( .A(G953), .ZN(n691) );
  INV_X1 U368 ( .A(n585), .ZN(n634) );
  NAND2_X1 U369 ( .A1(n619), .A2(n622), .ZN(n585) );
  OR2_X1 U370 ( .A1(n599), .A2(G902), .ZN(n394) );
  NOR2_X2 U371 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U372 ( .A1(G902), .A2(n667), .ZN(n444) );
  XNOR2_X2 U373 ( .A(n573), .B(KEYINPUT35), .ZN(n720) );
  XNOR2_X2 U374 ( .A(n460), .B(n461), .ZN(n482) );
  XNOR2_X2 U375 ( .A(n538), .B(KEYINPUT40), .ZN(n723) );
  NOR2_X1 U376 ( .A1(n569), .A2(n639), .ZN(n579) );
  XNOR2_X1 U377 ( .A(n398), .B(n354), .ZN(n690) );
  NAND2_X1 U378 ( .A1(n399), .A2(n347), .ZN(n398) );
  XNOR2_X1 U379 ( .A(n576), .B(n575), .ZN(n399) );
  XNOR2_X1 U380 ( .A(n369), .B(n414), .ZN(n722) );
  XNOR2_X1 U381 ( .A(n467), .B(KEYINPUT101), .ZN(n619) );
  XNOR2_X1 U382 ( .A(n579), .B(n364), .ZN(n570) );
  NAND2_X1 U383 ( .A1(n564), .A2(n556), .ZN(n639) );
  XNOR2_X1 U384 ( .A(n496), .B(n376), .ZN(n698) );
  XNOR2_X1 U385 ( .A(n433), .B(n432), .ZN(n459) );
  XNOR2_X1 U386 ( .A(G146), .B(KEYINPUT4), .ZN(n706) );
  XNOR2_X1 U387 ( .A(G107), .B(G110), .ZN(n700) );
  AND2_X1 U388 ( .A1(n595), .A2(n409), .ZN(n681) );
  NOR2_X2 U389 ( .A1(n687), .A2(G902), .ZN(n367) );
  XNOR2_X2 U390 ( .A(n421), .B(G143), .ZN(n433) );
  XNOR2_X2 U391 ( .A(G128), .B(KEYINPUT65), .ZN(n421) );
  XNOR2_X1 U392 ( .A(n567), .B(n566), .ZN(n577) );
  INV_X1 U393 ( .A(KEYINPUT86), .ZN(n566) );
  NAND2_X1 U394 ( .A1(n722), .A2(n611), .ZN(n567) );
  NOR2_X1 U395 ( .A1(G237), .A2(G953), .ZN(n450) );
  XNOR2_X1 U396 ( .A(n428), .B(n427), .ZN(n496) );
  XNOR2_X1 U397 ( .A(n705), .B(n435), .ZN(n498) );
  XNOR2_X1 U398 ( .A(n706), .B(n413), .ZN(n435) );
  INV_X1 U399 ( .A(G101), .ZN(n413) );
  XNOR2_X1 U400 ( .A(n412), .B(n411), .ZN(n558) );
  INV_X1 U401 ( .A(KEYINPUT0), .ZN(n411) );
  NAND2_X1 U402 ( .A1(n555), .A2(n554), .ZN(n412) );
  XNOR2_X1 U403 ( .A(n459), .B(n408), .ZN(n705) );
  XNOR2_X1 U404 ( .A(n434), .B(G137), .ZN(n408) );
  XOR2_X1 U405 ( .A(KEYINPUT69), .B(G131), .Z(n434) );
  XNOR2_X1 U406 ( .A(G122), .B(G104), .ZN(n447) );
  XOR2_X1 U407 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n461) );
  OR2_X1 U408 ( .A1(G237), .A2(G902), .ZN(n504) );
  XNOR2_X1 U409 ( .A(n548), .B(n402), .ZN(n630) );
  INV_X1 U410 ( .A(KEYINPUT38), .ZN(n402) );
  XNOR2_X1 U411 ( .A(n518), .B(KEYINPUT1), .ZN(n569) );
  OR2_X1 U412 ( .A1(n568), .A2(n506), .ZN(n407) );
  NAND2_X1 U413 ( .A1(n386), .A2(n587), .ZN(n388) );
  NOR2_X1 U414 ( .A1(n570), .A2(n391), .ZN(n386) );
  INV_X1 U415 ( .A(KEYINPUT34), .ZN(n392) );
  INV_X1 U416 ( .A(G472), .ZN(n393) );
  AND2_X1 U417 ( .A1(n396), .A2(n418), .ZN(n715) );
  XNOR2_X1 U418 ( .A(G137), .B(G128), .ZN(n479) );
  XNOR2_X1 U419 ( .A(G119), .B(G110), .ZN(n475) );
  XNOR2_X1 U420 ( .A(n451), .B(n361), .ZN(n677) );
  XNOR2_X1 U421 ( .A(n452), .B(n352), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n374), .B(n373), .ZN(n372) );
  XNOR2_X1 U423 ( .A(n426), .B(n698), .ZN(n375) );
  XNOR2_X1 U424 ( .A(n439), .B(n435), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n559), .B(n371), .ZN(n370) );
  INV_X1 U426 ( .A(KEYINPUT22), .ZN(n371) );
  INV_X1 U427 ( .A(KEYINPUT82), .ZN(n359) );
  INV_X1 U428 ( .A(KEYINPUT44), .ZN(n575) );
  XOR2_X1 U429 ( .A(KEYINPUT97), .B(G131), .Z(n446) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n445) );
  XOR2_X1 U431 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n449) );
  XNOR2_X1 U432 ( .A(G104), .B(G140), .ZN(n436) );
  XOR2_X1 U433 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n437) );
  XNOR2_X1 U434 ( .A(n700), .B(KEYINPUT71), .ZN(n439) );
  XOR2_X1 U435 ( .A(KEYINPUT77), .B(KEYINPUT18), .Z(n425) );
  XNOR2_X1 U436 ( .A(n422), .B(n346), .ZN(n374) );
  INV_X1 U437 ( .A(KEYINPUT104), .ZN(n364) );
  INV_X1 U438 ( .A(KEYINPUT33), .ZN(n391) );
  XNOR2_X1 U439 ( .A(n498), .B(n395), .ZN(n599) );
  XNOR2_X1 U440 ( .A(n497), .B(n499), .ZN(n395) );
  XNOR2_X1 U441 ( .A(n429), .B(n377), .ZN(n376) );
  INV_X1 U442 ( .A(KEYINPUT16), .ZN(n377) );
  XNOR2_X1 U443 ( .A(G116), .B(G107), .ZN(n456) );
  INV_X1 U444 ( .A(G134), .ZN(n432) );
  XNOR2_X1 U445 ( .A(n358), .B(n592), .ZN(n595) );
  AND2_X1 U446 ( .A1(n595), .A2(n594), .ZN(n674) );
  XNOR2_X1 U447 ( .A(n404), .B(KEYINPUT106), .ZN(n543) );
  XNOR2_X1 U448 ( .A(n407), .B(KEYINPUT105), .ZN(n406) );
  INV_X1 U449 ( .A(n619), .ZN(n405) );
  AND2_X1 U450 ( .A1(n388), .A2(n558), .ZN(n385) );
  OR2_X1 U451 ( .A1(n521), .A2(n520), .ZN(n536) );
  OR2_X1 U452 ( .A1(n501), .A2(n673), .ZN(n403) );
  XNOR2_X1 U453 ( .A(n455), .B(n454), .ZN(n529) );
  XNOR2_X1 U454 ( .A(n453), .B(G475), .ZN(n454) );
  NOR2_X1 U455 ( .A1(n518), .A2(n639), .ZN(n583) );
  XNOR2_X1 U456 ( .A(n486), .B(n485), .ZN(n687) );
  XNOR2_X1 U457 ( .A(n484), .B(n483), .ZN(n485) );
  BUF_X1 U458 ( .A(n681), .Z(n685) );
  XNOR2_X1 U459 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n724) );
  XNOR2_X1 U461 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n400) );
  OR2_X1 U462 ( .A1(n662), .A2(n534), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n562), .B(n415), .ZN(n414) );
  INV_X1 U464 ( .A(KEYINPUT66), .ZN(n415) );
  NAND2_X1 U465 ( .A1(n588), .A2(n565), .ZN(n611) );
  XNOR2_X1 U466 ( .A(n379), .B(n378), .ZN(G51) );
  INV_X1 U467 ( .A(KEYINPUT56), .ZN(n378) );
  NAND2_X1 U468 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U469 ( .A(n382), .B(n355), .ZN(n381) );
  XNOR2_X1 U470 ( .A(n666), .B(n368), .ZN(G75) );
  XNOR2_X1 U471 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n368) );
  NOR2_X1 U472 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U473 ( .A(n515), .B(n500), .ZN(n568) );
  AND2_X1 U474 ( .A1(n388), .A2(n387), .ZN(n345) );
  XOR2_X1 U475 ( .A(n423), .B(KEYINPUT88), .Z(n346) );
  AND2_X1 U476 ( .A1(n591), .A2(n419), .ZN(n347) );
  XOR2_X1 U477 ( .A(G125), .B(G140), .Z(n348) );
  XOR2_X1 U478 ( .A(n449), .B(n448), .Z(n349) );
  XNOR2_X1 U479 ( .A(n511), .B(KEYINPUT19), .ZN(n555) );
  INV_X1 U480 ( .A(n558), .ZN(n581) );
  XOR2_X1 U481 ( .A(n561), .B(KEYINPUT79), .Z(n350) );
  XOR2_X1 U482 ( .A(n503), .B(n502), .Z(n351) );
  AND2_X1 U483 ( .A1(G214), .A2(n494), .ZN(n352) );
  AND2_X1 U484 ( .A1(n389), .A2(n390), .ZN(n353) );
  BUF_X1 U485 ( .A(n569), .Z(n640) );
  XOR2_X1 U486 ( .A(KEYINPUT45), .B(KEYINPUT85), .Z(n354) );
  XOR2_X1 U487 ( .A(n431), .B(n430), .Z(n355) );
  XNOR2_X1 U488 ( .A(n375), .B(n372), .ZN(n501) );
  NOR2_X1 U489 ( .A1(n716), .A2(G952), .ZN(n689) );
  INV_X1 U490 ( .A(n689), .ZN(n380) );
  XOR2_X1 U491 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n356) );
  XOR2_X1 U492 ( .A(n603), .B(KEYINPUT63), .Z(n357) );
  XNOR2_X1 U493 ( .A(G902), .B(KEYINPUT15), .ZN(n596) );
  NAND2_X1 U494 ( .A1(n690), .A2(n715), .ZN(n358) );
  XNOR2_X1 U495 ( .A(n360), .B(n359), .ZN(n542) );
  AND2_X1 U496 ( .A1(n526), .A2(n527), .ZN(n360) );
  NAND2_X1 U497 ( .A1(n362), .A2(n392), .ZN(n384) );
  NAND2_X1 U498 ( .A1(n353), .A2(n385), .ZN(n362) );
  INV_X1 U499 ( .A(n674), .ZN(n410) );
  NAND2_X1 U500 ( .A1(n674), .A2(n675), .ZN(n679) );
  XNOR2_X1 U501 ( .A(n363), .B(n356), .ZN(G60) );
  NAND2_X1 U502 ( .A1(n680), .A2(n380), .ZN(n363) );
  AND2_X1 U503 ( .A1(n365), .A2(n416), .ZN(n397) );
  NOR2_X1 U504 ( .A1(n541), .A2(n542), .ZN(n365) );
  XNOR2_X1 U505 ( .A(n366), .B(n357), .ZN(G57) );
  NAND2_X1 U506 ( .A1(n602), .A2(n380), .ZN(n366) );
  XNOR2_X2 U507 ( .A(n367), .B(n487), .ZN(n564) );
  NAND2_X1 U508 ( .A1(n482), .A2(G221), .ZN(n483) );
  AND2_X1 U509 ( .A1(n370), .A2(n640), .ZN(n588) );
  NAND2_X1 U510 ( .A1(n370), .A2(n350), .ZN(n369) );
  NAND2_X1 U511 ( .A1(n681), .A2(G210), .ZN(n382) );
  NAND2_X1 U512 ( .A1(n384), .A2(n383), .ZN(n572) );
  NAND2_X1 U513 ( .A1(n345), .A2(n353), .ZN(n383) );
  NAND2_X1 U514 ( .A1(n568), .A2(n391), .ZN(n390) );
  NAND2_X1 U515 ( .A1(n353), .A2(n388), .ZN(n661) );
  NOR2_X1 U516 ( .A1(n581), .A2(n392), .ZN(n387) );
  NAND2_X1 U517 ( .A1(n570), .A2(n391), .ZN(n389) );
  XNOR2_X2 U518 ( .A(n394), .B(n393), .ZN(n515) );
  XNOR2_X1 U519 ( .A(n397), .B(KEYINPUT48), .ZN(n396) );
  NOR2_X1 U520 ( .A1(n723), .A2(n724), .ZN(n540) );
  XNOR2_X2 U521 ( .A(n403), .B(n351), .ZN(n548) );
  NAND2_X1 U522 ( .A1(n406), .A2(n405), .ZN(n404) );
  AND2_X1 U523 ( .A1(n673), .A2(n594), .ZN(n409) );
  NAND2_X1 U524 ( .A1(n410), .A2(n660), .ZN(n664) );
  NOR2_X1 U525 ( .A1(n624), .A2(n417), .ZN(n416) );
  AND2_X1 U526 ( .A1(n514), .A2(n513), .ZN(n417) );
  NOR2_X1 U527 ( .A1(n628), .A2(n550), .ZN(n418) );
  AND2_X1 U528 ( .A1(n590), .A2(n604), .ZN(n419) );
  XOR2_X1 U529 ( .A(KEYINPUT36), .B(n505), .Z(n420) );
  INV_X1 U530 ( .A(KEYINPUT46), .ZN(n539) );
  INV_X1 U531 ( .A(n433), .ZN(n422) );
  AND2_X1 U532 ( .A1(n720), .A2(KEYINPUT67), .ZN(n578) );
  XNOR2_X1 U533 ( .A(n496), .B(n495), .ZN(n497) );
  INV_X1 U534 ( .A(n626), .ZN(n550) );
  INV_X1 U535 ( .A(n447), .ZN(n429) );
  INV_X1 U536 ( .A(KEYINPUT62), .ZN(n598) );
  INV_X1 U537 ( .A(KEYINPUT89), .ZN(n502) );
  XNOR2_X1 U538 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n431) );
  XNOR2_X1 U539 ( .A(G125), .B(KEYINPUT17), .ZN(n423) );
  XNOR2_X2 U540 ( .A(KEYINPUT64), .B(n691), .ZN(n716) );
  NAND2_X1 U541 ( .A1(G224), .A2(n716), .ZN(n424) );
  XNOR2_X1 U542 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U543 ( .A(G119), .B(KEYINPUT3), .Z(n428) );
  XNOR2_X1 U544 ( .A(G116), .B(G113), .ZN(n427) );
  XNOR2_X1 U545 ( .A(n501), .B(KEYINPUT81), .ZN(n430) );
  XNOR2_X1 U546 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U547 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U548 ( .A1(G227), .A2(n716), .ZN(n440) );
  XNOR2_X1 U549 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U550 ( .A(n498), .B(n442), .ZN(n667) );
  XNOR2_X1 U551 ( .A(KEYINPUT70), .B(G469), .ZN(n443) );
  XNOR2_X2 U552 ( .A(n444), .B(n443), .ZN(n518) );
  XNOR2_X1 U553 ( .A(n446), .B(n445), .ZN(n452) );
  XOR2_X1 U554 ( .A(n447), .B(KEYINPUT11), .Z(n448) );
  XNOR2_X1 U555 ( .A(KEYINPUT10), .B(n348), .ZN(n709) );
  XNOR2_X1 U556 ( .A(G146), .B(n709), .ZN(n478) );
  XNOR2_X1 U557 ( .A(n349), .B(n478), .ZN(n451) );
  XNOR2_X1 U558 ( .A(n450), .B(KEYINPUT72), .ZN(n494) );
  NOR2_X1 U559 ( .A1(G902), .A2(n677), .ZN(n455) );
  XNOR2_X1 U560 ( .A(KEYINPUT13), .B(KEYINPUT99), .ZN(n453) );
  XOR2_X1 U561 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n457) );
  XNOR2_X1 U562 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U563 ( .A(n459), .B(n458), .ZN(n465) );
  XOR2_X1 U564 ( .A(G122), .B(KEYINPUT7), .Z(n463) );
  NAND2_X1 U565 ( .A1(G234), .A2(n716), .ZN(n460) );
  NAND2_X1 U566 ( .A1(G217), .A2(n482), .ZN(n462) );
  XNOR2_X1 U567 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U568 ( .A(n465), .B(n464), .ZN(n683) );
  NOR2_X1 U569 ( .A1(G902), .A2(n683), .ZN(n466) );
  XNOR2_X1 U570 ( .A(G478), .B(n466), .ZN(n528) );
  INV_X1 U571 ( .A(n528), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n529), .A2(n512), .ZN(n467) );
  XOR2_X1 U573 ( .A(KEYINPUT21), .B(KEYINPUT94), .Z(n470) );
  NAND2_X1 U574 ( .A1(G234), .A2(n596), .ZN(n468) );
  XNOR2_X1 U575 ( .A(KEYINPUT20), .B(n468), .ZN(n471) );
  NAND2_X1 U576 ( .A1(n471), .A2(G221), .ZN(n469) );
  XOR2_X1 U577 ( .A(n470), .B(n469), .Z(n643) );
  INV_X1 U578 ( .A(n643), .ZN(n556) );
  XOR2_X1 U579 ( .A(KEYINPUT74), .B(KEYINPUT25), .Z(n473) );
  NAND2_X1 U580 ( .A1(n471), .A2(G217), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U582 ( .A(KEYINPUT93), .B(n474), .ZN(n487) );
  XOR2_X1 U583 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n476) );
  XNOR2_X1 U584 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U585 ( .A(n478), .B(n477), .ZN(n486) );
  XOR2_X1 U586 ( .A(KEYINPUT24), .B(KEYINPUT83), .Z(n480) );
  XNOR2_X1 U587 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U588 ( .A(KEYINPUT91), .B(n481), .Z(n484) );
  NAND2_X1 U589 ( .A1(G234), .A2(G237), .ZN(n488) );
  XOR2_X1 U590 ( .A(n488), .B(KEYINPUT14), .Z(n657) );
  INV_X1 U591 ( .A(n657), .ZN(n492) );
  NOR2_X1 U592 ( .A1(n716), .A2(G900), .ZN(n489) );
  NAND2_X1 U593 ( .A1(G902), .A2(n489), .ZN(n490) );
  NAND2_X1 U594 ( .A1(G952), .A2(n691), .ZN(n551) );
  NAND2_X1 U595 ( .A1(n490), .A2(n551), .ZN(n491) );
  NAND2_X1 U596 ( .A1(n492), .A2(n491), .ZN(n517) );
  NOR2_X1 U597 ( .A1(n564), .A2(n517), .ZN(n493) );
  NAND2_X1 U598 ( .A1(n556), .A2(n493), .ZN(n506) );
  NAND2_X1 U599 ( .A1(n494), .A2(G210), .ZN(n499) );
  XOR2_X1 U600 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n495) );
  INV_X1 U601 ( .A(KEYINPUT6), .ZN(n500) );
  INV_X1 U602 ( .A(n596), .ZN(n673) );
  NAND2_X1 U603 ( .A1(G210), .A2(n504), .ZN(n503) );
  NAND2_X1 U604 ( .A1(G214), .A2(n504), .ZN(n629) );
  NAND2_X1 U605 ( .A1(n548), .A2(n629), .ZN(n511) );
  NOR2_X1 U606 ( .A1(n543), .A2(n511), .ZN(n505) );
  NOR2_X1 U607 ( .A1(n640), .A2(n420), .ZN(n624) );
  XOR2_X1 U608 ( .A(KEYINPUT47), .B(KEYINPUT68), .Z(n514) );
  NOR2_X1 U609 ( .A1(n506), .A2(n515), .ZN(n508) );
  XNOR2_X1 U610 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n507) );
  XNOR2_X1 U611 ( .A(n508), .B(n507), .ZN(n510) );
  XNOR2_X1 U612 ( .A(KEYINPUT108), .B(n518), .ZN(n509) );
  NOR2_X1 U613 ( .A1(n510), .A2(n509), .ZN(n533) );
  NAND2_X1 U614 ( .A1(n533), .A2(n555), .ZN(n616) );
  NAND2_X1 U615 ( .A1(n529), .A2(n512), .ZN(n622) );
  NOR2_X1 U616 ( .A1(n616), .A2(n634), .ZN(n513) );
  NAND2_X1 U617 ( .A1(n616), .A2(KEYINPUT47), .ZN(n527) );
  NAND2_X1 U618 ( .A1(n634), .A2(KEYINPUT47), .ZN(n524) );
  INV_X2 U619 ( .A(n515), .ZN(n646) );
  NAND2_X1 U620 ( .A1(n646), .A2(n629), .ZN(n516) );
  XNOR2_X1 U621 ( .A(n516), .B(KEYINPUT30), .ZN(n521) );
  INV_X1 U622 ( .A(n517), .ZN(n519) );
  NAND2_X1 U623 ( .A1(n519), .A2(n583), .ZN(n520) );
  NOR2_X1 U624 ( .A1(n528), .A2(n529), .ZN(n571) );
  INV_X1 U625 ( .A(n571), .ZN(n522) );
  NOR2_X1 U626 ( .A1(n536), .A2(n522), .ZN(n523) );
  NAND2_X1 U627 ( .A1(n548), .A2(n523), .ZN(n615) );
  NAND2_X1 U628 ( .A1(n524), .A2(n615), .ZN(n525) );
  XOR2_X1 U629 ( .A(KEYINPUT80), .B(n525), .Z(n526) );
  NAND2_X1 U630 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U631 ( .A(n530), .B(KEYINPUT102), .ZN(n632) );
  NAND2_X1 U632 ( .A1(n630), .A2(n629), .ZN(n633) );
  NOR2_X1 U633 ( .A1(n632), .A2(n633), .ZN(n532) );
  XNOR2_X1 U634 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n531) );
  XNOR2_X1 U635 ( .A(n532), .B(n531), .ZN(n662) );
  INV_X1 U636 ( .A(n533), .ZN(n534) );
  INV_X1 U637 ( .A(n630), .ZN(n535) );
  XNOR2_X1 U638 ( .A(n537), .B(KEYINPUT39), .ZN(n549) );
  NOR2_X1 U639 ( .A1(n549), .A2(n619), .ZN(n538) );
  XNOR2_X1 U640 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U641 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n546) );
  INV_X1 U642 ( .A(n640), .ZN(n563) );
  NOR2_X1 U643 ( .A1(n563), .A2(n543), .ZN(n544) );
  NAND2_X1 U644 ( .A1(n544), .A2(n629), .ZN(n545) );
  XOR2_X1 U645 ( .A(n546), .B(n545), .Z(n547) );
  NOR2_X1 U646 ( .A1(n548), .A2(n547), .ZN(n628) );
  OR2_X1 U647 ( .A1(n549), .A2(n622), .ZN(n626) );
  XNOR2_X1 U648 ( .A(KEYINPUT90), .B(G898), .ZN(n693) );
  NOR2_X1 U649 ( .A1(n691), .A2(n693), .ZN(n702) );
  NAND2_X1 U650 ( .A1(n702), .A2(G902), .ZN(n552) );
  AND2_X1 U651 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U652 ( .A1(n553), .A2(n657), .ZN(n554) );
  NOR2_X1 U653 ( .A1(n632), .A2(n643), .ZN(n557) );
  NAND2_X1 U654 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U655 ( .A(n564), .B(KEYINPUT103), .ZN(n642) );
  NAND2_X1 U656 ( .A1(n568), .A2(n642), .ZN(n560) );
  NOR2_X1 U657 ( .A1(n640), .A2(n560), .ZN(n561) );
  XOR2_X1 U658 ( .A(KEYINPUT78), .B(KEYINPUT32), .Z(n562) );
  NOR2_X1 U659 ( .A1(n564), .A2(n646), .ZN(n565) );
  INV_X1 U660 ( .A(n568), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U662 ( .A1(n720), .A2(KEYINPUT67), .ZN(n574) );
  NAND2_X1 U663 ( .A1(n577), .A2(n574), .ZN(n576) );
  NAND2_X1 U664 ( .A1(n578), .A2(n577), .ZN(n591) );
  NAND2_X1 U665 ( .A1(n646), .A2(n579), .ZN(n649) );
  NOR2_X1 U666 ( .A1(n581), .A2(n649), .ZN(n580) );
  XNOR2_X1 U667 ( .A(KEYINPUT31), .B(n580), .ZN(n621) );
  NOR2_X1 U668 ( .A1(n646), .A2(n581), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n583), .A2(n582), .ZN(n607) );
  NAND2_X1 U670 ( .A1(n621), .A2(n607), .ZN(n584) );
  XNOR2_X1 U671 ( .A(n584), .B(KEYINPUT96), .ZN(n586) );
  NAND2_X1 U672 ( .A1(n586), .A2(n585), .ZN(n590) );
  NOR2_X1 U673 ( .A1(n587), .A2(n642), .ZN(n589) );
  NAND2_X1 U674 ( .A1(n589), .A2(n588), .ZN(n604) );
  INV_X1 U675 ( .A(KEYINPUT2), .ZN(n593) );
  NOR2_X1 U676 ( .A1(KEYINPUT73), .A2(n593), .ZN(n592) );
  NAND2_X1 U677 ( .A1(KEYINPUT73), .A2(n593), .ZN(n594) );
  AND2_X1 U678 ( .A1(n673), .A2(G472), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n674), .A2(n597), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U681 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U682 ( .A(KEYINPUT87), .B(KEYINPUT112), .ZN(n603) );
  XNOR2_X1 U683 ( .A(G101), .B(n604), .ZN(G3) );
  NOR2_X1 U684 ( .A1(n619), .A2(n607), .ZN(n606) );
  XNOR2_X1 U685 ( .A(G104), .B(KEYINPUT113), .ZN(n605) );
  XNOR2_X1 U686 ( .A(n606), .B(n605), .ZN(G6) );
  NOR2_X1 U687 ( .A1(n622), .A2(n607), .ZN(n609) );
  XNOR2_X1 U688 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U690 ( .A(G107), .B(n610), .ZN(G9) );
  XNOR2_X1 U691 ( .A(G110), .B(n611), .ZN(G12) );
  NOR2_X1 U692 ( .A1(n622), .A2(n616), .ZN(n613) );
  XNOR2_X1 U693 ( .A(KEYINPUT114), .B(KEYINPUT29), .ZN(n612) );
  XNOR2_X1 U694 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U695 ( .A(G128), .B(n614), .ZN(G30) );
  XNOR2_X1 U696 ( .A(G143), .B(n615), .ZN(G45) );
  NOR2_X1 U697 ( .A1(n619), .A2(n616), .ZN(n618) );
  XNOR2_X1 U698 ( .A(G146), .B(KEYINPUT115), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n618), .B(n617), .ZN(G48) );
  NOR2_X1 U700 ( .A1(n619), .A2(n621), .ZN(n620) );
  XOR2_X1 U701 ( .A(G113), .B(n620), .Z(G15) );
  NOR2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U703 ( .A(G116), .B(n623), .Z(G18) );
  XNOR2_X1 U704 ( .A(G125), .B(n624), .ZN(n625) );
  XNOR2_X1 U705 ( .A(n625), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U706 ( .A(G134), .B(KEYINPUT116), .ZN(n627) );
  XNOR2_X1 U707 ( .A(n627), .B(n626), .ZN(G36) );
  XOR2_X1 U708 ( .A(G140), .B(n628), .Z(G42) );
  NOR2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n636) );
  NOR2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT117), .B(n637), .Z(n638) );
  NOR2_X1 U714 ( .A1(n661), .A2(n638), .ZN(n654) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n641), .B(KEYINPUT50), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U718 ( .A(KEYINPUT49), .B(n644), .ZN(n645) );
  NOR2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT51), .B(n651), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n662), .A2(n652), .ZN(n653) );
  NOR2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U725 ( .A(n655), .B(KEYINPUT52), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n656), .B(KEYINPUT118), .ZN(n658) );
  NOR2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U728 ( .A1(G952), .A2(n659), .ZN(n660) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n691), .A2(n665), .ZN(n666) );
  XNOR2_X1 U731 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n669) );
  XNOR2_X1 U732 ( .A(n667), .B(KEYINPUT57), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n669), .B(n668), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n681), .A2(G469), .ZN(n670) );
  XOR2_X1 U735 ( .A(n671), .B(n670), .Z(n672) );
  NOR2_X1 U736 ( .A1(n689), .A2(n672), .ZN(G54) );
  AND2_X1 U737 ( .A1(n673), .A2(G475), .ZN(n675) );
  XOR2_X1 U738 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n676) );
  XNOR2_X1 U739 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U740 ( .A1(G478), .A2(n685), .ZN(n682) );
  XNOR2_X1 U741 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U742 ( .A1(n689), .A2(n684), .ZN(G63) );
  NAND2_X1 U743 ( .A1(G217), .A2(n685), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n689), .A2(n688), .ZN(G66) );
  NAND2_X1 U746 ( .A1(n691), .A2(n690), .ZN(n697) );
  NAND2_X1 U747 ( .A1(G953), .A2(G224), .ZN(n692) );
  XNOR2_X1 U748 ( .A(n692), .B(KEYINPUT61), .ZN(n694) );
  NAND2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U750 ( .A(KEYINPUT123), .B(n695), .Z(n696) );
  NAND2_X1 U751 ( .A1(n697), .A2(n696), .ZN(n704) );
  XOR2_X1 U752 ( .A(G101), .B(n698), .Z(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n704), .B(n703), .ZN(G69) );
  XNOR2_X1 U756 ( .A(G227), .B(KEYINPUT126), .ZN(n711) );
  XNOR2_X1 U757 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n708) );
  XNOR2_X1 U758 ( .A(n705), .B(n706), .ZN(n707) );
  XNOR2_X1 U759 ( .A(n708), .B(n707), .ZN(n710) );
  XNOR2_X1 U760 ( .A(n709), .B(n710), .ZN(n714) );
  XOR2_X1 U761 ( .A(n711), .B(n714), .Z(n712) );
  NAND2_X1 U762 ( .A1(n712), .A2(G900), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n713), .A2(G953), .ZN(n719) );
  XNOR2_X1 U764 ( .A(n715), .B(n714), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U766 ( .A1(n719), .A2(n718), .ZN(G72) );
  XNOR2_X1 U767 ( .A(n720), .B(G122), .ZN(n721) );
  XNOR2_X1 U768 ( .A(n721), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U769 ( .A(n722), .B(G119), .ZN(G21) );
  XOR2_X1 U770 ( .A(n723), .B(G131), .Z(G33) );
  XOR2_X1 U771 ( .A(G137), .B(n724), .Z(G39) );
endmodule

