

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U552 ( .A(n690), .B(KEYINPUT98), .ZN(n692) );
  NOR2_X1 U553 ( .A1(G651), .A2(n581), .ZN(n786) );
  NOR2_X1 U554 ( .A1(n680), .A2(n679), .ZN(n515) );
  INV_X1 U555 ( .A(KEYINPUT93), .ZN(n630) );
  XNOR2_X1 U556 ( .A(n630), .B(KEYINPUT27), .ZN(n631) );
  XNOR2_X1 U557 ( .A(n632), .B(n631), .ZN(n635) );
  AND2_X1 U558 ( .A1(n654), .A2(n653), .ZN(n657) );
  INV_X1 U559 ( .A(KEYINPUT97), .ZN(n662) );
  NOR2_X1 U560 ( .A1(G2084), .A2(n649), .ZN(n668) );
  INV_X1 U561 ( .A(n705), .ZN(n597) );
  NAND2_X1 U562 ( .A1(n706), .A2(n597), .ZN(n649) );
  INV_X1 U563 ( .A(n1014), .ZN(n691) );
  AND2_X1 U564 ( .A1(n692), .A2(n691), .ZN(n697) );
  AND2_X1 U565 ( .A1(n550), .A2(G2104), .ZN(n889) );
  NOR2_X2 U566 ( .A1(G2104), .A2(n550), .ZN(n896) );
  XOR2_X1 U567 ( .A(KEYINPUT15), .B(n622), .Z(n997) );
  XNOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .ZN(n516) );
  XOR2_X1 U569 ( .A(n516), .B(KEYINPUT68), .Z(n581) );
  NAND2_X1 U570 ( .A1(n786), .A2(G51), .ZN(n520) );
  INV_X1 U571 ( .A(G651), .ZN(n524) );
  NOR2_X1 U572 ( .A1(G543), .A2(n524), .ZN(n517) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n517), .Z(n518) );
  XNOR2_X1 U574 ( .A(KEYINPUT70), .B(n518), .ZN(n788) );
  NAND2_X1 U575 ( .A1(G63), .A2(n788), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U577 ( .A(KEYINPUT6), .B(n521), .ZN(n530) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n791) );
  NAND2_X1 U579 ( .A1(G89), .A2(n791), .ZN(n522) );
  XNOR2_X1 U580 ( .A(n522), .B(KEYINPUT4), .ZN(n523) );
  XNOR2_X1 U581 ( .A(n523), .B(KEYINPUT76), .ZN(n527) );
  OR2_X1 U582 ( .A1(n524), .A2(n581), .ZN(n525) );
  XNOR2_X2 U583 ( .A(KEYINPUT69), .B(n525), .ZN(n792) );
  NAND2_X1 U584 ( .A1(G76), .A2(n792), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U586 ( .A(n528), .B(KEYINPUT5), .Z(n529) );
  NOR2_X1 U587 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U588 ( .A(KEYINPUT77), .B(n531), .Z(n532) );
  XOR2_X1 U589 ( .A(KEYINPUT7), .B(n532), .Z(G168) );
  XOR2_X1 U590 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U591 ( .A1(n786), .A2(G52), .ZN(n533) );
  XNOR2_X1 U592 ( .A(KEYINPUT71), .B(n533), .ZN(n541) );
  NAND2_X1 U593 ( .A1(G90), .A2(n791), .ZN(n535) );
  NAND2_X1 U594 ( .A1(G77), .A2(n792), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U596 ( .A(n536), .B(KEYINPUT72), .ZN(n537) );
  XNOR2_X1 U597 ( .A(n537), .B(KEYINPUT9), .ZN(n539) );
  NAND2_X1 U598 ( .A1(G64), .A2(n788), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U600 ( .A1(n541), .A2(n540), .ZN(G171) );
  INV_X1 U601 ( .A(G171), .ZN(G301) );
  NAND2_X1 U602 ( .A1(n792), .A2(G72), .ZN(n543) );
  NAND2_X1 U603 ( .A1(G60), .A2(n788), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G85), .A2(n791), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G47), .A2(n786), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n546) );
  OR2_X1 U608 ( .A1(n547), .A2(n546), .ZN(G290) );
  INV_X1 U609 ( .A(G2105), .ZN(n550) );
  NAND2_X1 U610 ( .A1(G101), .A2(n889), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n548), .B(KEYINPUT23), .ZN(n549) );
  XOR2_X1 U612 ( .A(n549), .B(KEYINPUT64), .Z(n594) );
  NAND2_X1 U613 ( .A1(G125), .A2(n896), .ZN(n558) );
  XNOR2_X1 U614 ( .A(KEYINPUT66), .B(KEYINPUT17), .ZN(n552) );
  NOR2_X1 U615 ( .A1(G2105), .A2(G2104), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(KEYINPUT65), .B(n553), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n559), .A2(G137), .ZN(n555) );
  AND2_X1 U619 ( .A1(G2105), .A2(G2104), .ZN(n895) );
  NAND2_X1 U620 ( .A1(G113), .A2(n895), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT67), .ZN(n557) );
  AND2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n595) );
  AND2_X1 U624 ( .A1(n594), .A2(n595), .ZN(G160) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  INV_X1 U628 ( .A(G120), .ZN(G236) );
  INV_X1 U629 ( .A(G69), .ZN(G235) );
  INV_X1 U630 ( .A(G108), .ZN(G238) );
  NAND2_X1 U631 ( .A1(G138), .A2(n559), .ZN(n562) );
  NAND2_X1 U632 ( .A1(G126), .A2(n896), .ZN(n560) );
  XOR2_X1 U633 ( .A(KEYINPUT83), .B(n560), .Z(n561) );
  NAND2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U635 ( .A1(G114), .A2(n895), .ZN(n564) );
  NAND2_X1 U636 ( .A1(G102), .A2(n889), .ZN(n563) );
  NAND2_X1 U637 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U638 ( .A1(n566), .A2(n565), .ZN(G164) );
  NAND2_X1 U639 ( .A1(G88), .A2(n791), .ZN(n568) );
  NAND2_X1 U640 ( .A1(G62), .A2(n788), .ZN(n567) );
  NAND2_X1 U641 ( .A1(n568), .A2(n567), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G75), .A2(n792), .ZN(n569) );
  XOR2_X1 U643 ( .A(KEYINPUT81), .B(n569), .Z(n571) );
  NAND2_X1 U644 ( .A1(n786), .A2(G50), .ZN(n570) );
  NAND2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U646 ( .A1(n573), .A2(n572), .ZN(G166) );
  INV_X1 U647 ( .A(G166), .ZN(G303) );
  NAND2_X1 U648 ( .A1(G91), .A2(n791), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G65), .A2(n788), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U651 ( .A1(G53), .A2(n786), .ZN(n576) );
  XNOR2_X1 U652 ( .A(KEYINPUT73), .B(n576), .ZN(n577) );
  NOR2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n792), .A2(G78), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(G299) );
  NAND2_X1 U656 ( .A1(G49), .A2(n786), .ZN(n583) );
  NAND2_X1 U657 ( .A1(G87), .A2(n581), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n584) );
  NOR2_X1 U659 ( .A1(n788), .A2(n584), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G651), .A2(G74), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(G288) );
  NAND2_X1 U662 ( .A1(G86), .A2(n791), .ZN(n588) );
  NAND2_X1 U663 ( .A1(G61), .A2(n788), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G73), .A2(n792), .ZN(n589) );
  XOR2_X1 U666 ( .A(KEYINPUT2), .B(n589), .Z(n590) );
  NOR2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n786), .A2(G48), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n593), .A2(n592), .ZN(G305) );
  NOR2_X1 U670 ( .A1(G164), .A2(G1384), .ZN(n706) );
  AND2_X1 U671 ( .A1(G40), .A2(n594), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n596), .A2(n595), .ZN(n705) );
  NAND2_X1 U673 ( .A1(G8), .A2(n649), .ZN(n704) );
  NOR2_X1 U674 ( .A1(G1971), .A2(n704), .ZN(n599) );
  NOR2_X1 U675 ( .A1(G2090), .A2(n649), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G303), .A2(n600), .ZN(n665) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n602) );
  NAND2_X1 U679 ( .A1(G56), .A2(n788), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n602), .B(n601), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n791), .A2(G81), .ZN(n603) );
  XNOR2_X1 U682 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U683 ( .A1(G68), .A2(n792), .ZN(n604) );
  NAND2_X1 U684 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U685 ( .A(KEYINPUT13), .B(n606), .Z(n607) );
  NOR2_X1 U686 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n786), .A2(G43), .ZN(n609) );
  NAND2_X1 U688 ( .A1(n610), .A2(n609), .ZN(n1007) );
  INV_X1 U689 ( .A(G1996), .ZN(n715) );
  NOR2_X1 U690 ( .A1(n649), .A2(n715), .ZN(n611) );
  XOR2_X1 U691 ( .A(n611), .B(KEYINPUT26), .Z(n613) );
  NAND2_X1 U692 ( .A1(n649), .A2(G1341), .ZN(n612) );
  NAND2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U694 ( .A1(n1007), .A2(n614), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n786), .A2(G54), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n792), .A2(G79), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G66), .A2(n788), .ZN(n615) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G92), .A2(n791), .ZN(n617) );
  XNOR2_X1 U700 ( .A(KEYINPUT75), .B(n617), .ZN(n618) );
  NOR2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G1348), .A2(n649), .ZN(n624) );
  INV_X1 U704 ( .A(n649), .ZN(n643) );
  NAND2_X1 U705 ( .A1(G2067), .A2(n643), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n627) );
  NOR2_X1 U707 ( .A1(n997), .A2(n627), .ZN(n625) );
  OR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n997), .A2(n627), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n637) );
  INV_X1 U711 ( .A(G299), .ZN(n802) );
  NAND2_X1 U712 ( .A1(n643), .A2(G2072), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G1956), .A2(n649), .ZN(n633) );
  XOR2_X1 U714 ( .A(KEYINPUT94), .B(n633), .Z(n634) );
  NOR2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n802), .A2(n638), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n641) );
  NOR2_X1 U718 ( .A1(n802), .A2(n638), .ZN(n639) );
  XOR2_X1 U719 ( .A(n639), .B(KEYINPUT28), .Z(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(KEYINPUT29), .ZN(n647) );
  XOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .Z(n929) );
  NOR2_X1 U723 ( .A1(n929), .A2(n649), .ZN(n645) );
  NOR2_X1 U724 ( .A1(n643), .A2(G1961), .ZN(n644) );
  NOR2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n655) );
  NOR2_X1 U726 ( .A1(G301), .A2(n655), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n704), .A2(G1966), .ZN(n648) );
  XNOR2_X1 U729 ( .A(n648), .B(KEYINPUT92), .ZN(n671) );
  XNOR2_X1 U730 ( .A(n668), .B(KEYINPUT91), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G8), .A2(n650), .ZN(n651) );
  NOR2_X1 U732 ( .A1(n671), .A2(n651), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n652), .B(KEYINPUT30), .ZN(n654) );
  INV_X1 U734 ( .A(G168), .ZN(n653) );
  AND2_X1 U735 ( .A1(G301), .A2(n655), .ZN(n656) );
  NOR2_X1 U736 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n658), .B(KEYINPUT31), .ZN(n659) );
  NOR2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT95), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n670), .A2(G286), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n666), .A2(G8), .ZN(n667) );
  XNOR2_X1 U744 ( .A(KEYINPUT32), .B(n667), .ZN(n698) );
  XOR2_X1 U745 ( .A(KEYINPUT91), .B(n668), .Z(n669) );
  NAND2_X1 U746 ( .A1(G8), .A2(n669), .ZN(n674) );
  INV_X1 U747 ( .A(n670), .ZN(n672) );
  NOR2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U750 ( .A(n675), .B(KEYINPUT96), .ZN(n699) );
  INV_X1 U751 ( .A(KEYINPUT33), .ZN(n676) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  AND2_X1 U753 ( .A1(n676), .A2(n1001), .ZN(n681) );
  AND2_X1 U754 ( .A1(n699), .A2(n681), .ZN(n677) );
  NAND2_X1 U755 ( .A1(n698), .A2(n677), .ZN(n689) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n683) );
  INV_X1 U757 ( .A(n704), .ZN(n679) );
  NAND2_X1 U758 ( .A1(n683), .A2(n679), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n678), .A2(KEYINPUT33), .ZN(n685) );
  INV_X1 U760 ( .A(n685), .ZN(n680) );
  INV_X1 U761 ( .A(n681), .ZN(n684) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U763 ( .A1(n683), .A2(n682), .ZN(n1002) );
  OR2_X1 U764 ( .A1(n684), .A2(n1002), .ZN(n686) );
  AND2_X1 U765 ( .A1(n686), .A2(n685), .ZN(n687) );
  OR2_X1 U766 ( .A1(n515), .A2(n687), .ZN(n688) );
  NAND2_X1 U767 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U768 ( .A(G1981), .B(G305), .ZN(n1014) );
  NOR2_X1 U769 ( .A1(G1981), .A2(G305), .ZN(n693) );
  XOR2_X1 U770 ( .A(n693), .B(KEYINPUT24), .Z(n694) );
  NOR2_X1 U771 ( .A1(n704), .A2(n694), .ZN(n695) );
  XNOR2_X1 U772 ( .A(n695), .B(KEYINPUT90), .ZN(n696) );
  NOR2_X1 U773 ( .A1(n697), .A2(n696), .ZN(n750) );
  NAND2_X1 U774 ( .A1(n699), .A2(n698), .ZN(n702) );
  NOR2_X1 U775 ( .A1(G2090), .A2(G303), .ZN(n700) );
  NAND2_X1 U776 ( .A1(G8), .A2(n700), .ZN(n701) );
  NAND2_X1 U777 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U778 ( .A1(n704), .A2(n703), .ZN(n748) );
  NOR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n755) );
  NAND2_X1 U780 ( .A1(G105), .A2(n889), .ZN(n707) );
  XNOR2_X1 U781 ( .A(n707), .B(KEYINPUT38), .ZN(n709) );
  BUF_X1 U782 ( .A(n559), .Z(n891) );
  NAND2_X1 U783 ( .A1(G141), .A2(n891), .ZN(n708) );
  NAND2_X1 U784 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U785 ( .A1(G117), .A2(n895), .ZN(n711) );
  NAND2_X1 U786 ( .A1(G129), .A2(n896), .ZN(n710) );
  NAND2_X1 U787 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U788 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U789 ( .A(KEYINPUT89), .B(n714), .Z(n869) );
  AND2_X1 U790 ( .A1(n715), .A2(n869), .ZN(n951) );
  NOR2_X1 U791 ( .A1(n869), .A2(n715), .ZN(n725) );
  NAND2_X1 U792 ( .A1(n895), .A2(G107), .ZN(n716) );
  XOR2_X1 U793 ( .A(KEYINPUT87), .B(n716), .Z(n718) );
  NAND2_X1 U794 ( .A1(n896), .A2(G119), .ZN(n717) );
  NAND2_X1 U795 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U796 ( .A(KEYINPUT88), .B(n719), .Z(n723) );
  NAND2_X1 U797 ( .A1(n891), .A2(G131), .ZN(n721) );
  NAND2_X1 U798 ( .A1(n889), .A2(G95), .ZN(n720) );
  AND2_X1 U799 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n870) );
  AND2_X1 U801 ( .A1(G1991), .A2(n870), .ZN(n724) );
  NOR2_X1 U802 ( .A1(n725), .A2(n724), .ZN(n947) );
  INV_X1 U803 ( .A(n755), .ZN(n726) );
  NOR2_X1 U804 ( .A1(n947), .A2(n726), .ZN(n751) );
  NOR2_X1 U805 ( .A1(G1986), .A2(G290), .ZN(n727) );
  NOR2_X1 U806 ( .A1(G1991), .A2(n870), .ZN(n945) );
  NOR2_X1 U807 ( .A1(n727), .A2(n945), .ZN(n728) );
  NOR2_X1 U808 ( .A1(n751), .A2(n728), .ZN(n729) );
  NOR2_X1 U809 ( .A1(n951), .A2(n729), .ZN(n730) );
  XNOR2_X1 U810 ( .A(n730), .B(KEYINPUT39), .ZN(n742) );
  XNOR2_X1 U811 ( .A(KEYINPUT37), .B(G2067), .ZN(n743) );
  NAND2_X1 U812 ( .A1(G116), .A2(n895), .ZN(n732) );
  NAND2_X1 U813 ( .A1(G128), .A2(n896), .ZN(n731) );
  NAND2_X1 U814 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U815 ( .A(n733), .B(KEYINPUT35), .ZN(n739) );
  NAND2_X1 U816 ( .A1(n889), .A2(G104), .ZN(n734) );
  XOR2_X1 U817 ( .A(KEYINPUT85), .B(n734), .Z(n736) );
  NAND2_X1 U818 ( .A1(G140), .A2(n891), .ZN(n735) );
  NAND2_X1 U819 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U820 ( .A(KEYINPUT34), .B(n737), .Z(n738) );
  NAND2_X1 U821 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U822 ( .A(n740), .B(KEYINPUT36), .Z(n903) );
  OR2_X1 U823 ( .A1(n743), .A2(n903), .ZN(n741) );
  XOR2_X1 U824 ( .A(KEYINPUT86), .B(n741), .Z(n954) );
  NAND2_X1 U825 ( .A1(n755), .A2(n954), .ZN(n752) );
  NAND2_X1 U826 ( .A1(n742), .A2(n752), .ZN(n744) );
  NAND2_X1 U827 ( .A1(n743), .A2(n903), .ZN(n958) );
  NAND2_X1 U828 ( .A1(n744), .A2(n958), .ZN(n745) );
  NAND2_X1 U829 ( .A1(n755), .A2(n745), .ZN(n746) );
  XNOR2_X1 U830 ( .A(n746), .B(KEYINPUT99), .ZN(n759) );
  INV_X1 U831 ( .A(n759), .ZN(n747) );
  AND2_X1 U832 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U833 ( .A1(n750), .A2(n749), .ZN(n761) );
  INV_X1 U834 ( .A(n751), .ZN(n753) );
  AND2_X1 U835 ( .A1(n753), .A2(n752), .ZN(n757) );
  XNOR2_X1 U836 ( .A(KEYINPUT84), .B(G1986), .ZN(n754) );
  XNOR2_X1 U837 ( .A(n754), .B(G290), .ZN(n1011) );
  NAND2_X1 U838 ( .A1(n755), .A2(n1011), .ZN(n756) );
  AND2_X1 U839 ( .A1(n757), .A2(n756), .ZN(n758) );
  OR2_X1 U840 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U841 ( .A1(n761), .A2(n760), .ZN(n763) );
  INV_X1 U842 ( .A(KEYINPUT40), .ZN(n762) );
  XNOR2_X1 U843 ( .A(n763), .B(n762), .ZN(G329) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U845 ( .A(n764), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U846 ( .A(G223), .ZN(n836) );
  NAND2_X1 U847 ( .A1(n836), .A2(G567), .ZN(n765) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n765), .Z(G234) );
  INV_X1 U849 ( .A(G860), .ZN(n799) );
  OR2_X1 U850 ( .A1(n1007), .A2(n799), .ZN(G153) );
  NAND2_X1 U851 ( .A1(G868), .A2(G301), .ZN(n767) );
  INV_X1 U852 ( .A(G868), .ZN(n768) );
  NAND2_X1 U853 ( .A1(n997), .A2(n768), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(G284) );
  NOR2_X1 U855 ( .A1(G286), .A2(n768), .ZN(n770) );
  NOR2_X1 U856 ( .A1(G868), .A2(G299), .ZN(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(G297) );
  NAND2_X1 U858 ( .A1(G559), .A2(n799), .ZN(n771) );
  XNOR2_X1 U859 ( .A(KEYINPUT78), .B(n771), .ZN(n772) );
  INV_X1 U860 ( .A(n997), .ZN(n797) );
  NAND2_X1 U861 ( .A1(n772), .A2(n797), .ZN(n773) );
  XNOR2_X1 U862 ( .A(KEYINPUT16), .B(n773), .ZN(G148) );
  NOR2_X1 U863 ( .A1(G868), .A2(n1007), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G868), .A2(n797), .ZN(n774) );
  NOR2_X1 U865 ( .A1(G559), .A2(n774), .ZN(n775) );
  NOR2_X1 U866 ( .A1(n776), .A2(n775), .ZN(G282) );
  NAND2_X1 U867 ( .A1(G123), .A2(n896), .ZN(n777) );
  XNOR2_X1 U868 ( .A(n777), .B(KEYINPUT18), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n895), .A2(G111), .ZN(n778) );
  NAND2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n889), .A2(G99), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G135), .A2(n891), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n944) );
  XNOR2_X1 U875 ( .A(G2096), .B(n944), .ZN(n785) );
  INV_X1 U876 ( .A(G2100), .ZN(n784) );
  NAND2_X1 U877 ( .A1(n785), .A2(n784), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G55), .A2(n786), .ZN(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT80), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G67), .A2(n788), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G93), .A2(n791), .ZN(n794) );
  NAND2_X1 U883 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U884 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n810) );
  NAND2_X1 U886 ( .A1(G559), .A2(n797), .ZN(n798) );
  XOR2_X1 U887 ( .A(n1007), .B(n798), .Z(n808) );
  NAND2_X1 U888 ( .A1(n799), .A2(n808), .ZN(n800) );
  XNOR2_X1 U889 ( .A(n800), .B(KEYINPUT79), .ZN(n801) );
  XNOR2_X1 U890 ( .A(n810), .B(n801), .ZN(G145) );
  XNOR2_X1 U891 ( .A(G166), .B(G305), .ZN(n807) );
  XNOR2_X1 U892 ( .A(n802), .B(n810), .ZN(n805) );
  XOR2_X1 U893 ( .A(KEYINPUT19), .B(G288), .Z(n803) );
  XNOR2_X1 U894 ( .A(G290), .B(n803), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n805), .B(n804), .ZN(n806) );
  XNOR2_X1 U896 ( .A(n807), .B(n806), .ZN(n909) );
  XNOR2_X1 U897 ( .A(n808), .B(n909), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n809), .A2(G868), .ZN(n812) );
  OR2_X1 U899 ( .A1(G868), .A2(n810), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n812), .A2(n811), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n813) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n813), .Z(n814) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n814), .ZN(n815) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n815), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n816), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U907 ( .A1(G235), .A2(G236), .ZN(n817) );
  XOR2_X1 U908 ( .A(KEYINPUT82), .B(n817), .Z(n818) );
  NOR2_X1 U909 ( .A1(G238), .A2(n818), .ZN(n819) );
  NAND2_X1 U910 ( .A1(G57), .A2(n819), .ZN(n919) );
  NAND2_X1 U911 ( .A1(n919), .A2(G567), .ZN(n824) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U914 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U915 ( .A1(G96), .A2(n822), .ZN(n920) );
  NAND2_X1 U916 ( .A1(n920), .A2(G2106), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n840) );
  NAND2_X1 U918 ( .A1(G483), .A2(G661), .ZN(n825) );
  NOR2_X1 U919 ( .A1(n840), .A2(n825), .ZN(n839) );
  NAND2_X1 U920 ( .A1(n839), .A2(G36), .ZN(G176) );
  XNOR2_X1 U921 ( .A(G2454), .B(G2451), .ZN(n834) );
  XNOR2_X1 U922 ( .A(G2430), .B(G2446), .ZN(n832) );
  XOR2_X1 U923 ( .A(G2435), .B(G2427), .Z(n827) );
  XNOR2_X1 U924 ( .A(KEYINPUT100), .B(G2438), .ZN(n826) );
  XNOR2_X1 U925 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U926 ( .A(n828), .B(G2443), .Z(n830) );
  XNOR2_X1 U927 ( .A(G1341), .B(G1348), .ZN(n829) );
  XNOR2_X1 U928 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U931 ( .A1(n835), .A2(G14), .ZN(n913) );
  XNOR2_X1 U932 ( .A(KEYINPUT101), .B(n913), .ZN(G401) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U935 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U938 ( .A(G96), .B(KEYINPUT102), .Z(G221) );
  INV_X1 U939 ( .A(n840), .ZN(G319) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2090), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n841), .B(KEYINPUT43), .ZN(n851) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2678), .Z(n843) );
  XNOR2_X1 U943 ( .A(KEYINPUT104), .B(G2096), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G2100), .B(G2084), .Z(n845) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2072), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U948 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT103), .B(KEYINPUT105), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U952 ( .A(G1956), .B(G1961), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1976), .B(G1966), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(G2474), .Z(n856) );
  XNOR2_X1 U956 ( .A(G1971), .B(G1986), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(KEYINPUT41), .B(G1981), .Z(n858) );
  XNOR2_X1 U959 ( .A(G1991), .B(G1996), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G100), .A2(n889), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n861), .B(KEYINPUT106), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G124), .A2(n896), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n862), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G112), .A2(n895), .ZN(n866) );
  NAND2_X1 U968 ( .A1(G136), .A2(n891), .ZN(n865) );
  NAND2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U970 ( .A1(n868), .A2(n867), .ZN(G162) );
  XOR2_X1 U971 ( .A(G162), .B(G164), .Z(n872) );
  XOR2_X1 U972 ( .A(n870), .B(n869), .Z(n871) );
  XNOR2_X1 U973 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U974 ( .A(KEYINPUT109), .B(KEYINPUT48), .Z(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(n876), .B(n875), .Z(n888) );
  NAND2_X1 U978 ( .A1(G118), .A2(n895), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G130), .A2(n896), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n885) );
  XNOR2_X1 U981 ( .A(KEYINPUT45), .B(KEYINPUT108), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n889), .A2(G106), .ZN(n881) );
  NAND2_X1 U983 ( .A1(G142), .A2(n891), .ZN(n879) );
  XOR2_X1 U984 ( .A(KEYINPUT107), .B(n879), .Z(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U986 ( .A(n883), .B(n882), .Z(n884) );
  NOR2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n944), .B(n886), .ZN(n887) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n902) );
  NAND2_X1 U990 ( .A1(n889), .A2(G103), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n890), .B(KEYINPUT110), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G139), .A2(n891), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(KEYINPUT111), .B(n894), .Z(n901) );
  NAND2_X1 U995 ( .A1(G115), .A2(n895), .ZN(n898) );
  NAND2_X1 U996 ( .A1(G127), .A2(n896), .ZN(n897) );
  NAND2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n899), .Z(n900) );
  NOR2_X1 U999 ( .A1(n901), .A2(n900), .ZN(n960) );
  XOR2_X1 U1000 ( .A(n902), .B(n960), .Z(n905) );
  XOR2_X1 U1001 ( .A(G160), .B(n903), .Z(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n906), .ZN(n907) );
  XOR2_X1 U1004 ( .A(KEYINPUT113), .B(n907), .Z(G395) );
  XNOR2_X1 U1005 ( .A(G286), .B(G301), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(n997), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n1007), .B(n909), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n912), .ZN(G397) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n913), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(G225) );
  XOR2_X1 U1016 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1019 ( .A(G325), .ZN(G261) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1021 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n939) );
  XNOR2_X1 U1022 ( .A(G2090), .B(G35), .ZN(n934) );
  XNOR2_X1 U1023 ( .A(G1996), .B(G32), .ZN(n922) );
  XNOR2_X1 U1024 ( .A(G33), .B(G2072), .ZN(n921) );
  NOR2_X1 U1025 ( .A1(n922), .A2(n921), .ZN(n928) );
  XOR2_X1 U1026 ( .A(G2067), .B(G26), .Z(n923) );
  NAND2_X1 U1027 ( .A1(n923), .A2(G28), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(G25), .B(G1991), .ZN(n924) );
  XNOR2_X1 U1029 ( .A(KEYINPUT118), .B(n924), .ZN(n925) );
  NOR2_X1 U1030 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n931) );
  XNOR2_X1 U1032 ( .A(G27), .B(n929), .ZN(n930) );
  NOR2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(KEYINPUT53), .B(n932), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1036 ( .A(G2084), .B(G34), .Z(n935) );
  XNOR2_X1 U1037 ( .A(KEYINPUT54), .B(n935), .ZN(n936) );
  NAND2_X1 U1038 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(n939), .B(n938), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(G29), .A2(n940), .ZN(n941) );
  XOR2_X1 U1041 ( .A(KEYINPUT120), .B(n941), .Z(n942) );
  NAND2_X1 U1042 ( .A1(n942), .A2(G11), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT121), .ZN(n973) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n949) );
  XOR2_X1 U1046 ( .A(G160), .B(G2084), .Z(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n956) );
  XOR2_X1 U1048 ( .A(G2090), .B(G162), .Z(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(n952), .B(KEYINPUT51), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(n957), .B(KEYINPUT115), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n967) );
  XNOR2_X1 U1055 ( .A(G2072), .B(n960), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G164), .B(G2078), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(n961), .B(KEYINPUT116), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1059 ( .A(KEYINPUT117), .B(n964), .Z(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT50), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT52), .B(n968), .ZN(n970) );
  INV_X1 U1063 ( .A(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n971), .A2(G29), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n1027) );
  XOR2_X1 U1067 ( .A(G1348), .B(KEYINPUT59), .Z(n974) );
  XNOR2_X1 U1068 ( .A(G4), .B(n974), .ZN(n981) );
  XOR2_X1 U1069 ( .A(G1981), .B(G6), .Z(n978) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G1956), .B(G20), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT125), .B(n979), .Z(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT60), .B(n982), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G21), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(G1961), .B(G5), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n994) );
  XNOR2_X1 U1081 ( .A(G1976), .B(G23), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G1986), .B(G24), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1084 ( .A(G1971), .B(KEYINPUT126), .Z(n989) );
  XNOR2_X1 U1085 ( .A(G22), .B(n989), .ZN(n990) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT58), .B(n992), .ZN(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1089 ( .A(KEYINPUT61), .B(n995), .Z(n996) );
  NOR2_X1 U1090 ( .A1(G16), .A2(n996), .ZN(n1024) );
  XOR2_X1 U1091 ( .A(G16), .B(KEYINPUT56), .Z(n1022) );
  XNOR2_X1 U1092 ( .A(G301), .B(G1961), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(n997), .B(G1348), .ZN(n998) );
  NOR2_X1 U1094 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(n1000), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1097 ( .A(G1956), .B(G299), .ZN(n1003) );
  NOR2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1099 ( .A1(n1006), .A2(n1005), .ZN(n1020) );
  NAND2_X1 U1100 ( .A1(G1971), .A2(G303), .ZN(n1009) );
  XOR2_X1 U1101 ( .A(G1341), .B(n1007), .Z(n1008) );
  NAND2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(G1966), .B(G168), .Z(n1012) );
  XNOR2_X1 U1105 ( .A(KEYINPUT122), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(KEYINPUT57), .B(KEYINPUT123), .ZN(n1015) );
  XNOR2_X1 U1108 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(n1025), .B(KEYINPUT127), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

