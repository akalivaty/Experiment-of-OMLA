//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  OR2_X1    g004(.A1(KEYINPUT70), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT70), .A2(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(G116), .A3(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT71), .ZN(new_n195));
  INV_X1    g009(.A(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT71), .A2(G116), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(G119), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n193), .A2(new_n199), .A3(KEYINPUT5), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n200), .A3(G113), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT2), .B(G113), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n193), .A3(new_n199), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G104), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G107), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n209), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n205), .A2(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n208), .A2(G104), .ZN(new_n214));
  OAI21_X1  g028(.A(G101), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n201), .A2(new_n204), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n193), .A2(new_n199), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n202), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n204), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(KEYINPUT72), .A3(new_n202), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT4), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n228), .A3(G101), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n218), .B1(new_n224), .B2(new_n230), .ZN(new_n231));
  XOR2_X1   g045(.A(G110), .B(G122), .Z(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n232), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n234), .B(new_n218), .C1(new_n224), .C2(new_n230), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(KEYINPUT6), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G953), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G224), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT79), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G125), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G146), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G146), .ZN(new_n250));
  AOI21_X1  g064(.A(G143), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n242), .B(new_n246), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n248), .A2(new_n250), .A3(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT66), .B1(new_n247), .B2(G143), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT64), .B(G146), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G143), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n243), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n248), .A2(new_n250), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n253), .B1(new_n265), .B2(new_n252), .ZN(new_n266));
  INV_X1    g080(.A(new_n246), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT65), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n241), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n253), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n270), .B1(new_n260), .B2(G143), .ZN(new_n271));
  XNOR2_X1  g085(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(G143), .B2(new_n260), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(new_n274), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n257), .B1(new_n260), .B2(G143), .ZN(new_n282));
  AND4_X1   g096(.A1(new_n261), .A2(new_n248), .A3(new_n250), .A4(G143), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n275), .A2(new_n241), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n240), .B1(new_n269), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n244), .B1(new_n282), .B2(new_n283), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n268), .A2(new_n288), .A3(new_n254), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G125), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n285), .A3(new_n239), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n231), .A2(new_n293), .A3(new_n232), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n236), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT80), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n285), .A4(new_n239), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT81), .B(KEYINPUT8), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n232), .B(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n201), .A2(new_n204), .A3(new_n217), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n217), .B1(new_n201), .B2(new_n204), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND3_X1   g117(.A1(new_n298), .A2(new_n235), .A3(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n239), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT82), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n290), .B2(new_n285), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n286), .A2(KEYINPUT82), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(G902), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n236), .A2(new_n292), .A3(KEYINPUT80), .A4(new_n294), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n190), .B1(new_n297), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n295), .A2(new_n296), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(new_n189), .A3(new_n313), .A4(new_n312), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n188), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT9), .B(G234), .ZN(new_n319));
  OAI21_X1  g133(.A(G221), .B1(new_n319), .B2(G902), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G469), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G140), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n237), .A2(G227), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT11), .ZN(new_n328));
  INV_X1    g142(.A(G134), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(G137), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(G137), .ZN(new_n331));
  INV_X1    g145(.A(G137), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT11), .A3(G134), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G131), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(G131), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n330), .A2(new_n333), .A3(new_n337), .A4(new_n331), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(G128), .B1(new_n253), .B2(new_n276), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n259), .A2(new_n262), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n272), .A2(G128), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n259), .B2(new_n262), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n217), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n275), .A2(new_n284), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n216), .A2(new_n346), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n345), .A2(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n264), .A2(new_n268), .A3(new_n229), .A4(new_n227), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n256), .A2(new_n280), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n265), .A2(new_n252), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n352), .A2(G128), .B1(new_n353), .B2(new_n270), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n348), .B1(new_n354), .B2(new_n344), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n259), .A2(new_n262), .A3(new_n341), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n216), .B1(new_n284), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n357), .B2(KEYINPUT10), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n289), .A2(new_n230), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n358), .A2(new_n359), .A3(new_n339), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n327), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n345), .A2(new_n346), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n350), .A2(new_n362), .A3(new_n340), .A4(new_n355), .ZN(new_n363));
  INV_X1    g177(.A(new_n327), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n275), .A2(new_n284), .A3(new_n216), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n345), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT12), .B1(new_n366), .B2(new_n339), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT12), .ZN(new_n368));
  AOI211_X1 g182(.A(new_n368), .B(new_n340), .C1(new_n345), .C2(new_n365), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n363), .B(new_n364), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(G902), .B1(new_n361), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n324), .B1(new_n371), .B2(new_n322), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n363), .B1(new_n367), .B2(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n327), .ZN(new_n374));
  INV_X1    g188(.A(new_n351), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n363), .A3(new_n364), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n376), .A3(G469), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n321), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n318), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(G234), .B2(new_n323), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n241), .A2(G140), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT16), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT16), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n382), .A3(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n386), .A3(new_n382), .A4(G125), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n385), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n247), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n385), .A2(new_n388), .A3(G146), .A4(new_n390), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(KEYINPUT70), .A2(G119), .ZN(new_n395));
  NOR2_X1   g209(.A1(KEYINPUT70), .A2(G119), .ZN(new_n396));
  OAI21_X1  g210(.A(G128), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G119), .A2(G128), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n397), .A2(KEYINPUT23), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n274), .B1(new_n395), .B2(new_n396), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT23), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G110), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n191), .A2(new_n192), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n398), .B1(new_n406), .B2(G128), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT24), .B(G110), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n394), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G110), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n400), .A2(new_n411), .A3(new_n403), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(new_n408), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n383), .A2(new_n384), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n260), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n393), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT22), .B(G137), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n237), .A2(G221), .A3(G234), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n410), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n410), .B2(new_n418), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT25), .B1(new_n424), .B2(new_n323), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n410), .A2(new_n418), .ZN(new_n426));
  INV_X1    g240(.A(new_n421), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n410), .A2(new_n418), .A3(new_n421), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n428), .A2(KEYINPUT25), .A3(new_n323), .A4(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n381), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT77), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n428), .A2(new_n323), .A3(new_n429), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT25), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n430), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT77), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n381), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n381), .A2(G902), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT78), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n424), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n433), .A2(new_n439), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n224), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT30), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(KEYINPUT69), .A2(KEYINPUT30), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n268), .A2(new_n288), .A3(new_n339), .A4(new_n254), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n334), .A2(G131), .ZN(new_n451));
  INV_X1    g265(.A(G131), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n332), .A2(G134), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n452), .B1(new_n453), .B2(new_n331), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n354), .B2(new_n344), .ZN(new_n456));
  AOI211_X1 g270(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n456), .ZN(new_n457));
  AND4_X1   g271(.A1(new_n446), .A2(new_n450), .A3(new_n456), .A4(new_n447), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n445), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n450), .A2(new_n224), .A3(new_n456), .ZN(new_n460));
  NOR2_X1   g274(.A1(G237), .A2(G953), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G210), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT27), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT26), .B(G101), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n459), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT31), .ZN(new_n467));
  INV_X1    g281(.A(new_n465), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT28), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n450), .A2(new_n456), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n445), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n471), .B2(new_n460), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n460), .A2(new_n469), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n468), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n466), .A2(new_n467), .A3(new_n475), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n450), .A2(new_n224), .A3(new_n456), .ZN(new_n477));
  INV_X1    g291(.A(new_n448), .ZN(new_n478));
  INV_X1    g292(.A(new_n449), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n450), .A2(new_n456), .A3(new_n446), .A4(new_n447), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n477), .B1(new_n482), .B2(new_n445), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT31), .A3(new_n465), .ZN(new_n484));
  NOR2_X1   g298(.A1(G472), .A2(G902), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT73), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n476), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT32), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT32), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n476), .A2(new_n489), .A3(new_n484), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n224), .B1(new_n450), .B2(new_n456), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT28), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n493), .A2(KEYINPUT29), .A3(new_n473), .A4(new_n465), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n494), .A2(KEYINPUT75), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(KEYINPUT75), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n323), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT74), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n493), .A2(new_n498), .A3(new_n473), .A4(new_n465), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT29), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n498), .B1(new_n483), .B2(new_n465), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n493), .A2(new_n473), .A3(new_n465), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G472), .B1(new_n497), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n444), .B1(new_n491), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT87), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n205), .ZN(new_n511));
  INV_X1    g325(.A(G237), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n237), .A3(G214), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT85), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n252), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n461), .B(G214), .C1(KEYINPUT85), .C2(G143), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G131), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n452), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n415), .B(KEYINPUT19), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n393), .B(new_n520), .C1(new_n522), .C2(new_n265), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n517), .B1(new_n524), .B2(new_n452), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n515), .A2(KEYINPUT18), .A3(new_n516), .A4(G131), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n415), .A2(new_n247), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n416), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n511), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n517), .A2(KEYINPUT17), .A3(G131), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n532), .A2(new_n392), .A3(KEYINPUT86), .A4(new_n393), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(new_n534), .A3(new_n519), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n392), .A3(new_n393), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT86), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n536), .A2(new_n539), .B1(new_n529), .B2(new_n527), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n531), .B1(new_n540), .B2(new_n511), .ZN(new_n541));
  OR2_X1    g355(.A1(G475), .A2(G902), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n507), .B(new_n509), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n523), .A2(new_n530), .ZN(new_n544));
  INV_X1    g358(.A(new_n511), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n537), .A2(new_n538), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n533), .A2(new_n535), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n511), .B(new_n530), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n542), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT87), .B1(new_n550), .B2(new_n508), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT20), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n543), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n540), .A2(new_n511), .ZN(new_n555));
  INV_X1    g369(.A(new_n549), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n323), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT15), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G478), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n197), .A2(G122), .A3(new_n198), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n196), .A2(G122), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n208), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n252), .A2(G128), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n274), .A2(G143), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G134), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n566), .A3(new_n329), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT14), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n562), .A2(new_n571), .A3(new_n563), .ZN(new_n572));
  OAI21_X1  g386(.A(G107), .B1(new_n562), .B2(new_n571), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n564), .B(new_n570), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n319), .A2(new_n380), .A3(G953), .ZN(new_n575));
  INV_X1    g389(.A(new_n564), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n208), .B1(new_n562), .B2(new_n563), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT13), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n566), .B1(new_n565), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT13), .B1(new_n252), .B2(G128), .ZN(new_n581));
  OAI21_X1  g395(.A(G134), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n569), .A2(KEYINPUT88), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT88), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n565), .A2(new_n566), .A3(new_n584), .A4(new_n329), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n574), .B(new_n575), .C1(new_n578), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT89), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n583), .A2(new_n585), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n589), .B(new_n582), .C1(new_n576), .C2(new_n577), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT89), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n574), .A4(new_n575), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n574), .B1(new_n578), .B2(new_n586), .ZN(new_n593));
  INV_X1    g407(.A(new_n575), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n588), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n323), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n561), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n596), .A2(KEYINPUT90), .A3(new_n323), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT90), .B1(new_n596), .B2(new_n323), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n560), .B(G478), .C1(new_n597), .C2(KEYINPUT91), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G952), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(G953), .ZN(new_n607));
  INV_X1    g421(.A(G234), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n607), .B1(new_n608), .B2(new_n512), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT92), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(G902), .B(G953), .C1(new_n608), .C2(new_n512), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT93), .Z(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT21), .B(G898), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n559), .A2(new_n605), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n379), .A2(new_n506), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT94), .B(G101), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G3));
  INV_X1    g434(.A(new_n616), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n318), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n487), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n476), .A2(KEYINPUT95), .A3(new_n323), .A4(new_n484), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n625), .A2(G472), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n476), .A2(new_n323), .A3(new_n484), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n624), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n361), .A2(new_n370), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n322), .A3(new_n323), .ZN(new_n632));
  INV_X1    g446(.A(new_n324), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n377), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n320), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n444), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n623), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n593), .B2(new_n594), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n596), .A2(new_n638), .B1(new_n587), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(G478), .A3(new_n323), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n600), .A2(new_n601), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(G478), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n559), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT34), .B(G104), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT96), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n645), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n550), .A2(new_n508), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n543), .A2(new_n551), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n605), .A2(new_n558), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n637), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT35), .B(G107), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  AND2_X1   g468(.A1(new_n554), .A2(new_n558), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n427), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT97), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n426), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n442), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n433), .A2(new_n439), .A3(new_n659), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n655), .A2(new_n604), .A3(new_n621), .A4(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n379), .A2(new_n630), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n491), .A2(new_n505), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n650), .A2(new_n558), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n611), .B1(new_n667), .B2(new_n614), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n666), .A2(new_n604), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n438), .B1(new_n437), .B2(new_n381), .ZN(new_n670));
  INV_X1    g484(.A(new_n381), .ZN(new_n671));
  AOI211_X1 g485(.A(KEYINPUT77), .B(new_n671), .C1(new_n436), .C2(new_n430), .ZN(new_n672));
  INV_X1    g486(.A(new_n659), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n635), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n665), .A2(new_n669), .A3(new_n675), .A4(new_n318), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT98), .B(G128), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G30));
  XNOR2_X1  g492(.A(new_n668), .B(KEYINPUT39), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n635), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT100), .Z(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n315), .A2(new_n317), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT38), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n468), .B1(new_n477), .B2(new_n492), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  INV_X1    g501(.A(new_n466), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n323), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G472), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n491), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n604), .B1(new_n554), .B2(new_n558), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n660), .A2(new_n188), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n685), .A2(new_n691), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n682), .A2(new_n683), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n252), .ZN(G45));
  INV_X1    g510(.A(new_n668), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n559), .A2(new_n643), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n665), .A2(new_n675), .A3(new_n699), .A4(new_n318), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NOR2_X1   g515(.A1(new_n622), .A2(new_n644), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n371), .A2(new_n322), .ZN(new_n703));
  AOI211_X1 g517(.A(G469), .B(G902), .C1(new_n361), .C2(new_n370), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n321), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n506), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NOR2_X1   g522(.A1(new_n622), .A2(new_n651), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n506), .A3(new_n705), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  AND3_X1   g525(.A1(new_n684), .A2(new_n705), .A3(new_n187), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n661), .A2(new_n712), .A3(new_n665), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n713), .A2(KEYINPUT101), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(KEYINPUT101), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  AND3_X1   g531(.A1(new_n692), .A2(new_n187), .A3(new_n684), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n433), .A2(new_n439), .A3(new_n443), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n627), .A2(G472), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(new_n487), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n703), .A2(new_n704), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n320), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n616), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n718), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND2_X1  g540(.A1(new_n698), .A2(KEYINPUT102), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT102), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n559), .A2(new_n643), .A3(new_n728), .A4(new_n697), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n720), .A2(new_n660), .A3(new_n487), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n712), .A2(new_n727), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n729), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n377), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n374), .A2(new_n376), .A3(KEYINPUT103), .A4(G469), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n372), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n321), .A2(new_n188), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n315), .A2(new_n317), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n734), .A2(KEYINPUT42), .A3(new_n506), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n506), .A2(new_n741), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n743), .B1(new_n744), .B2(new_n733), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NAND3_X1  g561(.A1(new_n506), .A2(new_n669), .A3(new_n741), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND2_X1  g563(.A1(new_n655), .A2(new_n643), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n630), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n660), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n374), .A2(new_n376), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n322), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n758), .B2(new_n757), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT46), .B1(new_n760), .B2(new_n633), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n704), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(KEYINPUT46), .A3(new_n633), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n321), .B(new_n679), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n754), .A2(new_n755), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n684), .A2(new_n188), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n756), .A2(new_n764), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT104), .B(G137), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G39));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n444), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n770), .A2(new_n665), .A3(new_n698), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT106), .ZN(new_n772));
  XNOR2_X1  g586(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n321), .B(new_n773), .C1(new_n762), .C2(new_n763), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n321), .B1(new_n762), .B2(new_n763), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n775), .B1(KEYINPUT105), .B2(new_n776), .ZN(new_n777));
  OR3_X1    g591(.A1(new_n772), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  XNOR2_X1  g593(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n780));
  INV_X1    g594(.A(new_n721), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n752), .A2(new_n611), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n752), .A2(KEYINPUT114), .A3(new_n611), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n685), .A2(new_n187), .A3(new_n723), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT116), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n722), .B(KEYINPUT107), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT115), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT115), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n321), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n796), .B1(new_n777), .B2(new_n774), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n766), .A3(new_n786), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n722), .A2(new_n315), .A3(new_n317), .A4(new_n739), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n784), .B2(new_n785), .ZN(new_n800));
  NOR4_X1   g614(.A1(new_n691), .A2(new_n799), .A3(new_n444), .A4(new_n610), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n559), .A2(new_n643), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n800), .A2(new_n730), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n790), .A2(KEYINPUT116), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n780), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n801), .A2(new_n559), .A3(new_n643), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n607), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n786), .B2(new_n712), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT48), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n800), .A2(new_n811), .A3(new_n506), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(new_n800), .B2(new_n506), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n790), .A2(new_n804), .A3(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n807), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n618), .A2(new_n662), .A3(new_n725), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n714), .B2(new_n715), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n741), .A2(new_n727), .A3(new_n730), .A4(new_n729), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n666), .A2(new_n605), .A3(new_n668), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n665), .A2(new_n675), .A3(new_n766), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n748), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n742), .B2(new_n745), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n644), .B1(new_n559), .B2(new_n604), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n623), .A2(new_n630), .A3(new_n636), .A4(new_n828), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n706), .A2(new_n710), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n822), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT108), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n320), .B1(new_n697), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n832), .B2(new_n697), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n433), .A2(new_n439), .A3(new_n659), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT109), .B1(new_n738), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n372), .A2(new_n736), .A3(new_n737), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n674), .A2(new_n837), .A3(new_n838), .A4(new_n834), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n718), .A2(new_n836), .A3(new_n691), .A4(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(new_n731), .A3(new_n676), .A4(new_n700), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n318), .A2(new_n378), .A3(new_n660), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n844), .B(new_n665), .C1(new_n669), .C2(new_n699), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT52), .A3(new_n731), .A4(new_n840), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n820), .B1(new_n831), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT110), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n822), .A2(new_n827), .A3(new_n830), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n843), .B2(new_n846), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n843), .A2(new_n846), .A3(new_n851), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n850), .B(KEYINPUT53), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT110), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n855), .B(new_n820), .C1(new_n831), .C2(new_n847), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n849), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT54), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n853), .A2(new_n852), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n820), .B1(new_n859), .B2(new_n831), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n843), .A2(new_n846), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(KEYINPUT111), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n843), .A2(new_n846), .A3(new_n851), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n831), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n863), .B(new_n861), .C1(new_n867), .C2(KEYINPUT53), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n858), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n819), .A2(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n792), .B(KEYINPUT49), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n719), .A2(new_n655), .A3(new_n643), .A4(new_n739), .ZN(new_n874));
  OR4_X1    g688(.A1(new_n691), .A2(new_n873), .A3(new_n685), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n872), .A2(new_n875), .ZN(G75));
  NAND2_X1  g690(.A1(new_n606), .A2(G953), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT119), .Z(new_n878));
  NAND2_X1  g692(.A1(new_n860), .A2(new_n863), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n323), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT56), .B1(new_n881), .B2(G210), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n236), .A2(new_n294), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(new_n292), .Z(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT55), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n878), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT118), .B1(new_n881), .B2(G210), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n879), .A2(KEYINPUT118), .A3(G210), .A4(G902), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n885), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n886), .A2(new_n891), .ZN(G51));
  INV_X1    g706(.A(new_n878), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n879), .A2(KEYINPUT54), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n868), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n324), .B(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n631), .B(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n880), .A2(new_n323), .A3(new_n760), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n893), .B1(new_n899), .B2(new_n900), .ZN(G54));
  NAND3_X1  g715(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n902));
  INV_X1    g716(.A(new_n541), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n893), .B1(new_n904), .B2(new_n905), .ZN(G60));
  NAND2_X1  g720(.A1(G478), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT59), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n640), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n893), .B1(new_n895), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n640), .B1(new_n871), .B2(new_n908), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(KEYINPUT121), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n913), .B(new_n640), .C1(new_n871), .C2(new_n908), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(G217), .A2(G902), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT122), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT60), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n879), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n424), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n893), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n658), .B(KEYINPUT123), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n879), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  OR2_X1    g739(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(KEYINPUT124), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n921), .A2(KEYINPUT124), .A3(new_n925), .A4(new_n923), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  NAND2_X1  g744(.A1(new_n822), .A2(new_n830), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT125), .Z(new_n932));
  NAND2_X1  g746(.A1(G224), .A2(G953), .ZN(new_n933));
  OAI22_X1  g747(.A1(new_n932), .A2(G953), .B1(new_n615), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(G898), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n883), .B1(new_n935), .B2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n934), .B(new_n936), .ZN(G69));
  AOI21_X1  g751(.A(new_n237), .B1(G227), .B2(G900), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n778), .A2(new_n767), .ZN(new_n942));
  INV_X1    g756(.A(new_n748), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n845), .A2(new_n731), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n506), .A2(new_n718), .ZN(new_n945));
  AOI211_X1 g759(.A(new_n943), .B(new_n944), .C1(new_n764), .C2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n746), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n942), .A2(new_n947), .A3(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n482), .B(new_n522), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(G900), .B2(G953), .ZN(new_n950));
  AOI22_X1  g764(.A1(new_n948), .A2(new_n950), .B1(new_n939), .B2(new_n938), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n695), .A2(new_n944), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n506), .A2(new_n766), .A3(new_n828), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n681), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n953), .A2(new_n767), .A3(new_n778), .A4(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n237), .ZN(new_n957));
  INV_X1    g771(.A(new_n949), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n941), .B(new_n951), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n938), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n956), .B2(new_n237), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n948), .A2(new_n950), .ZN(new_n962));
  OAI211_X1 g776(.A(KEYINPUT126), .B(new_n960), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n959), .A2(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(G472), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT63), .Z(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n956), .B2(new_n932), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n483), .A2(new_n468), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n893), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n483), .A2(new_n468), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n942), .A2(new_n947), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n966), .B1(new_n972), .B2(new_n932), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n973), .B2(KEYINPUT127), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(KEYINPUT127), .B2(new_n973), .ZN(new_n975));
  INV_X1    g789(.A(new_n968), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n857), .A2(new_n971), .A3(new_n966), .A4(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n969), .A2(new_n975), .A3(new_n977), .ZN(G57));
endmodule


