//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032;
  INV_X1    g000(.A(G134gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G127gat), .ZN(new_n203));
  INV_X1    g002(.A(G127gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G134gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n207), .B1(KEYINPUT71), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  INV_X1    g010(.A(G113gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G120gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n206), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n202), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(G127gat), .B(G134gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT70), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n209), .A2(new_n216), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT68), .B(KEYINPUT26), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT26), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n228), .A2(new_n231), .A3(KEYINPUT67), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(new_n223), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238));
  INV_X1    g037(.A(G183gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT27), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT27), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G183gat), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G190gat), .ZN(new_n244));
  AND2_X1   g043(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n240), .A2(new_n242), .A3(new_n244), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n249), .A2(new_n245), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n237), .A2(new_n238), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n248), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n225), .A2(new_n226), .B1(new_n232), .B2(new_n235), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n239), .A2(new_n244), .A3(KEYINPUT24), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n244), .A2(G183gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n256), .B1(KEYINPUT24), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n223), .B1(KEYINPUT23), .B2(new_n229), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n260), .A2(KEYINPUT25), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT23), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n266), .A2(G169gat), .A3(G176gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n265), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n266), .B1(G169gat), .B2(G176gat), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT64), .B(new_n269), .C1(new_n270), .C2(new_n223), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n268), .A2(new_n260), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n263), .A2(new_n264), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n222), .B1(new_n255), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G227gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n273), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n262), .A4(new_n260), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT71), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n206), .A3(new_n219), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n208), .A2(KEYINPUT71), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n203), .A2(new_n205), .A3(new_n220), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n202), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n288));
  OAI22_X1  g087(.A1(new_n283), .A2(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n281), .A2(new_n289), .A3(new_n254), .A4(new_n251), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n278), .A3(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G71gat), .B(G99gat), .Z(new_n292));
  XNOR2_X1  g091(.A(G15gat), .B(G43gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT73), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n291), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n275), .A2(new_n278), .A3(new_n290), .A4(new_n294), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT73), .B1(new_n299), .B2(new_n296), .ZN(new_n300));
  AND2_X1   g099(.A1(new_n291), .A2(KEYINPUT32), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT34), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n275), .A2(new_n290), .ZN(new_n304));
  INV_X1    g103(.A(new_n278), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g105(.A(KEYINPUT34), .B(new_n278), .C1(new_n275), .C2(new_n290), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n308), .B(new_n298), .C1(new_n301), .C2(new_n300), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT36), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n313), .A2(KEYINPUT36), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n310), .A2(new_n311), .A3(new_n313), .A4(KEYINPUT36), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n252), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n237), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n281), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT75), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n325), .A3(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n281), .A2(new_n254), .A3(new_n251), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n323), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n279), .A2(new_n280), .B1(new_n319), .B2(new_n237), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n339), .B(new_n322), .C1(new_n340), .C2(KEYINPUT29), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n324), .A2(new_n336), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT37), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n323), .A2(KEYINPUT29), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n337), .A2(new_n344), .B1(new_n323), .B2(new_n340), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n345), .B2(new_n335), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT38), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  NAND4_X1  g149(.A1(new_n324), .A2(new_n335), .A3(new_n338), .A4(new_n341), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n336), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n350), .A2(new_n343), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n356));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(G141gat), .A2(G148gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT78), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n362));
  INV_X1    g161(.A(G141gat), .ZN(new_n363));
  INV_X1    g162(.A(G148gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n358), .B1(new_n361), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n357), .A2(KEYINPUT77), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(G155gat), .A3(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT81), .B(G162gat), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT2), .B1(new_n379), .B2(new_n373), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT80), .A3(new_n366), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n357), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(new_n359), .B2(new_n360), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n380), .A2(new_n381), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n216), .A2(new_n206), .A3(new_n219), .A4(new_n282), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n221), .A2(new_n217), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n378), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT78), .B1(new_n359), .B2(new_n360), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n365), .A2(new_n362), .A3(new_n366), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n376), .B1(new_n391), .B2(new_n358), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n384), .A2(new_n381), .A3(new_n382), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT2), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n374), .A2(KEYINPUT81), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G162gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n394), .B1(new_n398), .B2(G155gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n289), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n388), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n389), .A2(new_n390), .B1(new_n356), .B2(new_n357), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n406), .A2(new_n376), .B1(new_n393), .B2(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT82), .A3(new_n289), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n403), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT5), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(KEYINPUT3), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n378), .A2(new_n412), .A3(new_n385), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n413), .A3(new_n289), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n407), .B2(new_n289), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n378), .A4(new_n385), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(new_n404), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n410), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT0), .ZN(new_n421));
  XNOR2_X1  g220(.A(G57gat), .B(G85gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n421), .B(new_n422), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AND3_X1   g223(.A1(new_n411), .A2(new_n413), .A3(new_n289), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n416), .A2(new_n417), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n427), .A2(KEYINPUT5), .A3(new_n404), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n351), .A2(new_n352), .ZN(new_n432));
  INV_X1    g231(.A(new_n350), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n353), .ZN(new_n436));
  INV_X1    g235(.A(new_n354), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n436), .A2(new_n437), .B1(KEYINPUT37), .B2(new_n432), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n355), .B(new_n435), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n427), .A2(new_n404), .B1(new_n409), .B2(KEYINPUT5), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT5), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n418), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n419), .A2(KEYINPUT86), .A3(new_n428), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n424), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT87), .A4(new_n424), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n419), .A2(new_n428), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT6), .B1(new_n453), .B2(new_n423), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT88), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n456));
  INV_X1    g255(.A(new_n454), .ZN(new_n457));
  AOI211_X1 g256(.A(new_n456), .B(new_n457), .C1(new_n450), .C2(new_n451), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n441), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(G22gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n335), .B1(new_n413), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n407), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT3), .B1(new_n335), .B2(new_n463), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(G228gat), .B(G233gat), .C1(new_n464), .C2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n407), .B2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n336), .ZN(new_n470));
  NAND2_X1  g269(.A1(G228gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n334), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(KEYINPUT29), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n333), .A2(new_n472), .A3(new_n334), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT3), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n470), .B(new_n471), .C1(new_n465), .C2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT31), .B(G50gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n468), .B2(new_n477), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n462), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n468), .A2(new_n477), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n478), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n477), .A3(new_n479), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n461), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n403), .A2(new_n408), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n404), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n405), .B1(new_n425), .B2(new_n426), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT39), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n423), .B1(new_n490), .B2(KEYINPUT39), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  OAI22_X1  g292(.A1(new_n491), .A2(new_n492), .B1(KEYINPUT85), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT85), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(KEYINPUT40), .ZN(new_n496));
  OAI211_X1 g295(.A(KEYINPUT85), .B(new_n493), .C1(new_n491), .C2(new_n492), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n450), .B2(new_n451), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n434), .A2(KEYINPUT30), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT30), .A4(new_n350), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(new_n353), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n487), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n318), .B1(new_n459), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n434), .A2(KEYINPUT30), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n424), .B1(new_n419), .B2(new_n428), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n423), .B1(new_n443), .B2(new_n445), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(KEYINPUT83), .A3(new_n430), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n512), .A3(new_n429), .ZN(new_n513));
  INV_X1    g312(.A(new_n431), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT76), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n502), .B2(new_n353), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n436), .A2(KEYINPUT76), .A3(new_n501), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n487), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n514), .B1(new_n455), .B2(new_n458), .ZN(new_n523));
  INV_X1    g322(.A(new_n487), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n312), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n525), .A2(new_n504), .A3(KEYINPUT35), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n487), .B1(new_n310), .B2(new_n311), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI211_X1 g329(.A(KEYINPUT89), .B(new_n487), .C1(new_n310), .C2(new_n311), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT35), .B1(new_n532), .B2(new_n521), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n506), .A2(new_n522), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G1gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n537), .A3(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT16), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(G8gat), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT91), .B(G29gat), .Z(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT92), .B(G36gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT14), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  XNOR2_X1  g351(.A(G43gat), .B(G50gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT15), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n552), .B1(new_n551), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n553), .A2(KEYINPUT15), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n551), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(KEYINPUT94), .A2(KEYINPUT17), .ZN(new_n561));
  NOR2_X1   g360(.A1(KEYINPUT94), .A2(KEYINPUT17), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n559), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n555), .B2(new_n556), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT94), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n545), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G8gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n544), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT96), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n545), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n576), .A2(new_n566), .ZN(new_n577));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n570), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT97), .B(KEYINPUT18), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n535), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G113gat), .B(G141gat), .Z(new_n584));
  XNOR2_X1  g383(.A(G169gat), .B(G197gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT12), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n564), .A2(new_n569), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n572), .ZN(new_n592));
  INV_X1    g391(.A(new_n577), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n592), .A2(KEYINPUT18), .A3(new_n578), .A4(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n578), .B(KEYINPUT13), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n576), .A2(new_n566), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n596), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n592), .A2(new_n578), .A3(new_n593), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n581), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n590), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n598), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n602), .B(new_n594), .C1(new_n580), .C2(new_n582), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(new_n583), .A3(new_n589), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT99), .B1(new_n534), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n601), .A2(new_n604), .ZN(new_n608));
  AOI221_X4 g407(.A(new_n318), .B1(new_n521), .B2(new_n487), .C1(new_n459), .C2(new_n505), .ZN(new_n609));
  INV_X1    g408(.A(new_n429), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n610), .B1(new_n454), .B2(KEYINPUT83), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n431), .B1(new_n611), .B2(new_n510), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n612), .A2(new_n507), .A3(new_n519), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n530), .B2(new_n531), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n614), .A2(KEYINPUT35), .B1(new_n523), .B2(new_n526), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n607), .B(new_n608), .C1(new_n609), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n606), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT7), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  INV_X1    g419(.A(G85gat), .ZN(new_n621));
  INV_X1    g420(.A(G92gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(KEYINPUT8), .A2(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G99gat), .B(G106gat), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n619), .A3(new_n623), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G57gat), .B(G64gat), .Z(new_n630));
  INV_X1    g429(.A(KEYINPUT9), .ZN(new_n631));
  INV_X1    g430(.A(G71gat), .ZN(new_n632));
  INV_X1    g431(.A(G78gat), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G71gat), .B(G78gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n630), .A2(new_n636), .A3(new_n634), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(KEYINPUT100), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT100), .B1(new_n638), .B2(new_n639), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n629), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n629), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  AND3_X1   g450(.A1(new_n645), .A2(new_n628), .A3(new_n626), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n640), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n652), .B1(new_n655), .B2(new_n629), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n651), .B1(new_n656), .B2(KEYINPUT10), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n647), .A2(KEYINPUT103), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n629), .A2(new_n658), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n657), .A2(new_n659), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n648), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n650), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n655), .A2(new_n660), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT103), .B1(new_n647), .B2(new_n658), .ZN(new_n665));
  AOI211_X1 g464(.A(new_n651), .B(KEYINPUT10), .C1(new_n643), .C2(new_n646), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(KEYINPUT104), .A3(new_n648), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n649), .B1(new_n663), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G120gat), .B(G148gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(G176gat), .B(G204gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(KEYINPUT105), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n669), .B2(new_n673), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n667), .A2(new_n648), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n649), .A2(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(G190gat), .B(G218gat), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n591), .A2(new_n629), .ZN(new_n685));
  AND2_X1   g484(.A1(G232gat), .A2(G233gat), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n560), .A2(new_n644), .B1(KEYINPUT41), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n684), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n685), .A2(new_n684), .A3(new_n687), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n686), .A2(KEYINPUT41), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G134gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n374), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n694), .B1(new_n688), .B2(KEYINPUT102), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n655), .A2(KEYINPUT21), .ZN(new_n700));
  XOR2_X1   g499(.A(G127gat), .B(G155gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n573), .A2(new_n575), .B1(KEYINPUT21), .B2(new_n655), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(G231gat), .A2(G233gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT101), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(G183gat), .B(G211gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n704), .B(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n682), .A2(new_n699), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n617), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n617), .A2(KEYINPUT106), .A3(new_n713), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n612), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g519(.A(new_n571), .B1(new_n718), .B2(new_n504), .ZN(new_n721));
  INV_X1    g520(.A(new_n504), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT16), .B(G8gat), .ZN(new_n723));
  AOI211_X1 g522(.A(new_n722), .B(new_n723), .C1(new_n716), .C2(new_n717), .ZN(new_n724));
  OAI21_X1  g523(.A(KEYINPUT42), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n718), .A2(new_n504), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n723), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(G1325gat));
  INV_X1    g528(.A(new_n718), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n318), .B(KEYINPUT107), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G15gat), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(G15gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n734), .A3(new_n312), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1326gat));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n617), .B2(new_n713), .ZN(new_n737));
  INV_X1    g536(.A(new_n713), .ZN(new_n738));
  AOI211_X1 g537(.A(new_n715), .B(new_n738), .C1(new_n606), .C2(new_n616), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n487), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT108), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT108), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n742), .B(new_n487), .C1(new_n737), .C2(new_n739), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT43), .B(G22gat), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n741), .B2(new_n743), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1327gat));
  NOR2_X1   g546(.A1(new_n682), .A2(new_n711), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n698), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n617), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n751), .A2(new_n612), .A3(new_n546), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n749), .A2(new_n605), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT109), .B1(new_n613), .B2(new_n524), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n521), .A2(new_n760), .A3(new_n487), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n318), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n423), .B1(new_n453), .B2(new_n442), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT87), .B1(new_n764), .B2(new_n447), .ZN(new_n765));
  AND4_X1   g564(.A1(KEYINPUT87), .A2(new_n446), .A3(new_n424), .A4(new_n447), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n454), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n456), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n452), .A2(KEYINPUT88), .A3(new_n454), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n440), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n452), .A2(new_n496), .A3(new_n497), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n524), .B1(new_n771), .B2(new_n722), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n763), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(KEYINPUT110), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n760), .B1(new_n521), .B2(new_n487), .ZN(new_n775));
  AOI211_X1 g574(.A(KEYINPUT109), .B(new_n524), .C1(new_n515), .C2(new_n520), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n506), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n527), .A2(new_n533), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n758), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n783));
  INV_X1    g582(.A(new_n534), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n699), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n756), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n612), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n754), .B(new_n755), .C1(new_n546), .C2(new_n788), .ZN(G1328gat));
  AND3_X1   g588(.A1(new_n751), .A2(new_n504), .A3(new_n547), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n786), .A2(new_n722), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n793), .C1(new_n547), .C2(new_n794), .ZN(G1329gat));
  OAI21_X1  g594(.A(G43gat), .B1(new_n786), .B2(new_n763), .ZN(new_n796));
  INV_X1    g595(.A(G43gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n751), .A2(new_n797), .A3(new_n312), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(KEYINPUT47), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n731), .B(new_n756), .C1(new_n782), .C2(new_n785), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G43gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n798), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT111), .B(KEYINPUT47), .C1(new_n802), .C2(new_n798), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n799), .B1(new_n805), .B2(new_n806), .ZN(G1330gat));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n487), .B(new_n756), .C1(new_n782), .C2(new_n785), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(G50gat), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n524), .A2(G50gat), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n617), .A2(new_n750), .A3(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n808), .B(new_n809), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n809), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n813), .B1(G50gat), .B2(new_n810), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(KEYINPUT112), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n814), .A2(new_n817), .ZN(G1331gat));
  AOI21_X1  g617(.A(new_n615), .B1(new_n774), .B2(new_n779), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n675), .A2(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n605), .A2(new_n698), .A3(new_n711), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n612), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g623(.A(new_n504), .B(KEYINPUT114), .Z(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT115), .ZN(new_n828));
  NOR2_X1   g627(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n828), .B(new_n829), .ZN(G1333gat));
  NAND3_X1  g629(.A1(new_n822), .A2(new_n632), .A3(new_n312), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n822), .A2(new_n731), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n632), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g633(.A1(new_n822), .A2(new_n487), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g635(.A1(new_n780), .A2(new_n781), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n608), .A2(new_n711), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n699), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(KEYINPUT51), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT51), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n842), .B1(new_n819), .B2(new_n839), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n820), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n621), .A3(new_n612), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n820), .A2(new_n608), .A3(new_n711), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n782), .B2(new_n785), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT116), .B1(new_n847), .B2(new_n787), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G85gat), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n847), .A2(KEYINPUT116), .A3(new_n787), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(G1336gat));
  INV_X1    g650(.A(new_n825), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n852), .B(new_n846), .C1(new_n782), .C2(new_n785), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G92gat), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n622), .A3(new_n682), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT117), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n837), .B2(new_n840), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n819), .A2(new_n842), .A3(new_n839), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n854), .A2(new_n855), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n504), .B(new_n846), .C1(new_n782), .C2(new_n785), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G92gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n855), .B1(new_n863), .B2(new_n860), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT118), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n854), .A2(new_n855), .A3(new_n860), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n841), .A2(new_n843), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n868), .A2(new_n857), .B1(new_n862), .B2(G92gat), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n866), .B(new_n867), .C1(new_n869), .C2(new_n855), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n865), .A2(new_n870), .ZN(G1337gat));
  INV_X1    g670(.A(G99gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n844), .A2(new_n872), .A3(new_n312), .ZN(new_n873));
  OAI21_X1  g672(.A(G99gat), .B1(new_n847), .B2(new_n732), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1338gat));
  AOI21_X1  g674(.A(G106gat), .B1(new_n844), .B2(new_n487), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n877));
  INV_X1    g676(.A(G106gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n847), .A2(new_n878), .A3(new_n524), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n876), .B2(new_n879), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1339gat));
  NAND2_X1  g681(.A1(new_n713), .A2(new_n605), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n603), .A2(new_n589), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n578), .B1(new_n592), .B2(new_n593), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n593), .A2(new_n597), .A3(new_n596), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n588), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n889), .B1(new_n667), .B2(new_n648), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n662), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n673), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n663), .A2(new_n668), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT55), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT55), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n681), .A3(new_n897), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n888), .A2(new_n698), .A3(new_n898), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n605), .A2(new_n898), .B1(new_n820), .B2(new_n888), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n698), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n883), .B1(new_n901), .B2(new_n711), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n902), .A2(new_n528), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n852), .A2(new_n787), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(new_n212), .A3(new_n605), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n902), .A2(new_n612), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(new_n532), .A3(new_n852), .ZN(new_n908));
  AOI21_X1  g707(.A(G113gat), .B1(new_n908), .B2(new_n608), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n906), .A2(new_n909), .ZN(G1340gat));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n210), .A3(new_n682), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n903), .A2(new_n682), .A3(new_n904), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(KEYINPUT119), .A3(G120gat), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT119), .B1(new_n912), .B2(G120gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1341gat));
  OAI21_X1  g714(.A(G127gat), .B1(new_n905), .B2(new_n712), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n908), .A2(new_n204), .A3(new_n711), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1342gat));
  INV_X1    g717(.A(new_n907), .ZN(new_n919));
  INV_X1    g718(.A(new_n532), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n698), .A2(new_n504), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n919), .A2(new_n202), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n923));
  OAI21_X1  g722(.A(G134gat), .B1(new_n905), .B2(new_n698), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G1343gat));
  NOR3_X1   g725(.A1(new_n852), .A2(new_n787), .A3(new_n318), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n898), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n896), .A2(KEYINPUT120), .A3(new_n681), .A4(new_n897), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n930), .A2(new_n608), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n682), .A2(new_n887), .A3(new_n884), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n699), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n712), .B1(new_n934), .B2(new_n899), .ZN(new_n935));
  AOI211_X1 g734(.A(new_n928), .B(new_n524), .C1(new_n935), .C2(new_n883), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT57), .B1(new_n902), .B2(new_n487), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n608), .B(new_n927), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(G141gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n732), .A2(new_n487), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n605), .A2(G141gat), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(new_n825), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n919), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n919), .A2(KEYINPUT122), .A3(new_n942), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT58), .B1(new_n939), .B2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT58), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n919), .A2(new_n942), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT123), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT123), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n919), .A2(new_n954), .A3(new_n942), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n953), .A2(new_n825), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(new_n943), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n950), .B1(new_n939), .B2(new_n958), .ZN(G1344gat));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n927), .B1(new_n936), .B2(new_n937), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n960), .B(G148gat), .C1(new_n961), .C2(new_n820), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n902), .A2(KEYINPUT57), .A3(new_n487), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n524), .B1(new_n935), .B2(new_n883), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(KEYINPUT57), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n927), .A2(new_n682), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n364), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n962), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n682), .A2(new_n364), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n956), .B2(new_n969), .ZN(G1345gat));
  OAI21_X1  g769(.A(G155gat), .B1(new_n961), .B2(new_n712), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n711), .A2(new_n373), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n956), .B2(new_n972), .ZN(G1346gat));
  NAND4_X1  g772(.A1(new_n953), .A2(new_n379), .A3(new_n921), .A4(new_n955), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n398), .B1(new_n961), .B2(new_n698), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT124), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n974), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1347gat));
  NOR2_X1   g779(.A1(new_n722), .A2(new_n612), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n903), .A2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(G169gat), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n982), .A2(new_n983), .A3(new_n605), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n902), .A2(new_n787), .ZN(new_n985));
  AND3_X1   g784(.A1(new_n985), .A2(new_n920), .A3(new_n852), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(new_n608), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n984), .B1(new_n987), .B2(new_n983), .ZN(G1348gat));
  INV_X1    g787(.A(G176gat), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n986), .A2(new_n989), .A3(new_n682), .ZN(new_n990));
  OAI21_X1  g789(.A(G176gat), .B1(new_n982), .B2(new_n820), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT125), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n992), .B(new_n993), .ZN(G1349gat));
  NAND3_X1  g793(.A1(new_n986), .A2(new_n243), .A3(new_n711), .ZN(new_n995));
  OAI21_X1  g794(.A(G183gat), .B1(new_n982), .B2(new_n712), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g796(.A(new_n997), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g797(.A1(new_n986), .A2(new_n244), .A3(new_n699), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n903), .A2(new_n699), .A3(new_n981), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT61), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n1000), .A2(new_n1001), .A3(G190gat), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n1001), .B1(new_n1000), .B2(G190gat), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n999), .B1(new_n1002), .B2(new_n1003), .ZN(G1351gat));
  NAND2_X1  g803(.A1(new_n902), .A2(new_n787), .ZN(new_n1005));
  NOR3_X1   g804(.A1(new_n1005), .A2(new_n825), .A3(new_n940), .ZN(new_n1006));
  INV_X1    g805(.A(G197gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1006), .A2(new_n1007), .A3(new_n608), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n732), .A2(new_n608), .A3(new_n981), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n965), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g810(.A(KEYINPUT126), .B(new_n963), .C1(new_n964), .C2(KEYINPUT57), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014));
  OAI21_X1  g813(.A(G197gat), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g814(.A(KEYINPUT127), .B(new_n1009), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1008), .B1(new_n1015), .B2(new_n1016), .ZN(G1352gat));
  INV_X1    g816(.A(G204gat), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1006), .A2(new_n1018), .A3(new_n682), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT62), .ZN(new_n1020));
  XNOR2_X1  g819(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n732), .A2(new_n981), .ZN(new_n1022));
  AOI21_X1  g821(.A(new_n1022), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1023));
  AND2_X1   g822(.A1(new_n1023), .A2(new_n682), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1024), .B2(new_n1018), .ZN(G1353gat));
  NOR2_X1   g824(.A1(new_n1022), .A2(new_n712), .ZN(new_n1026));
  AOI21_X1  g825(.A(new_n327), .B1(new_n965), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g826(.A(new_n1027), .B(KEYINPUT63), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1006), .A2(new_n327), .A3(new_n711), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1028), .A2(new_n1029), .ZN(G1354gat));
  AOI21_X1  g829(.A(G218gat), .B1(new_n1006), .B2(new_n699), .ZN(new_n1031));
  NOR2_X1   g830(.A1(new_n698), .A2(new_n328), .ZN(new_n1032));
  AOI21_X1  g831(.A(new_n1031), .B1(new_n1023), .B2(new_n1032), .ZN(G1355gat));
endmodule


