

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743;

  XNOR2_X1 U366 ( .A(G101), .B(KEYINPUT85), .ZN(n388) );
  BUF_X1 U367 ( .A(n717), .Z(n342) );
  NOR2_X2 U368 ( .A1(n596), .A2(n595), .ZN(n597) );
  AND2_X2 U369 ( .A1(n362), .A2(n366), .ZN(n351) );
  NOR2_X2 U370 ( .A1(n367), .A2(n404), .ZN(n358) );
  NAND2_X2 U371 ( .A1(n708), .A2(n402), .ZN(n367) );
  OR2_X2 U372 ( .A1(n708), .A2(n363), .ZN(n362) );
  XNOR2_X2 U373 ( .A(n591), .B(n398), .ZN(n708) );
  XNOR2_X2 U374 ( .A(n445), .B(n431), .ZN(n580) );
  INV_X1 U375 ( .A(G953), .ZN(n679) );
  INV_X2 U376 ( .A(G146), .ZN(n439) );
  NOR2_X1 U377 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U378 ( .A1(n647), .A2(n657), .ZN(n368) );
  BUF_X1 U379 ( .A(n482), .Z(n605) );
  NAND2_X1 U380 ( .A1(n536), .A2(n537), .ZN(n369) );
  XNOR2_X1 U381 ( .A(n412), .B(n411), .ZN(n581) );
  XNOR2_X1 U382 ( .A(G110), .B(G107), .ZN(n350) );
  NOR2_X1 U383 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U384 ( .A1(n381), .A2(n598), .ZN(n380) );
  XNOR2_X1 U385 ( .A(n369), .B(KEYINPUT100), .ZN(n647) );
  XNOR2_X1 U386 ( .A(n528), .B(n527), .ZN(n531) );
  XNOR2_X1 U387 ( .A(n479), .B(n478), .ZN(n536) );
  OR2_X1 U388 ( .A1(n726), .A2(G902), .ZN(n438) );
  XNOR2_X1 U389 ( .A(n421), .B(n420), .ZN(n719) );
  XNOR2_X1 U390 ( .A(n581), .B(n385), .ZN(n421) );
  XNOR2_X1 U391 ( .A(n350), .B(G104), .ZN(n435) );
  XNOR2_X1 U392 ( .A(n399), .B(G902), .ZN(n686) );
  XNOR2_X1 U393 ( .A(G116), .B(G113), .ZN(n389) );
  XNOR2_X1 U394 ( .A(KEYINPUT84), .B(KEYINPUT15), .ZN(n399) );
  XNOR2_X2 U395 ( .A(n380), .B(KEYINPUT33), .ZN(n652) );
  BUF_X1 U396 ( .A(n638), .Z(n343) );
  BUF_X1 U397 ( .A(n726), .Z(n344) );
  BUF_X1 U398 ( .A(n722), .Z(n345) );
  INV_X1 U399 ( .A(n378), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n597), .B(KEYINPUT35), .ZN(n717) );
  NAND2_X1 U401 ( .A1(n362), .A2(n361), .ZN(n360) );
  AND2_X1 U402 ( .A1(n366), .A2(n643), .ZN(n361) );
  NOR2_X1 U403 ( .A1(n354), .A2(KEYINPUT78), .ZN(n353) );
  INV_X1 U404 ( .A(n367), .ZN(n354) );
  XNOR2_X1 U405 ( .A(n422), .B(KEYINPUT20), .ZN(n425) );
  NAND2_X1 U406 ( .A1(n425), .A2(G217), .ZN(n384) );
  XNOR2_X1 U407 ( .A(n454), .B(n460), .ZN(n372) );
  XNOR2_X1 U408 ( .A(G140), .B(G137), .ZN(n431) );
  NAND2_X1 U409 ( .A1(n400), .A2(n402), .ZN(n366) );
  NAND2_X1 U410 ( .A1(n365), .A2(n364), .ZN(n363) );
  XNOR2_X1 U411 ( .A(n463), .B(G475), .ZN(n464) );
  XNOR2_X1 U412 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n411) );
  NAND2_X1 U413 ( .A1(n526), .A2(n643), .ZN(n528) );
  INV_X1 U414 ( .A(KEYINPUT30), .ZN(n527) );
  NAND2_X1 U415 ( .A1(n355), .A2(n353), .ZN(n352) );
  INV_X1 U416 ( .A(n360), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n384), .B(n383), .ZN(n382) );
  XNOR2_X1 U418 ( .A(n423), .B(KEYINPUT87), .ZN(n383) );
  XNOR2_X1 U419 ( .A(G119), .B(G128), .ZN(n413) );
  XOR2_X1 U420 ( .A(KEYINPUT76), .B(KEYINPUT8), .Z(n415) );
  XNOR2_X1 U421 ( .A(n371), .B(n370), .ZN(n702) );
  XNOR2_X1 U422 ( .A(n462), .B(n461), .ZN(n370) );
  XNOR2_X1 U423 ( .A(n372), .B(n581), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n580), .B(n437), .ZN(n726) );
  XOR2_X1 U425 ( .A(n368), .B(KEYINPUT101), .Z(n347) );
  XNOR2_X1 U426 ( .A(n428), .B(KEYINPUT66), .ZN(n660) );
  AND2_X1 U427 ( .A1(n379), .A2(n378), .ZN(n348) );
  INV_X1 U428 ( .A(KEYINPUT78), .ZN(n404) );
  XNOR2_X1 U429 ( .A(KEYINPUT81), .B(KEYINPUT0), .ZN(n349) );
  XNOR2_X2 U430 ( .A(n522), .B(KEYINPUT22), .ZN(n602) );
  XNOR2_X2 U431 ( .A(n429), .B(G134), .ZN(n472) );
  XNOR2_X2 U432 ( .A(n472), .B(n430), .ZN(n445) );
  NAND2_X1 U433 ( .A1(n351), .A2(n367), .ZN(n556) );
  NAND2_X2 U434 ( .A1(n356), .A2(n352), .ZN(n495) );
  AND2_X2 U435 ( .A1(n359), .A2(n357), .ZN(n356) );
  INV_X1 U436 ( .A(n358), .ZN(n357) );
  NAND2_X1 U437 ( .A1(n360), .A2(KEYINPUT78), .ZN(n359) );
  INV_X1 U438 ( .A(n402), .ZN(n364) );
  INV_X1 U439 ( .A(n400), .ZN(n365) );
  NOR2_X1 U440 ( .A1(n702), .A2(G902), .ZN(n465) );
  NAND2_X1 U441 ( .A1(n375), .A2(n373), .ZN(n381) );
  NAND2_X1 U442 ( .A1(n374), .A2(n379), .ZN(n373) );
  INV_X1 U443 ( .A(n660), .ZN(n379) );
  NOR2_X1 U444 ( .A1(n510), .A2(n592), .ZN(n374) );
  AND2_X1 U445 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U446 ( .A1(n510), .A2(n592), .ZN(n376) );
  NAND2_X1 U447 ( .A1(n660), .A2(n592), .ZN(n377) );
  INV_X1 U448 ( .A(n510), .ZN(n378) );
  XNOR2_X2 U449 ( .A(n424), .B(n382), .ZN(n482) );
  INV_X1 U450 ( .A(n593), .ZN(n511) );
  AND2_X2 U451 ( .A1(n593), .A2(n347), .ZN(n522) );
  XNOR2_X2 U452 ( .A(n410), .B(n349), .ZN(n593) );
  XNOR2_X2 U453 ( .A(n495), .B(KEYINPUT19), .ZN(n548) );
  XNOR2_X1 U454 ( .A(n413), .B(n431), .ZN(n385) );
  AND2_X1 U455 ( .A1(n554), .A2(n553), .ZN(n386) );
  INV_X1 U456 ( .A(n569), .ZN(n570) );
  NOR2_X1 U457 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U458 ( .A1(n386), .A2(n572), .ZN(n574) );
  BUF_X1 U459 ( .A(n652), .Z(n677) );
  XNOR2_X1 U460 ( .A(n465), .B(n464), .ZN(n537) );
  INV_X1 U461 ( .A(KEYINPUT105), .ZN(n534) );
  INV_X1 U462 ( .A(KEYINPUT39), .ZN(n558) );
  XNOR2_X1 U463 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n562) );
  XNOR2_X1 U464 ( .A(n563), .B(n562), .ZN(n742) );
  XNOR2_X1 U465 ( .A(KEYINPUT16), .B(G122), .ZN(n387) );
  XNOR2_X1 U466 ( .A(n435), .B(n387), .ZN(n392) );
  XNOR2_X1 U467 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U468 ( .A(KEYINPUT3), .B(G119), .ZN(n390) );
  XNOR2_X1 U469 ( .A(n391), .B(n390), .ZN(n444) );
  XNOR2_X1 U470 ( .A(n392), .B(n444), .ZN(n591) );
  XNOR2_X1 U471 ( .A(n439), .B(G125), .ZN(n412) );
  NAND2_X1 U472 ( .A1(n679), .A2(G224), .ZN(n393) );
  XNOR2_X1 U473 ( .A(n393), .B(KEYINPUT4), .ZN(n394) );
  XNOR2_X1 U474 ( .A(n412), .B(n394), .ZN(n397) );
  XNOR2_X2 U475 ( .A(G143), .B(G128), .ZN(n429) );
  XNOR2_X1 U476 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n395) );
  XNOR2_X1 U477 ( .A(n429), .B(n395), .ZN(n396) );
  XNOR2_X1 U478 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X1 U479 ( .A(n686), .ZN(n400) );
  INV_X1 U480 ( .A(G902), .ZN(n476) );
  INV_X1 U481 ( .A(G237), .ZN(n401) );
  NAND2_X1 U482 ( .A1(n476), .A2(n401), .ZN(n403) );
  NAND2_X1 U483 ( .A1(n403), .A2(G210), .ZN(n402) );
  NAND2_X1 U484 ( .A1(n403), .A2(G214), .ZN(n643) );
  NAND2_X1 U485 ( .A1(G237), .A2(G234), .ZN(n405) );
  XOR2_X1 U486 ( .A(KEYINPUT14), .B(n405), .Z(n486) );
  INV_X1 U487 ( .A(G952), .ZN(n694) );
  NOR2_X1 U488 ( .A1(n694), .A2(G953), .ZN(n407) );
  NAND2_X1 U489 ( .A1(G953), .A2(G902), .ZN(n483) );
  NOR2_X1 U490 ( .A1(G898), .A2(n483), .ZN(n406) );
  NOR2_X1 U491 ( .A1(n407), .A2(n406), .ZN(n408) );
  NOR2_X1 U492 ( .A1(n486), .A2(n408), .ZN(n409) );
  NAND2_X1 U493 ( .A1(n548), .A2(n409), .ZN(n410) );
  NAND2_X1 U494 ( .A1(n679), .A2(G234), .ZN(n414) );
  XNOR2_X1 U495 ( .A(n415), .B(n414), .ZN(n471) );
  NAND2_X1 U496 ( .A1(n471), .A2(G221), .ZN(n419) );
  XOR2_X1 U497 ( .A(KEYINPUT70), .B(KEYINPUT24), .Z(n417) );
  XNOR2_X1 U498 ( .A(G110), .B(KEYINPUT23), .ZN(n416) );
  XNOR2_X1 U499 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U500 ( .A(n419), .B(n418), .ZN(n420) );
  NAND2_X1 U501 ( .A1(n719), .A2(n476), .ZN(n424) );
  NAND2_X1 U502 ( .A1(n686), .A2(G234), .ZN(n422) );
  XOR2_X1 U503 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n423) );
  NAND2_X1 U504 ( .A1(n425), .A2(G221), .ZN(n426) );
  XNOR2_X1 U505 ( .A(n426), .B(KEYINPUT21), .ZN(n657) );
  INV_X1 U506 ( .A(n657), .ZN(n427) );
  NAND2_X1 U507 ( .A1(n482), .A2(n427), .ZN(n428) );
  XNOR2_X1 U508 ( .A(KEYINPUT4), .B(G131), .ZN(n430) );
  NAND2_X1 U509 ( .A1(n679), .A2(G227), .ZN(n432) );
  XNOR2_X1 U510 ( .A(n432), .B(KEYINPUT86), .ZN(n434) );
  XNOR2_X1 U511 ( .A(n439), .B(G101), .ZN(n433) );
  XNOR2_X1 U512 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U513 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X2 U514 ( .A(n438), .B(G469), .ZN(n500) );
  INV_X1 U515 ( .A(n500), .ZN(n545) );
  NOR2_X2 U516 ( .A1(G953), .A2(G237), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n459), .A2(G210), .ZN(n440) );
  XNOR2_X1 U518 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U519 ( .A(KEYINPUT5), .B(G137), .Z(n441) );
  XNOR2_X1 U520 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U521 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U522 ( .A(n446), .B(n445), .ZN(n691) );
  NAND2_X1 U523 ( .A1(n691), .A2(n476), .ZN(n449) );
  INV_X1 U524 ( .A(KEYINPUT71), .ZN(n447) );
  XNOR2_X1 U525 ( .A(n447), .B(G472), .ZN(n448) );
  XNOR2_X1 U526 ( .A(n449), .B(n448), .ZN(n526) );
  BUF_X1 U527 ( .A(n526), .Z(n664) );
  NOR2_X1 U528 ( .A1(n545), .A2(n664), .ZN(n450) );
  NAND2_X1 U529 ( .A1(n379), .A2(n450), .ZN(n451) );
  NOR2_X1 U530 ( .A1(n511), .A2(n451), .ZN(n619) );
  XOR2_X1 U531 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n453) );
  XNOR2_X1 U532 ( .A(G143), .B(G122), .ZN(n452) );
  XNOR2_X1 U533 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U534 ( .A(G140), .B(G104), .Z(n456) );
  XNOR2_X1 U535 ( .A(G113), .B(G131), .ZN(n455) );
  XNOR2_X1 U536 ( .A(n456), .B(n455), .ZN(n462) );
  XOR2_X1 U537 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n458) );
  XNOR2_X1 U538 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n457) );
  XNOR2_X1 U539 ( .A(n458), .B(n457), .ZN(n461) );
  NAND2_X1 U540 ( .A1(G214), .A2(n459), .ZN(n460) );
  XNOR2_X1 U541 ( .A(KEYINPUT93), .B(KEYINPUT13), .ZN(n463) );
  XOR2_X1 U542 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n467) );
  XNOR2_X1 U543 ( .A(G107), .B(G122), .ZN(n466) );
  XNOR2_X1 U544 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U545 ( .A(n468), .B(KEYINPUT94), .Z(n470) );
  XNOR2_X1 U546 ( .A(G116), .B(KEYINPUT95), .ZN(n469) );
  XNOR2_X1 U547 ( .A(n470), .B(n469), .ZN(n475) );
  NAND2_X1 U548 ( .A1(n471), .A2(G217), .ZN(n473) );
  XNOR2_X1 U549 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U550 ( .A(n475), .B(n474), .ZN(n724) );
  NAND2_X1 U551 ( .A1(n724), .A2(n476), .ZN(n479) );
  XOR2_X1 U552 ( .A(G478), .B(KEYINPUT97), .Z(n477) );
  XOR2_X1 U553 ( .A(KEYINPUT96), .B(n477), .Z(n478) );
  INV_X1 U554 ( .A(n536), .ZN(n505) );
  OR2_X1 U555 ( .A1(n537), .A2(n505), .ZN(n480) );
  XNOR2_X1 U556 ( .A(n480), .B(KEYINPUT98), .ZN(n560) );
  INV_X1 U557 ( .A(n560), .ZN(n736) );
  NAND2_X1 U558 ( .A1(n619), .A2(n736), .ZN(n481) );
  XNOR2_X1 U559 ( .A(n481), .B(G104), .ZN(G6) );
  NOR2_X1 U560 ( .A1(n486), .A2(n483), .ZN(n484) );
  XNOR2_X1 U561 ( .A(n484), .B(KEYINPUT103), .ZN(n485) );
  NOR2_X1 U562 ( .A1(G900), .A2(n485), .ZN(n489) );
  INV_X1 U563 ( .A(n486), .ZN(n487) );
  NAND2_X1 U564 ( .A1(n487), .A2(G952), .ZN(n674) );
  NOR2_X1 U565 ( .A1(n674), .A2(G953), .ZN(n488) );
  NOR2_X1 U566 ( .A1(n489), .A2(n488), .ZN(n529) );
  NOR2_X1 U567 ( .A1(n657), .A2(n529), .ZN(n490) );
  XNOR2_X1 U568 ( .A(n490), .B(KEYINPUT69), .ZN(n491) );
  NOR2_X1 U569 ( .A1(n605), .A2(n491), .ZN(n543) );
  INV_X1 U570 ( .A(KEYINPUT6), .ZN(n492) );
  XNOR2_X1 U571 ( .A(n664), .B(n492), .ZN(n598) );
  NAND2_X1 U572 ( .A1(n543), .A2(n598), .ZN(n493) );
  NOR2_X1 U573 ( .A1(n493), .A2(n560), .ZN(n494) );
  XNOR2_X1 U574 ( .A(KEYINPUT104), .B(n494), .ZN(n515) );
  INV_X1 U575 ( .A(n495), .ZN(n496) );
  NAND2_X1 U576 ( .A1(n515), .A2(n496), .ZN(n498) );
  XOR2_X1 U577 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n497) );
  XNOR2_X1 U578 ( .A(n498), .B(n497), .ZN(n501) );
  XNOR2_X1 U579 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n499) );
  XNOR2_X2 U580 ( .A(n500), .B(n499), .ZN(n510) );
  NAND2_X1 U581 ( .A1(n501), .A2(n378), .ZN(n569) );
  XOR2_X1 U582 ( .A(G125), .B(KEYINPUT37), .Z(n502) );
  XNOR2_X1 U583 ( .A(n569), .B(n502), .ZN(G27) );
  XOR2_X1 U584 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n504) );
  XNOR2_X1 U585 ( .A(G107), .B(KEYINPUT113), .ZN(n503) );
  XNOR2_X1 U586 ( .A(n504), .B(n503), .ZN(n509) );
  NAND2_X1 U587 ( .A1(n537), .A2(n505), .ZN(n507) );
  INV_X1 U588 ( .A(KEYINPUT99), .ZN(n506) );
  XNOR2_X1 U589 ( .A(n507), .B(n506), .ZN(n575) );
  INV_X1 U590 ( .A(n575), .ZN(n733) );
  NAND2_X1 U591 ( .A1(n619), .A2(n733), .ZN(n508) );
  XOR2_X1 U592 ( .A(n509), .B(n508), .Z(G9) );
  NAND2_X1 U593 ( .A1(n348), .A2(n664), .ZN(n667) );
  NOR2_X1 U594 ( .A1(n511), .A2(n667), .ZN(n513) );
  XOR2_X1 U595 ( .A(KEYINPUT88), .B(KEYINPUT31), .Z(n512) );
  XNOR2_X1 U596 ( .A(n513), .B(n512), .ZN(n620) );
  NAND2_X1 U597 ( .A1(n620), .A2(n736), .ZN(n514) );
  XNOR2_X1 U598 ( .A(n514), .B(G113), .ZN(G15) );
  NAND2_X1 U599 ( .A1(n515), .A2(n643), .ZN(n516) );
  NOR2_X1 U600 ( .A1(n516), .A2(n378), .ZN(n517) );
  XNOR2_X1 U601 ( .A(n517), .B(KEYINPUT43), .ZN(n519) );
  INV_X1 U602 ( .A(n556), .ZN(n518) );
  NOR2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n577) );
  XOR2_X1 U604 ( .A(G140), .B(n577), .Z(G42) );
  XNOR2_X1 U605 ( .A(G116), .B(KEYINPUT115), .ZN(n521) );
  NAND2_X1 U606 ( .A1(n620), .A2(n733), .ZN(n520) );
  XOR2_X1 U607 ( .A(n521), .B(n520), .Z(G18) );
  XNOR2_X1 U608 ( .A(G101), .B(KEYINPUT112), .ZN(n525) );
  INV_X1 U609 ( .A(n602), .ZN(n608) );
  INV_X1 U610 ( .A(n605), .ZN(n656) );
  NOR2_X1 U611 ( .A1(n598), .A2(n656), .ZN(n523) );
  NAND2_X1 U612 ( .A1(n346), .A2(n523), .ZN(n524) );
  NOR2_X1 U613 ( .A1(n608), .A2(n524), .ZN(n623) );
  XOR2_X1 U614 ( .A(n525), .B(n623), .Z(G3) );
  AND2_X1 U615 ( .A1(n560), .A2(n575), .ZN(n649) );
  NAND2_X1 U616 ( .A1(n649), .A2(KEYINPUT47), .ZN(n541) );
  INV_X1 U617 ( .A(n529), .ZN(n530) );
  NAND2_X1 U618 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U619 ( .A1(n532), .A2(n545), .ZN(n555) );
  NAND2_X1 U620 ( .A1(n555), .A2(n379), .ZN(n533) );
  NOR2_X1 U621 ( .A1(n533), .A2(n556), .ZN(n535) );
  XNOR2_X1 U622 ( .A(n535), .B(n534), .ZN(n539) );
  OR2_X1 U623 ( .A1(n537), .A2(n536), .ZN(n595) );
  INV_X1 U624 ( .A(n595), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U626 ( .A(KEYINPUT106), .B(n540), .ZN(n743) );
  NAND2_X1 U627 ( .A1(n541), .A2(n743), .ZN(n542) );
  XNOR2_X1 U628 ( .A(n542), .B(KEYINPUT75), .ZN(n554) );
  NAND2_X1 U629 ( .A1(n543), .A2(n664), .ZN(n544) );
  XNOR2_X1 U630 ( .A(KEYINPUT28), .B(n544), .ZN(n546) );
  NOR2_X1 U631 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U632 ( .A(n547), .B(KEYINPUT107), .ZN(n565) );
  INV_X1 U633 ( .A(n548), .ZN(n549) );
  OR2_X1 U634 ( .A1(n565), .A2(n549), .ZN(n550) );
  XNOR2_X1 U635 ( .A(n550), .B(KEYINPUT47), .ZN(n552) );
  INV_X1 U636 ( .A(n550), .ZN(n737) );
  NAND2_X1 U637 ( .A1(n737), .A2(n649), .ZN(n551) );
  NAND2_X1 U638 ( .A1(n552), .A2(n551), .ZN(n553) );
  AND2_X1 U639 ( .A1(n379), .A2(n555), .ZN(n557) );
  XNOR2_X1 U640 ( .A(n556), .B(KEYINPUT38), .ZN(n644) );
  NAND2_X1 U641 ( .A1(n557), .A2(n644), .ZN(n559) );
  XNOR2_X1 U642 ( .A(n559), .B(n558), .ZN(n576) );
  INV_X1 U643 ( .A(n576), .ZN(n561) );
  NAND2_X1 U644 ( .A1(n561), .A2(n736), .ZN(n563) );
  NAND2_X1 U645 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U646 ( .A1(n647), .A2(n648), .ZN(n564) );
  XNOR2_X1 U647 ( .A(n564), .B(KEYINPUT41), .ZN(n676) );
  NOR2_X1 U648 ( .A1(n565), .A2(n676), .ZN(n567) );
  XNOR2_X1 U649 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n566) );
  XNOR2_X1 U650 ( .A(n567), .B(n566), .ZN(n740) );
  NAND2_X1 U651 ( .A1(n742), .A2(n740), .ZN(n568) );
  XNOR2_X1 U652 ( .A(n568), .B(KEYINPUT46), .ZN(n571) );
  XOR2_X1 U653 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n573) );
  XNOR2_X1 U654 ( .A(n574), .B(n573), .ZN(n579) );
  NOR2_X1 U655 ( .A1(n576), .A2(n575), .ZN(n739) );
  NOR2_X1 U656 ( .A1(n577), .A2(n739), .ZN(n578) );
  NAND2_X1 U657 ( .A1(n579), .A2(n578), .ZN(n637) );
  XOR2_X1 U658 ( .A(n581), .B(n580), .Z(n583) );
  XNOR2_X1 U659 ( .A(n637), .B(n583), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n582), .A2(n679), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n583), .B(G227), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n584), .A2(G900), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n585), .A2(G953), .ZN(n586) );
  XNOR2_X1 U664 ( .A(n586), .B(KEYINPUT124), .ZN(n587) );
  NAND2_X1 U665 ( .A1(n588), .A2(n587), .ZN(G72) );
  INV_X1 U666 ( .A(G898), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n589), .A2(G953), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n636) );
  INV_X1 U669 ( .A(KEYINPUT102), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n652), .A2(n593), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n594), .B(KEYINPUT34), .ZN(n596) );
  NOR2_X1 U672 ( .A1(n717), .A2(KEYINPUT77), .ZN(n612) );
  INV_X1 U673 ( .A(n598), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n599), .A2(n656), .ZN(n600) );
  NOR2_X1 U675 ( .A1(n510), .A2(n600), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n604) );
  XNOR2_X1 U677 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n603) );
  XNOR2_X2 U678 ( .A(n604), .B(n603), .ZN(n700) );
  NOR2_X1 U679 ( .A1(n605), .A2(n664), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n346), .A2(n606), .ZN(n607) );
  NOR2_X2 U681 ( .A1(n608), .A2(n607), .ZN(n697) );
  INV_X1 U682 ( .A(KEYINPUT44), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n697), .A2(n609), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n700), .A2(n610), .ZN(n611) );
  NOR2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n614) );
  NOR2_X1 U686 ( .A1(KEYINPUT77), .A2(KEYINPUT44), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n627) );
  NOR2_X1 U688 ( .A1(n697), .A2(KEYINPUT44), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n700), .A2(n615), .ZN(n617) );
  INV_X1 U690 ( .A(KEYINPUT77), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n618), .A2(n342), .ZN(n625) );
  NOR2_X1 U693 ( .A1(n621), .A2(n649), .ZN(n622) );
  NOR2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U696 ( .A(n628), .B(KEYINPUT45), .ZN(n638) );
  NOR2_X1 U697 ( .A1(n343), .A2(G953), .ZN(n629) );
  XNOR2_X1 U698 ( .A(n629), .B(KEYINPUT123), .ZN(n634) );
  NAND2_X1 U699 ( .A1(G224), .A2(G953), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(KEYINPUT122), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n631), .B(KEYINPUT61), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n632), .A2(G898), .ZN(n633) );
  NAND2_X1 U703 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U704 ( .A(n636), .B(n635), .Z(G69) );
  NOR2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U706 ( .A1(KEYINPUT2), .A2(KEYINPUT72), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n640), .B(n639), .ZN(n642) );
  OR2_X1 U708 ( .A1(KEYINPUT2), .A2(KEYINPUT72), .ZN(n641) );
  NAND2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n687) );
  BUF_X1 U710 ( .A(n687), .Z(n684) );
  NOR2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U712 ( .A(n645), .B(KEYINPUT118), .ZN(n646) );
  NOR2_X1 U713 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U714 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U715 ( .A1(n651), .A2(n650), .ZN(n654) );
  INV_X1 U716 ( .A(n677), .ZN(n653) );
  NOR2_X1 U717 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U718 ( .A(KEYINPUT119), .B(n655), .Z(n672) );
  XOR2_X1 U719 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n659) );
  NAND2_X1 U720 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U721 ( .A(n659), .B(n658), .ZN(n666) );
  NAND2_X1 U722 ( .A1(n660), .A2(n346), .ZN(n661) );
  XNOR2_X1 U723 ( .A(n661), .B(KEYINPUT117), .ZN(n662) );
  XNOR2_X1 U724 ( .A(KEYINPUT50), .B(n662), .ZN(n663) );
  NOR2_X1 U725 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U726 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U727 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U728 ( .A(KEYINPUT51), .B(n669), .ZN(n670) );
  NOR2_X1 U729 ( .A1(n676), .A2(n670), .ZN(n671) );
  NOR2_X1 U730 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U731 ( .A(KEYINPUT52), .B(n673), .ZN(n675) );
  NOR2_X1 U732 ( .A1(n675), .A2(n674), .ZN(n682) );
  INV_X1 U733 ( .A(n676), .ZN(n678) );
  NAND2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n680) );
  NAND2_X1 U735 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U736 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U737 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U738 ( .A(KEYINPUT53), .B(n685), .Z(G75) );
  NOR2_X2 U739 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X2 U740 ( .A(n688), .B(KEYINPUT64), .ZN(n722) );
  NAND2_X1 U741 ( .A1(n722), .A2(G472), .ZN(n693) );
  XOR2_X1 U742 ( .A(KEYINPUT82), .B(KEYINPUT111), .Z(n689) );
  XNOR2_X1 U743 ( .A(n689), .B(KEYINPUT62), .ZN(n690) );
  XNOR2_X1 U744 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U745 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U746 ( .A1(n694), .A2(G953), .ZN(n720) );
  NAND2_X1 U747 ( .A1(n695), .A2(n720), .ZN(n696) );
  XNOR2_X1 U748 ( .A(n696), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U749 ( .A(G110), .B(KEYINPUT114), .Z(n698) );
  XNOR2_X1 U750 ( .A(n697), .B(n698), .ZN(G12) );
  XOR2_X1 U751 ( .A(G119), .B(KEYINPUT125), .Z(n699) );
  XNOR2_X1 U752 ( .A(n700), .B(n699), .ZN(G21) );
  NAND2_X1 U753 ( .A1(n722), .A2(G475), .ZN(n704) );
  XOR2_X1 U754 ( .A(KEYINPUT83), .B(KEYINPUT59), .Z(n701) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U756 ( .A(n704), .B(n703), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n705), .A2(n720), .ZN(n707) );
  XNOR2_X1 U758 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n707), .B(n706), .ZN(G60) );
  INV_X1 U760 ( .A(KEYINPUT56), .ZN(n716) );
  NAND2_X1 U761 ( .A1(n722), .A2(G210), .ZN(n713) );
  XOR2_X1 U762 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n710) );
  XNOR2_X1 U763 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n709) );
  XNOR2_X1 U764 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n708), .B(n711), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n714), .A2(n720), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n716), .B(n715), .ZN(G51) );
  XNOR2_X1 U769 ( .A(n342), .B(G122), .ZN(G24) );
  NAND2_X1 U770 ( .A1(n722), .A2(G217), .ZN(n718) );
  XOR2_X1 U771 ( .A(n719), .B(n718), .Z(n721) );
  INV_X1 U772 ( .A(n720), .ZN(n731) );
  NOR2_X1 U773 ( .A1(n721), .A2(n731), .ZN(G66) );
  AND2_X1 U774 ( .A1(n345), .A2(G478), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n725), .A2(n731), .ZN(G63) );
  NAND2_X1 U777 ( .A1(n345), .A2(G469), .ZN(n730) );
  XOR2_X1 U778 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n727) );
  XNOR2_X1 U779 ( .A(n727), .B(KEYINPUT58), .ZN(n728) );
  XNOR2_X1 U780 ( .A(n344), .B(n728), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n730), .B(n729), .ZN(n732) );
  NOR2_X1 U782 ( .A1(n732), .A2(n731), .ZN(G54) );
  XOR2_X1 U783 ( .A(G128), .B(KEYINPUT29), .Z(n735) );
  NAND2_X1 U784 ( .A1(n737), .A2(n733), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n735), .B(n734), .ZN(G30) );
  NAND2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n738), .B(G146), .ZN(G48) );
  XOR2_X1 U788 ( .A(G134), .B(n739), .Z(G36) );
  XNOR2_X1 U789 ( .A(G137), .B(n740), .ZN(n741) );
  XNOR2_X1 U790 ( .A(n741), .B(KEYINPUT126), .ZN(G39) );
  XNOR2_X1 U791 ( .A(n742), .B(G131), .ZN(G33) );
  XNOR2_X1 U792 ( .A(G143), .B(n743), .ZN(G45) );
endmodule

