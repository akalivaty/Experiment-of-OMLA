//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AND3_X1   g040(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(KEYINPUT67), .B2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n465), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n469), .A2(G136), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT68), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n468), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR3_X1   g058(.A1(new_n477), .A2(new_n480), .A3(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(KEYINPUT4), .B(G138), .C1(new_n466), .C2(new_n467), .ZN(new_n485));
  NAND2_X1  g060(.A1(G102), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G126), .B1(new_n466), .B2(new_n467), .ZN(new_n488));
  OR2_X1    g063(.A1(KEYINPUT69), .A2(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(KEYINPUT69), .A2(G114), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n489), .A2(G2104), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n481), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n481), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(KEYINPUT4), .B1(new_n461), .B2(new_n493), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n487), .A2(new_n492), .A3(new_n494), .ZN(G164));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(KEYINPUT70), .A2(G651), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(KEYINPUT6), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT71), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n499), .A2(new_n505), .A3(KEYINPUT6), .A4(new_n500), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n496), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT70), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT70), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NOR3_X1   g086(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n506), .B1(new_n512), .B2(new_n502), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(G88), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(new_n516), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n509), .A2(new_n510), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n508), .A2(new_n517), .A3(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  AOI21_X1  g102(.A(new_n520), .B1(new_n504), .B2(new_n506), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT73), .B(G89), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n507), .A2(G51), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n516), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n531), .A3(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G64), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n520), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n507), .A2(G52), .B1(new_n541), .B2(new_n524), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n528), .A2(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G43), .Z(new_n546));
  NAND2_X1  g121(.A1(new_n507), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n528), .A2(G81), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n523), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT76), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n514), .B2(new_n515), .ZN(new_n561));
  AND2_X1   g136(.A1(G78), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g140(.A(KEYINPUT77), .B(G651), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(new_n528), .B2(G91), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n507), .A2(new_n568), .A3(G53), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n568), .B1(new_n507), .B2(G53), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n498), .B1(new_n520), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n507), .B2(G49), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n528), .A2(KEYINPUT78), .A3(G87), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT78), .B1(new_n528), .B2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n520), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n507), .A2(G48), .B1(new_n581), .B2(new_n524), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n513), .A2(G86), .A3(new_n516), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n528), .A2(new_n585), .A3(G86), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n528), .A2(G85), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n513), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT80), .B(G47), .Z(new_n591));
  OAI221_X1 g166(.A(new_n588), .B1(new_n523), .B2(new_n589), .C1(new_n590), .C2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  OAI21_X1  g168(.A(G54), .B1(new_n507), .B2(KEYINPUT81), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n513), .A2(KEYINPUT81), .A3(G543), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n594), .A2(new_n595), .B1(new_n498), .B2(new_n596), .ZN(new_n597));
  AND4_X1   g172(.A1(KEYINPUT10), .A2(new_n513), .A3(G92), .A4(new_n516), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT10), .B1(new_n528), .B2(G92), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n593), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  OAI21_X1  g184(.A(KEYINPUT82), .B1(new_n552), .B2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n601), .A2(new_n608), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  MUX2_X1   g187(.A(KEYINPUT82), .B(new_n610), .S(new_n612), .Z(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n461), .A2(new_n472), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT84), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT13), .Z(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n469), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n482), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n481), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND3_X1  g202(.A1(new_n620), .A2(new_n621), .A3(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT87), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT86), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XOR2_X1   g215(.A(G1341), .B(G1348), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  OAI21_X1  g219(.A(G14), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(KEYINPUT17), .ZN(new_n653));
  INV_X1    g228(.A(new_n647), .ZN(new_n654));
  INV_X1    g229(.A(new_n648), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n650), .A3(new_n655), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(new_n649), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n652), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT88), .B(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n664), .A2(new_n665), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n663), .A2(new_n666), .A3(new_n670), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1981), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(G229));
  INV_X1    g256(.A(KEYINPUT104), .ZN(new_n682));
  NAND2_X1  g257(.A1(G305), .A2(G16), .ZN(new_n683));
  INV_X1    g258(.A(G6), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(G16), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(KEYINPUT92), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT92), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n683), .A2(new_n689), .A3(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT32), .B(G1981), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n691), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n689), .B1(new_n683), .B2(new_n686), .ZN(new_n694));
  AOI211_X1 g269(.A(KEYINPUT92), .B(new_n685), .C1(G305), .C2(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT95), .ZN(new_n700));
  NAND2_X1  g275(.A1(G303), .A2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT94), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n700), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  AOI211_X1 g281(.A(KEYINPUT95), .B(new_n704), .C1(G303), .C2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(G1971), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g283(.A1(new_n528), .A2(G88), .B1(new_n522), .B2(new_n524), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n702), .B1(new_n709), .B2(new_n508), .ZN(new_n710));
  OAI21_X1  g285(.A(KEYINPUT95), .B1(new_n710), .B2(new_n704), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n701), .A2(new_n700), .A3(new_n705), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n702), .A2(G23), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G288), .B2(G16), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI211_X1 g294(.A(KEYINPUT33), .B(new_n716), .C1(G288), .C2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(G1976), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n577), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n528), .A2(KEYINPUT78), .A3(G87), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n702), .B1(new_n724), .B2(new_n575), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT33), .B1(new_n725), .B2(new_n716), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n717), .A2(new_n718), .ZN(new_n727));
  INV_X1    g302(.A(G1976), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n715), .B1(new_n721), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n692), .A2(new_n696), .A3(KEYINPUT93), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n699), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT34), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT34), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n699), .A2(new_n730), .A3(new_n734), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n469), .A2(G131), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n482), .A2(G119), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n481), .A2(G107), .ZN(new_n738));
  OAI21_X1  g313(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n736), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G25), .B(new_n740), .S(G29), .Z(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT35), .B(G1991), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT91), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n741), .B(new_n743), .Z(new_n744));
  AND2_X1   g319(.A1(new_n702), .A2(G24), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G290), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1986), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n747), .B2(new_n746), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n733), .A2(new_n735), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(KEYINPUT36), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n733), .A2(new_n752), .A3(new_n735), .A4(new_n749), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G34), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n474), .B2(new_n757), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT100), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n757), .A2(G35), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G162), .B2(new_n757), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT29), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n766), .B(new_n763), .C1(G162), .C2(new_n757), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n757), .A2(G33), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n469), .A2(G139), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT97), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n461), .A2(G127), .ZN(new_n773));
  INV_X1    g348(.A(G115), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n471), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n776));
  NAND2_X1  g351(.A1(G103), .A2(G2104), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G2105), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n481), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n775), .A2(G2105), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n772), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n770), .B1(new_n782), .B2(G29), .ZN(new_n783));
  INV_X1    g358(.A(G2072), .ZN(new_n784));
  AOI22_X1  g359(.A1(G2090), .A2(new_n768), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n757), .A2(G32), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n469), .A2(G141), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n482), .A2(G129), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT26), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n791), .A2(new_n792), .B1(G105), .B2(new_n472), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n786), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT27), .B(G1996), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT31), .B(G11), .Z(new_n799));
  INV_X1    g374(.A(G28), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(KEYINPUT30), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT102), .Z(new_n802));
  AOI21_X1  g377(.A(G29), .B1(new_n800), .B2(KEYINPUT30), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n798), .B(new_n804), .C1(new_n757), .C2(new_n626), .ZN(new_n805));
  AOI211_X1 g380(.A(new_n797), .B(new_n805), .C1(new_n760), .C2(new_n759), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n757), .A2(G27), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G164), .B2(new_n757), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2078), .ZN(new_n809));
  NOR2_X1   g384(.A1(G171), .A2(new_n702), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G5), .B2(new_n702), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n762), .A2(new_n785), .A3(new_n806), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G16), .A2(G19), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n552), .B2(G16), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1341), .Z(new_n817));
  NAND2_X1  g392(.A1(new_n702), .A2(G21), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G168), .B2(new_n702), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G1966), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n757), .A2(G26), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT28), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n469), .A2(G140), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n482), .A2(G128), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n481), .A2(G116), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n823), .B1(new_n828), .B2(G29), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT96), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2067), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n811), .A2(new_n812), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n819), .A2(G1966), .ZN(new_n833));
  NOR4_X1   g408(.A1(new_n821), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n702), .A2(G20), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT23), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n605), .B2(new_n702), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1956), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n601), .A2(G16), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G4), .B2(G16), .ZN(new_n840));
  INV_X1    g415(.A(G1348), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n838), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OR3_X1    g419(.A1(new_n783), .A2(KEYINPUT101), .A3(new_n784), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT101), .B1(new_n783), .B2(new_n784), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n768), .B2(G2090), .ZN(new_n848));
  INV_X1    g423(.A(G2090), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n765), .A2(KEYINPUT103), .A3(new_n849), .A4(new_n767), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n845), .A2(new_n846), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n814), .A2(new_n834), .A3(new_n844), .A4(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n682), .B1(new_n754), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g429(.A(KEYINPUT104), .B(new_n852), .C1(new_n751), .C2(new_n753), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(G311));
  NAND2_X1  g431(.A1(new_n754), .A2(new_n853), .ZN(G150));
  AOI22_X1  g432(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT105), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(KEYINPUT105), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n524), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n528), .A2(G93), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n507), .A2(G55), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G860), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT37), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n601), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n551), .A2(KEYINPUT106), .ZN(new_n869));
  INV_X1    g444(.A(new_n864), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n551), .A2(KEYINPUT106), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n869), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n868), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(KEYINPUT39), .ZN(new_n877));
  INV_X1    g452(.A(G860), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n876), .B2(KEYINPUT39), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n866), .B1(new_n877), .B2(new_n879), .ZN(G145));
  INV_X1    g455(.A(G37), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n626), .B(new_n474), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(G162), .Z(new_n883));
  NAND2_X1  g458(.A1(KEYINPUT4), .A2(G138), .ZN(new_n884));
  NAND2_X1  g459(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT3), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(KEYINPUT67), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n486), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n481), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G126), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n887), .B2(new_n888), .ZN(new_n893));
  INV_X1    g468(.A(new_n490), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(KEYINPUT69), .B2(G114), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(G2105), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n494), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n891), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n828), .B(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n794), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n781), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n782), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n902), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n482), .A2(G130), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n481), .A2(G118), .ZN(new_n909));
  OAI21_X1  g484(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(G142), .B2(new_n469), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(new_n740), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n618), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n907), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n904), .A2(new_n914), .A3(new_n906), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n883), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n883), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n907), .A2(KEYINPUT107), .A3(new_n914), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n881), .B(new_n917), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g498(.A1(new_n597), .A2(new_n600), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(G299), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n601), .A2(new_n605), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n874), .A2(new_n611), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n874), .A2(new_n611), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n925), .A2(new_n926), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT41), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n930), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(G288), .B(G305), .ZN(new_n940));
  XNOR2_X1  g515(.A(G290), .B(G303), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(KEYINPUT108), .B2(KEYINPUT42), .ZN(new_n943));
  OAI221_X1 g518(.A(new_n930), .B1(KEYINPUT108), .B2(KEYINPUT42), .C1(new_n931), .C2(new_n936), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n939), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n870), .A2(G868), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(G331));
  XNOR2_X1  g525(.A(G168), .B(G301), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n874), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n951), .B1(new_n872), .B2(new_n873), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(KEYINPUT109), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n869), .A2(new_n871), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n864), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n956), .B1(new_n960), .B2(new_n951), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n953), .B1(new_n955), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n933), .A2(new_n935), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n960), .A2(new_n951), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n964), .A2(new_n934), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n962), .A2(new_n963), .B1(new_n954), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G37), .B1(new_n966), .B2(new_n942), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n953), .A2(new_n927), .A3(new_n954), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n954), .A2(KEYINPUT109), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n960), .A2(new_n956), .A3(new_n951), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n964), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n968), .B1(new_n971), .B2(new_n936), .ZN(new_n972));
  INV_X1    g547(.A(new_n942), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT43), .B1(new_n967), .B2(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n942), .B(new_n968), .C1(new_n971), .C2(new_n936), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n881), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n927), .A2(KEYINPUT110), .A3(new_n932), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n953), .A2(new_n954), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n978), .B(new_n979), .C1(new_n963), .C2(KEYINPUT110), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n965), .B1(new_n961), .B2(new_n955), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n942), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n977), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n975), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n967), .B2(new_n974), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n977), .A2(new_n982), .A3(KEYINPUT43), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n989), .ZN(G397));
  AOI21_X1  g565(.A(new_n481), .B1(new_n462), .B2(new_n463), .ZN(new_n991));
  INV_X1    g566(.A(G137), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n468), .A2(new_n992), .A3(G2105), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  INV_X1    g569(.A(new_n473), .ZN(new_n995));
  NOR4_X1   g570(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n899), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G1996), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT46), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1000), .B(KEYINPUT112), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n828), .B(G2067), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n901), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1003), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1004), .B1(new_n1009), .B2(new_n901), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n1003), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1001), .A2(new_n901), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT113), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n740), .A2(new_n743), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g591(.A1(new_n828), .A2(G2067), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1008), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n740), .A2(new_n743), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1003), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n1000), .A2(G290), .A3(G1986), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  AOI211_X1 g599(.A(new_n1007), .B(new_n1018), .C1(new_n1021), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G303), .A2(G8), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT55), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n492), .A2(new_n494), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n1028), .B2(new_n891), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n996), .B1(new_n1029), .B2(KEYINPUT45), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n899), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n713), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n465), .A2(G40), .A3(new_n470), .A4(new_n473), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n998), .B2(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n899), .A2(new_n1036), .A3(new_n997), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n849), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(KEYINPUT117), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G8), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1027), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1033), .A2(KEYINPUT115), .A3(new_n1038), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1027), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(G8), .A4(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1029), .B2(new_n996), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(G288), .B2(new_n728), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G288), .A2(new_n728), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1052), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n582), .A2(new_n583), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G1981), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n582), .A2(new_n584), .A3(new_n1059), .A4(new_n586), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1058), .A2(new_n1060), .A3(KEYINPUT49), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT49), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1050), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1056), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1042), .A2(new_n1048), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n996), .A3(new_n1037), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1034), .B1(new_n998), .B2(new_n999), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1031), .A3(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n567), .B(new_n1074), .C1(new_n570), .C2(new_n571), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1074), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G299), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1070), .A2(new_n1073), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1077), .A2(new_n1080), .A3(new_n1075), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1077), .B2(new_n1075), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n998), .A2(new_n1034), .A3(G2067), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1085), .B1(new_n1068), .B2(new_n841), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1084), .B1(new_n1086), .B2(new_n924), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1086), .A2(new_n1084), .A3(new_n924), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1078), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1071), .A2(new_n1031), .A3(new_n1072), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1956), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1077), .A2(new_n1075), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1091), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1083), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1348), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  NOR4_X1   g675(.A1(new_n1099), .A2(new_n601), .A3(new_n1100), .A4(new_n1085), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n924), .B1(new_n1086), .B2(KEYINPUT60), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1099), .B2(new_n1085), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n999), .B1(G164), .B2(G1384), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1105), .A2(new_n1009), .A3(new_n1031), .A4(new_n996), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n998), .B2(new_n1034), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1106), .A2(KEYINPUT123), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT123), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n552), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT59), .B(new_n552), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1098), .A2(new_n1104), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1079), .A2(KEYINPUT124), .A3(new_n1095), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1091), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1079), .A2(new_n1095), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT124), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1090), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1071), .A2(new_n1031), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(G2078), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1068), .A2(new_n812), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1029), .A2(KEYINPUT118), .A3(KEYINPUT45), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1031), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1071), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OR2_X1    g704(.A1(new_n1122), .A2(G2078), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1124), .B(new_n1125), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(G301), .B(KEYINPUT54), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1123), .A2(new_n1130), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1132), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1134), .A2(new_n1135), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n1139));
  INV_X1    g714(.A(G1966), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1129), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1035), .A2(new_n760), .A3(new_n1037), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1139), .B(new_n1049), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G286), .A2(G8), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT125), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1138), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1145), .B1(KEYINPUT126), .B2(new_n1138), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G8), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1147), .A2(new_n1149), .B1(new_n1148), .B2(new_n1145), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1137), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1121), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1049), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT126), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1144), .B(KEYINPUT125), .Z(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT51), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1148), .A2(new_n1145), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1139), .B2(KEYINPUT51), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n1153), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT62), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1146), .A2(new_n1150), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1160), .A2(new_n1162), .A3(G171), .A4(new_n1131), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1066), .B1(new_n1152), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1065), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1060), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n724), .A2(new_n728), .A3(new_n575), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT116), .Z(new_n1168));
  OR2_X1    g743(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1165), .A2(new_n1048), .B1(new_n1170), .B2(new_n1063), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1049), .B(G286), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1042), .A2(new_n1065), .A3(new_n1048), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1149), .A2(new_n1174), .A3(G286), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1045), .A2(new_n1046), .A3(G8), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1027), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1176), .A2(new_n1178), .A3(new_n1048), .A4(new_n1065), .ZN(new_n1179));
  AOI211_X1 g754(.A(KEYINPUT119), .B(new_n1171), .C1(new_n1175), .C2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT119), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1175), .A2(new_n1179), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1171), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1164), .A2(new_n1180), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(G290), .A2(G1986), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1022), .B1(new_n1000), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT111), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1021), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT114), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1025), .B1(new_n1185), .B2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g767(.A1(new_n459), .A2(G227), .ZN(new_n1194));
  NOR3_X1   g768(.A1(G229), .A2(G401), .A3(new_n1194), .ZN(new_n1195));
  OAI211_X1 g769(.A(new_n922), .B(new_n1195), .C1(new_n987), .C2(new_n988), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


