

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n384) );
  XNOR2_X1 U326 ( .A(n385), .B(n384), .ZN(n386) );
  NOR2_X1 U327 ( .A1(n578), .A2(n379), .ZN(n380) );
  XNOR2_X1 U328 ( .A(n331), .B(KEYINPUT32), .ZN(n332) );
  XNOR2_X1 U329 ( .A(n351), .B(n332), .ZN(n336) );
  NOR2_X1 U330 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U331 ( .A(n368), .B(n367), .ZN(n370) );
  XNOR2_X1 U332 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U333 ( .A(KEYINPUT36), .B(n543), .Z(n585) );
  NOR2_X1 U334 ( .A1(n523), .A2(n452), .ZN(n566) );
  XOR2_X1 U335 ( .A(n311), .B(n406), .Z(n523) );
  XNOR2_X1 U336 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n456) );
  XNOR2_X1 U337 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n294) );
  XNOR2_X1 U339 ( .A(G43GAT), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U341 ( .A(KEYINPUT65), .B(G176GAT), .Z(n296) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(G15GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U344 ( .A(n298), .B(n297), .Z(n303) );
  XOR2_X1 U345 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n300) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U348 ( .A(KEYINPUT89), .B(n301), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U350 ( .A(G120GAT), .B(G71GAT), .Z(n340) );
  XOR2_X1 U351 ( .A(n304), .B(n340), .Z(n307) );
  XOR2_X1 U352 ( .A(G190GAT), .B(G134GAT), .Z(n364) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n305), .B(G127GAT), .ZN(n423) );
  XNOR2_X1 U355 ( .A(n364), .B(n423), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U357 ( .A(KEYINPUT18), .B(KEYINPUT88), .Z(n309) );
  XNOR2_X1 U358 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U360 ( .A(KEYINPUT19), .B(n310), .Z(n406) );
  XOR2_X1 U361 ( .A(G43GAT), .B(G29GAT), .Z(n313) );
  XNOR2_X1 U362 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U364 ( .A(n314), .B(KEYINPUT70), .Z(n316) );
  XNOR2_X1 U365 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n375) );
  XOR2_X1 U367 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n318) );
  XNOR2_X1 U368 ( .A(KEYINPUT71), .B(KEYINPUT68), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n375), .B(n319), .ZN(n327) );
  XOR2_X1 U371 ( .A(G141GAT), .B(G22GAT), .Z(n437) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(G197GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n320), .B(G8GAT), .ZN(n398) );
  XOR2_X1 U374 ( .A(n437), .B(n398), .Z(n322) );
  NAND2_X1 U375 ( .A1(G229GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U377 ( .A(G15GAT), .B(G1GAT), .Z(n348) );
  XOR2_X1 U378 ( .A(n323), .B(n348), .Z(n325) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n573) );
  XNOR2_X1 U382 ( .A(n573), .B(KEYINPUT72), .ZN(n564) );
  INV_X1 U383 ( .A(KEYINPUT118), .ZN(n381) );
  XOR2_X1 U384 ( .A(KEYINPUT31), .B(KEYINPUT77), .Z(n329) );
  XNOR2_X1 U385 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n344) );
  XNOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n330), .B(KEYINPUT73), .ZN(n351) );
  AND2_X1 U389 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XOR2_X1 U390 ( .A(G176GAT), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U391 ( .A(KEYINPUT33), .B(n401), .ZN(n334) );
  XOR2_X1 U392 ( .A(G148GAT), .B(G78GAT), .Z(n432) );
  XNOR2_X1 U393 ( .A(G204GAT), .B(n432), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U396 ( .A(G92GAT), .B(KEYINPUT74), .Z(n338) );
  XNOR2_X1 U397 ( .A(G99GAT), .B(G85GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U399 ( .A(G106GAT), .B(n339), .Z(n369) );
  XNOR2_X1 U400 ( .A(n340), .B(n369), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U402 ( .A(n344), .B(n343), .Z(n458) );
  INV_X1 U403 ( .A(n458), .ZN(n578) );
  XOR2_X1 U404 ( .A(G155GAT), .B(G211GAT), .Z(n346) );
  XNOR2_X1 U405 ( .A(G183GAT), .B(G127GAT), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U407 ( .A(n347), .B(G78GAT), .Z(n350) );
  XNOR2_X1 U408 ( .A(n348), .B(G22GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U410 ( .A(n351), .B(KEYINPUT12), .Z(n353) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U413 ( .A(n355), .B(n354), .Z(n363) );
  XOR2_X1 U414 ( .A(KEYINPUT83), .B(G64GAT), .Z(n357) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G71GAT), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U417 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n359) );
  XNOR2_X1 U418 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U421 ( .A(n363), .B(n362), .Z(n581) );
  INV_X1 U422 ( .A(n581), .ZN(n491) );
  XOR2_X1 U423 ( .A(G218GAT), .B(G162GAT), .Z(n433) );
  XOR2_X1 U424 ( .A(n364), .B(n433), .Z(n368) );
  XOR2_X1 U425 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n366) );
  XNOR2_X1 U426 ( .A(KEYINPUT79), .B(KEYINPUT66), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n372) );
  NAND2_X1 U429 ( .A1(G232GAT), .A2(G233GAT), .ZN(n371) );
  XOR2_X1 U430 ( .A(n372), .B(n371), .Z(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n377) );
  XNOR2_X1 U432 ( .A(n375), .B(KEYINPUT9), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n559) );
  XNOR2_X1 U434 ( .A(KEYINPUT80), .B(n559), .ZN(n543) );
  NOR2_X1 U435 ( .A1(n491), .A2(n585), .ZN(n378) );
  XOR2_X1 U436 ( .A(KEYINPUT45), .B(n378), .Z(n379) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  NOR2_X1 U438 ( .A1(n564), .A2(n382), .ZN(n391) );
  XNOR2_X1 U439 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n383) );
  XOR2_X1 U440 ( .A(n578), .B(n383), .Z(n550) );
  NAND2_X1 U441 ( .A1(n550), .A2(n573), .ZN(n385) );
  NAND2_X1 U442 ( .A1(n386), .A2(n491), .ZN(n387) );
  XOR2_X1 U443 ( .A(KEYINPUT117), .B(n387), .Z(n388) );
  NOR2_X1 U444 ( .A1(n559), .A2(n388), .ZN(n389) );
  XOR2_X1 U445 ( .A(n389), .B(KEYINPUT47), .Z(n390) );
  XNOR2_X1 U446 ( .A(n392), .B(KEYINPUT48), .ZN(n529) );
  XOR2_X1 U447 ( .A(KEYINPUT99), .B(G190GAT), .Z(n394) );
  NAND2_X1 U448 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n397) );
  XOR2_X1 U450 ( .A(G204GAT), .B(G211GAT), .Z(n396) );
  XNOR2_X1 U451 ( .A(KEYINPUT91), .B(KEYINPUT21), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n442) );
  XOR2_X1 U453 ( .A(n397), .B(n442), .Z(n400) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(n398), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U456 ( .A(n402), .B(n401), .Z(n404) );
  XNOR2_X1 U457 ( .A(G218GAT), .B(G92GAT), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n521) );
  NOR2_X1 U460 ( .A1(n529), .A2(n521), .ZN(n407) );
  XNOR2_X1 U461 ( .A(KEYINPUT54), .B(n407), .ZN(n572) );
  NAND2_X1 U462 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XOR2_X1 U463 ( .A(G148GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G141GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U466 ( .A(G134GAT), .B(G85GAT), .Z(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n429) );
  XOR2_X1 U469 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n415) );
  XNOR2_X1 U470 ( .A(KEYINPUT5), .B(KEYINPUT98), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U472 ( .A(KEYINPUT96), .B(G57GAT), .Z(n417) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G120GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U475 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT95), .B(KEYINPUT97), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U479 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n422), .B(KEYINPUT2), .ZN(n440) );
  XNOR2_X1 U481 ( .A(n423), .B(n440), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n568) );
  XOR2_X1 U485 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n431) );
  XNOR2_X1 U486 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n448) );
  XOR2_X1 U488 ( .A(G106GAT), .B(n432), .Z(n435) );
  XNOR2_X1 U489 ( .A(G50GAT), .B(n433), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n446) );
  XOR2_X1 U492 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n439) );
  NAND2_X1 U493 ( .A1(G228GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U495 ( .A(n441), .B(n440), .Z(n444) );
  XNOR2_X1 U496 ( .A(G197GAT), .B(n442), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n467) );
  INV_X1 U500 ( .A(n467), .ZN(n449) );
  AND2_X1 U501 ( .A1(n568), .A2(n449), .ZN(n450) );
  AND2_X1 U502 ( .A1(n572), .A2(n450), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NAND2_X1 U504 ( .A1(n566), .A2(n550), .ZN(n455) );
  XOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  XNOR2_X1 U506 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  NAND2_X1 U508 ( .A1(n543), .A2(n566), .ZN(n457) );
  NAND2_X1 U509 ( .A1(n458), .A2(n564), .ZN(n494) );
  XOR2_X1 U510 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n460) );
  OR2_X1 U511 ( .A1(n543), .A2(n491), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n460), .B(n459), .ZN(n476) );
  INV_X1 U513 ( .A(n523), .ZN(n533) );
  XOR2_X1 U514 ( .A(KEYINPUT27), .B(KEYINPUT100), .Z(n461) );
  XOR2_X1 U515 ( .A(n521), .B(n461), .Z(n470) );
  INV_X1 U516 ( .A(n470), .ZN(n531) );
  XOR2_X1 U517 ( .A(KEYINPUT28), .B(n467), .Z(n534) );
  NAND2_X1 U518 ( .A1(n531), .A2(n534), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n533), .A2(n462), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n568), .A2(n463), .ZN(n474) );
  NOR2_X1 U521 ( .A1(n523), .A2(n521), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n467), .A2(n464), .ZN(n465) );
  XNOR2_X1 U523 ( .A(KEYINPUT25), .B(n465), .ZN(n466) );
  NAND2_X1 U524 ( .A1(n466), .A2(n568), .ZN(n472) );
  XOR2_X1 U525 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n469) );
  NAND2_X1 U526 ( .A1(n523), .A2(n467), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n469), .B(n468), .ZN(n570) );
  NOR2_X1 U528 ( .A1(n470), .A2(n570), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT102), .B(n475), .ZN(n490) );
  NAND2_X1 U532 ( .A1(n476), .A2(n490), .ZN(n508) );
  OR2_X1 U533 ( .A1(n494), .A2(n508), .ZN(n488) );
  NOR2_X1 U534 ( .A1(n568), .A2(n488), .ZN(n481) );
  XOR2_X1 U535 ( .A(KEYINPUT34), .B(KEYINPUT105), .Z(n478) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(KEYINPUT104), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U538 ( .A(KEYINPUT103), .B(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  NOR2_X1 U540 ( .A1(n521), .A2(n488), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n484), .ZN(G1325GAT) );
  NOR2_X1 U544 ( .A1(n523), .A2(n488), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT108), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U547 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n534), .A2(n488), .ZN(n489) );
  XOR2_X1 U549 ( .A(G22GAT), .B(n489), .Z(G1327GAT) );
  XNOR2_X1 U550 ( .A(KEYINPUT110), .B(KEYINPUT39), .ZN(n498) );
  NAND2_X1 U551 ( .A1(n491), .A2(n490), .ZN(n492) );
  NOR2_X1 U552 ( .A1(n492), .A2(n585), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT37), .ZN(n519) );
  NOR2_X1 U554 ( .A1(n519), .A2(n494), .ZN(n496) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(KEYINPUT109), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(n503) );
  NOR2_X1 U557 ( .A1(n568), .A2(n503), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n503), .A2(n521), .ZN(n500) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n500), .Z(G1329GAT) );
  NOR2_X1 U562 ( .A1(n523), .A2(n503), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT40), .B(n501), .Z(n502) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  NOR2_X1 U565 ( .A1(n503), .A2(n534), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT111), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  INV_X1 U568 ( .A(n550), .ZN(n506) );
  NOR2_X1 U569 ( .A1(n506), .A2(n573), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(KEYINPUT113), .ZN(n518) );
  OR2_X1 U571 ( .A1(n518), .A2(n508), .ZN(n514) );
  NOR2_X1 U572 ( .A1(n568), .A2(n514), .ZN(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n511), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n521), .A2(n514), .ZN(n512) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n523), .A2(n514), .ZN(n513) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n513), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n534), .A2(n514), .ZN(n516) );
  XNOR2_X1 U581 ( .A(KEYINPUT114), .B(KEYINPUT43), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(n517), .ZN(G1335GAT) );
  OR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U585 ( .A1(n568), .A2(n526), .ZN(n520) );
  XOR2_X1 U586 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n526), .ZN(n522) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n526), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U592 ( .A1(n534), .A2(n526), .ZN(n527) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(n527), .Z(n528) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(KEYINPUT120), .ZN(n537) );
  NOR2_X1 U596 ( .A1(n568), .A2(n529), .ZN(n530) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(KEYINPUT119), .B(n532), .ZN(n552) );
  AND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U600 ( .A1(n552), .A2(n535), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n544), .A2(n564), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1340GAT) );
  XNOR2_X1 U603 ( .A(KEYINPUT121), .B(KEYINPUT49), .ZN(n539) );
  AND2_X1 U604 ( .A1(n544), .A2(n550), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(G120GAT), .B(n540), .Z(G1341GAT) );
  NAND2_X1 U607 ( .A1(n581), .A2(n544), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n547), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT123), .Z(n549) );
  INV_X1 U615 ( .A(n570), .ZN(n551) );
  AND2_X1 U616 ( .A1(n551), .A2(n552), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n560), .A2(n573), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  AND2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n581), .A2(n560), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT124), .ZN(n558) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n558), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n562) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n566), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n581), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT127), .Z(n575) );
  INV_X1 U636 ( .A(n568), .ZN(n569) );
  NOR2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  AND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n583), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n583), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U648 ( .A(n583), .ZN(n584) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

