

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n779), .A2(n778), .ZN(n780) );
  AND2_X1 U550 ( .A1(n759), .A2(n758), .ZN(n760) );
  AND2_X1 U551 ( .A1(n733), .A2(G8), .ZN(n689) );
  XOR2_X2 U552 ( .A(KEYINPUT64), .B(G2104), .Z(n523) );
  NAND2_X1 U553 ( .A1(n871), .A2(G101), .ZN(n529) );
  NOR2_X2 U554 ( .A1(n535), .A2(n534), .ZN(G160) );
  XOR2_X1 U555 ( .A(KEYINPUT74), .B(n574), .Z(n516) );
  NOR2_X1 U556 ( .A1(n748), .A2(n724), .ZN(n517) );
  XOR2_X1 U557 ( .A(n745), .B(n744), .Z(n518) );
  INV_X1 U558 ( .A(G8), .ZN(n724) );
  AND2_X1 U559 ( .A1(n692), .A2(n691), .ZN(n718) );
  NOR2_X1 U560 ( .A1(G1966), .A2(n768), .ZN(n750) );
  INV_X1 U561 ( .A(KEYINPUT32), .ZN(n744) );
  XNOR2_X1 U562 ( .A(n753), .B(KEYINPUT101), .ZN(n754) );
  NAND2_X1 U563 ( .A1(n518), .A2(n754), .ZN(n770) );
  XNOR2_X1 U564 ( .A(n689), .B(KEYINPUT95), .ZN(n768) );
  NOR2_X1 U565 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n692) );
  NOR2_X1 U567 ( .A1(G543), .A2(n541), .ZN(n536) );
  XOR2_X1 U568 ( .A(KEYINPUT15), .B(n578), .Z(n702) );
  NOR2_X1 U569 ( .A1(G651), .A2(n648), .ZN(n643) );
  XNOR2_X1 U570 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U571 ( .A1(n523), .A2(G2105), .ZN(n519) );
  XNOR2_X2 U572 ( .A(n519), .B(KEYINPUT65), .ZN(n598) );
  NAND2_X1 U573 ( .A1(n598), .A2(G126), .ZN(n522) );
  NOR2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n520), .Z(n870) );
  NAND2_X1 U576 ( .A1(n870), .A2(G138), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n874) );
  NAND2_X1 U579 ( .A1(G114), .A2(n874), .ZN(n525) );
  NOR2_X4 U580 ( .A1(G2105), .A2(n523), .ZN(n871) );
  NAND2_X1 U581 ( .A1(G102), .A2(n871), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n527), .A2(n526), .ZN(G164) );
  NAND2_X1 U584 ( .A1(n870), .A2(G137), .ZN(n531) );
  INV_X1 U585 ( .A(KEYINPUT23), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U587 ( .A1(G125), .A2(n598), .ZN(n533) );
  NAND2_X1 U588 ( .A1(G113), .A2(n874), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  NAND2_X1 U591 ( .A1(G51), .A2(n643), .ZN(n538) );
  INV_X1 U592 ( .A(G651), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT1), .B(n536), .Z(n647) );
  NAND2_X1 U594 ( .A1(G63), .A2(n647), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U596 ( .A(KEYINPUT6), .B(n539), .ZN(n547) );
  NOR2_X1 U597 ( .A1(G543), .A2(G651), .ZN(n635) );
  NAND2_X1 U598 ( .A1(n635), .A2(G89), .ZN(n540) );
  XNOR2_X1 U599 ( .A(n540), .B(KEYINPUT4), .ZN(n543) );
  NOR2_X1 U600 ( .A1(n648), .A2(n541), .ZN(n634) );
  NAND2_X1 U601 ( .A1(G76), .A2(n634), .ZN(n542) );
  NAND2_X1 U602 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U603 ( .A(KEYINPUT75), .B(n544), .ZN(n545) );
  XNOR2_X1 U604 ( .A(KEYINPUT5), .B(n545), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(n548), .Z(G168) );
  XNOR2_X1 U607 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n553) );
  NAND2_X1 U608 ( .A1(G77), .A2(n634), .ZN(n550) );
  NAND2_X1 U609 ( .A1(G90), .A2(n635), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U611 ( .A(n551), .B(KEYINPUT9), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n553), .B(n552), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G52), .A2(n643), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G64), .A2(n647), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U616 ( .A1(n557), .A2(n556), .ZN(G171) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U621 ( .A(n558), .B(KEYINPUT10), .ZN(n559) );
  XNOR2_X1 U622 ( .A(KEYINPUT70), .B(n559), .ZN(G223) );
  INV_X1 U623 ( .A(G223), .ZN(n820) );
  NAND2_X1 U624 ( .A1(n820), .A2(G567), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U626 ( .A1(G81), .A2(n635), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT71), .B(n561), .Z(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G68), .A2(n634), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT13), .B(n565), .ZN(n571) );
  NAND2_X1 U632 ( .A1(G43), .A2(n643), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT72), .B(n566), .Z(n569) );
  NAND2_X1 U634 ( .A1(n647), .A2(G56), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(n567), .Z(n568) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n944) );
  INV_X1 U638 ( .A(G860), .ZN(n608) );
  OR2_X1 U639 ( .A1(n944), .A2(n608), .ZN(G153) );
  XNOR2_X1 U640 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G868), .A2(G301), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n643), .A2(G54), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G79), .A2(n634), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G92), .A2(n635), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n647), .A2(G66), .ZN(n574) );
  NOR2_X1 U647 ( .A1(n575), .A2(n516), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n578) );
  INV_X1 U649 ( .A(G868), .ZN(n660) );
  NAND2_X1 U650 ( .A1(n702), .A2(n660), .ZN(n579) );
  NAND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G91), .A2(n635), .ZN(n582) );
  NAND2_X1 U653 ( .A1(G53), .A2(n643), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G78), .A2(n634), .ZN(n583) );
  XNOR2_X1 U656 ( .A(KEYINPUT69), .B(n583), .ZN(n584) );
  NOR2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n647), .A2(G65), .ZN(n586) );
  NAND2_X1 U659 ( .A1(n587), .A2(n586), .ZN(G299) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n588), .B(KEYINPUT76), .ZN(n590) );
  NOR2_X1 U662 ( .A1(n660), .A2(G286), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n590), .A2(n589), .ZN(G297) );
  NAND2_X1 U664 ( .A1(n608), .A2(G559), .ZN(n591) );
  INV_X1 U665 ( .A(n702), .ZN(n943) );
  NAND2_X1 U666 ( .A1(n591), .A2(n943), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U668 ( .A1(G868), .A2(n944), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G868), .A2(n943), .ZN(n593) );
  NOR2_X1 U670 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U671 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G135), .A2(n870), .ZN(n597) );
  NAND2_X1 U673 ( .A1(G111), .A2(n874), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G123), .A2(n598), .ZN(n599) );
  XNOR2_X1 U676 ( .A(n599), .B(KEYINPUT18), .ZN(n600) );
  XNOR2_X1 U677 ( .A(n600), .B(KEYINPUT77), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n871), .A2(G99), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n914) );
  XNOR2_X1 U681 ( .A(G2096), .B(n914), .ZN(n605) );
  NOR2_X1 U682 ( .A1(G2100), .A2(n605), .ZN(n606) );
  XOR2_X1 U683 ( .A(KEYINPUT78), .B(n606), .Z(G156) );
  NAND2_X1 U684 ( .A1(G559), .A2(n943), .ZN(n607) );
  XOR2_X1 U685 ( .A(n944), .B(n607), .Z(n656) );
  NAND2_X1 U686 ( .A1(n608), .A2(n656), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G55), .A2(n643), .ZN(n609) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT80), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G80), .A2(n634), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G67), .A2(n647), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G93), .A2(n635), .ZN(n612) );
  XNOR2_X1 U693 ( .A(KEYINPUT79), .B(n612), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n659) );
  XNOR2_X1 U696 ( .A(n617), .B(n659), .ZN(G145) );
  NAND2_X1 U697 ( .A1(n643), .A2(G50), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G75), .A2(n634), .ZN(n619) );
  NAND2_X1 U699 ( .A1(G88), .A2(n635), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n647), .A2(G62), .ZN(n620) );
  XOR2_X1 U702 ( .A(KEYINPUT82), .B(n620), .Z(n621) );
  NOR2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U705 ( .A(KEYINPUT83), .B(n625), .Z(G303) );
  INV_X1 U706 ( .A(G303), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G73), .A2(n634), .ZN(n626) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n626), .Z(n631) );
  NAND2_X1 U709 ( .A1(G86), .A2(n635), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G61), .A2(n647), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U712 ( .A(KEYINPUT81), .B(n629), .Z(n630) );
  NOR2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n643), .A2(G48), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U716 ( .A1(G72), .A2(n634), .ZN(n637) );
  NAND2_X1 U717 ( .A1(G85), .A2(n635), .ZN(n636) );
  NAND2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G60), .A2(n647), .ZN(n638) );
  XOR2_X1 U720 ( .A(KEYINPUT66), .B(n638), .Z(n639) );
  NOR2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n643), .A2(G47), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U724 ( .A1(G49), .A2(n643), .ZN(n645) );
  NAND2_X1 U725 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U727 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(G288) );
  XNOR2_X1 U730 ( .A(G166), .B(G305), .ZN(n655) );
  XNOR2_X1 U731 ( .A(G290), .B(G299), .ZN(n653) );
  XOR2_X1 U732 ( .A(KEYINPUT19), .B(G288), .Z(n651) );
  XNOR2_X1 U733 ( .A(n659), .B(n651), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n890) );
  XNOR2_X1 U736 ( .A(n890), .B(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n657), .A2(G868), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(KEYINPUT84), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U740 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n663), .B(KEYINPUT20), .ZN(n664) );
  XNOR2_X1 U743 ( .A(n664), .B(KEYINPUT85), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n668), .B(KEYINPUT22), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(KEYINPUT86), .ZN(n670) );
  NOR2_X1 U751 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G96), .A2(n671), .ZN(n824) );
  NAND2_X1 U753 ( .A1(n824), .A2(G2106), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U755 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U756 ( .A1(G108), .A2(n673), .ZN(n825) );
  NAND2_X1 U757 ( .A1(n825), .A2(G567), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n675), .A2(n674), .ZN(n826) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U760 ( .A1(n826), .A2(n676), .ZN(n823) );
  NAND2_X1 U761 ( .A1(n823), .A2(G36), .ZN(G176) );
  XNOR2_X1 U762 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NAND2_X1 U763 ( .A1(G140), .A2(n870), .ZN(n678) );
  NAND2_X1 U764 ( .A1(G104), .A2(n871), .ZN(n677) );
  NAND2_X1 U765 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U766 ( .A(KEYINPUT34), .B(n679), .ZN(n685) );
  NAND2_X1 U767 ( .A1(n598), .A2(G128), .ZN(n680) );
  XNOR2_X1 U768 ( .A(n680), .B(KEYINPUT88), .ZN(n682) );
  NAND2_X1 U769 ( .A1(G116), .A2(n874), .ZN(n681) );
  NAND2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U771 ( .A(KEYINPUT35), .B(n683), .Z(n684) );
  NOR2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U773 ( .A(KEYINPUT36), .B(n686), .ZN(n885) );
  NOR2_X1 U774 ( .A1(n813), .A2(n885), .ZN(n928) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n688) );
  NOR2_X1 U776 ( .A1(n692), .A2(n688), .ZN(n816) );
  NAND2_X1 U777 ( .A1(n928), .A2(n816), .ZN(n687) );
  XOR2_X1 U778 ( .A(KEYINPUT89), .B(n687), .Z(n811) );
  INV_X1 U779 ( .A(n811), .ZN(n781) );
  INV_X1 U780 ( .A(n688), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n733) );
  NOR2_X1 U782 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NAND2_X1 U783 ( .A1(n756), .A2(KEYINPUT33), .ZN(n690) );
  OR2_X1 U784 ( .A1(n768), .A2(n690), .ZN(n764) );
  AND2_X1 U785 ( .A1(n718), .A2(G1996), .ZN(n693) );
  XOR2_X1 U786 ( .A(n693), .B(KEYINPUT26), .Z(n695) );
  NAND2_X1 U787 ( .A1(n733), .A2(G1341), .ZN(n694) );
  NAND2_X1 U788 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n696), .A2(n944), .ZN(n700) );
  NAND2_X1 U790 ( .A1(G1348), .A2(n733), .ZN(n698) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n718), .ZN(n697) );
  NAND2_X1 U792 ( .A1(n698), .A2(n697), .ZN(n701) );
  NOR2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n699) );
  NOR2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n704) );
  AND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n711) );
  NAND2_X1 U797 ( .A1(G2072), .A2(n718), .ZN(n706) );
  XOR2_X1 U798 ( .A(KEYINPUT98), .B(KEYINPUT27), .Z(n705) );
  XNOR2_X1 U799 ( .A(n706), .B(n705), .ZN(n709) );
  NAND2_X1 U800 ( .A1(G1956), .A2(n733), .ZN(n707) );
  XOR2_X1 U801 ( .A(KEYINPUT99), .B(n707), .Z(n708) );
  NAND2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U803 ( .A1(n713), .A2(G299), .ZN(n710) );
  NOR2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U805 ( .A(KEYINPUT100), .B(n712), .ZN(n716) );
  NAND2_X1 U806 ( .A1(G299), .A2(n713), .ZN(n714) );
  XOR2_X1 U807 ( .A(KEYINPUT28), .B(n714), .Z(n715) );
  NOR2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U809 ( .A(n717), .B(KEYINPUT29), .ZN(n723) );
  XOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .Z(n996) );
  NOR2_X1 U811 ( .A1(n996), .A2(n733), .ZN(n720) );
  NOR2_X1 U812 ( .A1(n718), .A2(G1961), .ZN(n719) );
  NOR2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U814 ( .A(KEYINPUT97), .B(n721), .ZN(n728) );
  NAND2_X1 U815 ( .A1(G171), .A2(n728), .ZN(n722) );
  NAND2_X1 U816 ( .A1(n723), .A2(n722), .ZN(n746) );
  INV_X1 U817 ( .A(n750), .ZN(n725) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n733), .ZN(n748) );
  NAND2_X1 U819 ( .A1(n725), .A2(n517), .ZN(n726) );
  XNOR2_X1 U820 ( .A(n726), .B(KEYINPUT30), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n727), .A2(G168), .ZN(n730) );
  NOR2_X1 U822 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n732) );
  INV_X1 U824 ( .A(KEYINPUT31), .ZN(n731) );
  XNOR2_X1 U825 ( .A(n732), .B(n731), .ZN(n747) );
  NOR2_X1 U826 ( .A1(G1971), .A2(n768), .ZN(n735) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U830 ( .A1(n724), .A2(n737), .ZN(n739) );
  AND2_X1 U831 ( .A1(n747), .A2(n739), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n746), .A2(n738), .ZN(n743) );
  INV_X1 U833 ( .A(n739), .ZN(n741) );
  AND2_X1 U834 ( .A1(G286), .A2(G8), .ZN(n740) );
  OR2_X1 U835 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U836 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n752) );
  AND2_X1 U838 ( .A1(G8), .A2(n748), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n952) );
  NAND2_X1 U843 ( .A1(n770), .A2(n952), .ZN(n759) );
  NAND2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n948) );
  INV_X1 U845 ( .A(n948), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n757), .A2(n768), .ZN(n758) );
  NOR2_X1 U847 ( .A1(KEYINPUT33), .A2(n760), .ZN(n762) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n958) );
  INV_X1 U849 ( .A(n958), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n765), .B(KEYINPUT102), .ZN(n779) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XNOR2_X1 U853 ( .A(n766), .B(KEYINPUT24), .ZN(n767) );
  XNOR2_X1 U854 ( .A(n767), .B(KEYINPUT96), .ZN(n769) );
  INV_X1 U855 ( .A(n768), .ZN(n775) );
  AND2_X1 U856 ( .A1(n769), .A2(n775), .ZN(n777) );
  INV_X1 U857 ( .A(n770), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G166), .A2(G8), .ZN(n771) );
  NOR2_X1 U859 ( .A1(G2090), .A2(n771), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n781), .A2(n780), .ZN(n804) );
  NAND2_X1 U864 ( .A1(G141), .A2(n870), .ZN(n783) );
  NAND2_X1 U865 ( .A1(G117), .A2(n874), .ZN(n782) );
  NAND2_X1 U866 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U867 ( .A1(n871), .A2(G105), .ZN(n784) );
  XOR2_X1 U868 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U869 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U870 ( .A1(n598), .A2(G129), .ZN(n787) );
  NAND2_X1 U871 ( .A1(n788), .A2(n787), .ZN(n863) );
  NAND2_X1 U872 ( .A1(G1996), .A2(n863), .ZN(n789) );
  XOR2_X1 U873 ( .A(KEYINPUT93), .B(n789), .Z(n799) );
  XNOR2_X1 U874 ( .A(KEYINPUT92), .B(G1991), .ZN(n1000) );
  NAND2_X1 U875 ( .A1(G131), .A2(n870), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G95), .A2(n871), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(KEYINPUT91), .B(n792), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G119), .A2(n598), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G107), .A2(n874), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U882 ( .A(KEYINPUT90), .B(n795), .Z(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n864) );
  NAND2_X1 U884 ( .A1(n1000), .A2(n864), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n920) );
  NAND2_X1 U886 ( .A1(n920), .A2(n816), .ZN(n800) );
  XOR2_X1 U887 ( .A(KEYINPUT94), .B(n800), .Z(n808) );
  XNOR2_X1 U888 ( .A(G1986), .B(G290), .ZN(n954) );
  NAND2_X1 U889 ( .A1(n816), .A2(n954), .ZN(n801) );
  XNOR2_X1 U890 ( .A(KEYINPUT87), .B(n801), .ZN(n802) );
  NOR2_X1 U891 ( .A1(n808), .A2(n802), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n818) );
  NOR2_X1 U893 ( .A1(G1996), .A2(n863), .ZN(n923) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U895 ( .A1(n1000), .A2(n864), .ZN(n916) );
  NOR2_X1 U896 ( .A1(n805), .A2(n916), .ZN(n806) );
  XOR2_X1 U897 ( .A(KEYINPUT103), .B(n806), .Z(n807) );
  NOR2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U899 ( .A1(n923), .A2(n809), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U902 ( .A1(n813), .A2(n885), .ZN(n930) );
  NAND2_X1 U903 ( .A1(n814), .A2(n930), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U905 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U906 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U909 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U911 ( .A1(n823), .A2(n822), .ZN(G188) );
  INV_X1 U913 ( .A(G132), .ZN(G219) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G82), .ZN(G220) );
  INV_X1 U916 ( .A(G69), .ZN(G235) );
  NOR2_X1 U917 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U918 ( .A(G325), .ZN(G261) );
  INV_X1 U919 ( .A(n826), .ZN(G319) );
  XNOR2_X1 U920 ( .A(G1996), .B(G2474), .ZN(n836) );
  XOR2_X1 U921 ( .A(G1981), .B(G1961), .Z(n828) );
  XNOR2_X1 U922 ( .A(G1991), .B(G1966), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U924 ( .A(G1976), .B(G1971), .Z(n830) );
  XNOR2_X1 U925 ( .A(G1986), .B(G1956), .ZN(n829) );
  XNOR2_X1 U926 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U927 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U928 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U930 ( .A(n836), .B(n835), .ZN(G229) );
  XOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .Z(n838) );
  XNOR2_X1 U932 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n837) );
  XNOR2_X1 U933 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U934 ( .A(KEYINPUT43), .B(G2090), .Z(n840) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U937 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U938 ( .A(G2096), .B(G2100), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n844), .B(n843), .ZN(n846) );
  XOR2_X1 U940 ( .A(G2078), .B(G2084), .Z(n845) );
  XNOR2_X1 U941 ( .A(n846), .B(n845), .ZN(G227) );
  NAND2_X1 U942 ( .A1(G100), .A2(n871), .ZN(n853) );
  NAND2_X1 U943 ( .A1(G136), .A2(n870), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G112), .A2(n874), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n851) );
  NAND2_X1 U946 ( .A1(n598), .A2(G124), .ZN(n849) );
  XOR2_X1 U947 ( .A(KEYINPUT44), .B(n849), .Z(n850) );
  NOR2_X1 U948 ( .A1(n851), .A2(n850), .ZN(n852) );
  NAND2_X1 U949 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n854), .B(KEYINPUT111), .ZN(G162) );
  NAND2_X1 U951 ( .A1(G130), .A2(n598), .ZN(n856) );
  NAND2_X1 U952 ( .A1(G118), .A2(n874), .ZN(n855) );
  NAND2_X1 U953 ( .A1(n856), .A2(n855), .ZN(n861) );
  NAND2_X1 U954 ( .A1(G142), .A2(n870), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G106), .A2(n871), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n859), .B(KEYINPUT45), .Z(n860) );
  NOR2_X1 U958 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n862), .B(n914), .ZN(n884) );
  XNOR2_X1 U960 ( .A(G160), .B(n863), .ZN(n865) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U962 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U965 ( .A(n869), .B(n868), .Z(n882) );
  NAND2_X1 U966 ( .A1(G139), .A2(n870), .ZN(n873) );
  NAND2_X1 U967 ( .A1(G103), .A2(n871), .ZN(n872) );
  NAND2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n880) );
  NAND2_X1 U969 ( .A1(G127), .A2(n598), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G115), .A2(n874), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U972 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  XNOR2_X1 U973 ( .A(KEYINPUT112), .B(n878), .ZN(n879) );
  NOR2_X1 U974 ( .A1(n880), .A2(n879), .ZN(n932) );
  XNOR2_X1 U975 ( .A(G164), .B(n932), .ZN(n881) );
  XNOR2_X1 U976 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U977 ( .A(n884), .B(n883), .ZN(n887) );
  XNOR2_X1 U978 ( .A(n885), .B(G162), .ZN(n886) );
  XNOR2_X1 U979 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U980 ( .A1(G37), .A2(n888), .ZN(n889) );
  XOR2_X1 U981 ( .A(KEYINPUT115), .B(n889), .Z(G395) );
  XNOR2_X1 U982 ( .A(n943), .B(G286), .ZN(n891) );
  XNOR2_X1 U983 ( .A(n891), .B(n890), .ZN(n893) );
  XNOR2_X1 U984 ( .A(n944), .B(G171), .ZN(n892) );
  XNOR2_X1 U985 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U986 ( .A1(G37), .A2(n894), .ZN(G397) );
  XOR2_X1 U987 ( .A(G2427), .B(KEYINPUT107), .Z(n896) );
  XNOR2_X1 U988 ( .A(G1341), .B(G1348), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n906) );
  XOR2_X1 U990 ( .A(G2451), .B(G2435), .Z(n898) );
  XNOR2_X1 U991 ( .A(G2430), .B(G2438), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U993 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n900) );
  XNOR2_X1 U994 ( .A(G2443), .B(G2454), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U996 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U997 ( .A(G2446), .B(KEYINPUT104), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n906), .B(n905), .ZN(n907) );
  NAND2_X1 U1000 ( .A1(n907), .A2(G14), .ZN(n913) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n913), .ZN(n910) );
  NOR2_X1 U1002 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n911) );
  NAND2_X1 U1006 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G96), .ZN(G221) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(n913), .ZN(G401) );
  XNOR2_X1 U1011 ( .A(G160), .B(G2084), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1014 ( .A(KEYINPUT116), .B(n918), .Z(n919) );
  NOR2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n926) );
  XNOR2_X1 U1016 ( .A(G2090), .B(G162), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n921), .B(KEYINPUT117), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n924), .Z(n925) );
  NAND2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(n929), .B(KEYINPUT118), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(n931), .A2(n930), .ZN(n938) );
  XOR2_X1 U1024 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n936) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n934) );
  XOR2_X1 U1026 ( .A(G2072), .B(n932), .Z(n933) );
  NOR2_X1 U1027 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1028 ( .A(n936), .B(n935), .Z(n937) );
  NOR2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n939), .ZN(n941) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1032 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1033 ( .A1(n942), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1034 ( .A(G16), .B(KEYINPUT56), .ZN(n967) );
  XNOR2_X1 U1035 ( .A(n943), .B(G1348), .ZN(n965) );
  XOR2_X1 U1036 ( .A(G171), .B(G1961), .Z(n946) );
  XNOR2_X1 U1037 ( .A(n944), .B(G1341), .ZN(n945) );
  NOR2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n957) );
  XOR2_X1 U1039 ( .A(G1956), .B(G299), .Z(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n950) );
  AND2_X1 U1041 ( .A1(G303), .A2(G1971), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1043 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1044 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(n955), .B(KEYINPUT124), .ZN(n956) );
  NAND2_X1 U1046 ( .A1(n957), .A2(n956), .ZN(n963) );
  XNOR2_X1 U1047 ( .A(G1966), .B(G168), .ZN(n959) );
  NAND2_X1 U1048 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1049 ( .A(KEYINPUT57), .B(n960), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(KEYINPUT123), .B(n961), .ZN(n962) );
  NOR2_X1 U1051 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1052 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1053 ( .A1(n967), .A2(n966), .ZN(n994) );
  INV_X1 U1054 ( .A(G16), .ZN(n992) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G21), .ZN(n969) );
  XNOR2_X1 U1056 ( .A(G1961), .B(G5), .ZN(n968) );
  NOR2_X1 U1057 ( .A1(n969), .A2(n968), .ZN(n979) );
  XOR2_X1 U1058 ( .A(G1348), .B(KEYINPUT59), .Z(n970) );
  XNOR2_X1 U1059 ( .A(G4), .B(n970), .ZN(n972) );
  XNOR2_X1 U1060 ( .A(G20), .B(G1956), .ZN(n971) );
  NOR2_X1 U1061 ( .A1(n972), .A2(n971), .ZN(n976) );
  XNOR2_X1 U1062 ( .A(G1341), .B(G19), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G6), .B(G1981), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1066 ( .A(KEYINPUT60), .B(n977), .Z(n978) );
  NAND2_X1 U1067 ( .A1(n979), .A2(n978), .ZN(n989) );
  XNOR2_X1 U1068 ( .A(KEYINPUT125), .B(G1976), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(n980), .B(G23), .ZN(n985) );
  XNOR2_X1 U1070 ( .A(G1986), .B(KEYINPUT126), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n981), .B(G24), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G22), .B(G1971), .ZN(n982) );
  NOR2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1075 ( .A(KEYINPUT127), .B(n986), .Z(n987) );
  XNOR2_X1 U1076 ( .A(KEYINPUT58), .B(n987), .ZN(n988) );
  NOR2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1078 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NAND2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1080 ( .A1(n994), .A2(n993), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(G2072), .B(G33), .Z(n995) );
  NAND2_X1 U1082 ( .A1(G28), .A2(n995), .ZN(n1006) );
  XNOR2_X1 U1083 ( .A(G1996), .B(G32), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(n996), .B(G27), .ZN(n997) );
  NOR2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(KEYINPUT120), .B(n999), .ZN(n1004) );
  XNOR2_X1 U1087 ( .A(n1000), .B(G25), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(G2067), .B(G26), .ZN(n1001) );
  NOR2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1091 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1092 ( .A(KEYINPUT53), .B(n1007), .Z(n1011) );
  XNOR2_X1 U1093 ( .A(KEYINPUT54), .B(G34), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(n1008), .B(KEYINPUT121), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G2084), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1097 ( .A(G35), .B(G2090), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1014), .B(KEYINPUT55), .ZN(n1016) );
  INV_X1 U1100 ( .A(G29), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT122), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

