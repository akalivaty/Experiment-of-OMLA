//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1194, new_n1195,
    new_n1196, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1247, new_n1248, new_n1249, new_n1250;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g0006(.A(KEYINPUT64), .B(G238), .Z(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT65), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n220), .A2(new_n204), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n206), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NOR4_X1   g0025(.A1(new_n218), .A2(new_n219), .A3(new_n222), .A4(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G250), .B(G257), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT66), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n230), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT67), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n208), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n208), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n204), .A2(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n221), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n246), .A2(new_n255), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n203), .A2(G20), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G68), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n248), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(KEYINPUT11), .B1(new_n253), .B2(new_n255), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G97), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n276), .A2(new_n232), .A3(new_n269), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n266), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n279));
  AND2_X1   g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  OAI21_X1  g0080(.A(G274), .B1(new_n280), .B2(new_n221), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n265), .A2(new_n282), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(new_n285), .B2(G238), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n278), .A2(new_n279), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n278), .A2(new_n286), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT13), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n289), .B2(KEYINPUT71), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n287), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n279), .B1(new_n278), .B2(new_n286), .ZN(new_n294));
  OAI21_X1  g0094(.A(G169), .B1(new_n287), .B2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n293), .A2(G179), .B1(KEYINPUT14), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT72), .B(KEYINPUT14), .ZN(new_n297));
  OAI211_X1 g0097(.A(G169), .B(new_n297), .C1(new_n287), .C2(new_n294), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT73), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n262), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n293), .A2(G190), .ZN(new_n302));
  OAI21_X1  g0102(.A(G200), .B1(new_n287), .B2(new_n294), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(new_n262), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(KEYINPUT8), .B(G58), .ZN(new_n306));
  INV_X1    g0106(.A(G150), .ZN(new_n307));
  INV_X1    g0107(.A(new_n249), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n306), .A2(new_n252), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(G50), .A2(G58), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n204), .B1(new_n310), .B2(new_n208), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n255), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G50), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n203), .B2(G20), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n257), .A2(new_n314), .B1(new_n313), .B2(new_n246), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n268), .A2(G1698), .ZN(new_n318));
  INV_X1    g0118(.A(G223), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n317), .B1(new_n251), .B2(new_n268), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n266), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n283), .B1(new_n285), .B2(G226), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n316), .B1(new_n324), .B2(G169), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(G179), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(G200), .B2(new_n323), .ZN(new_n330));
  XNOR2_X1  g0130(.A(new_n316), .B(KEYINPUT69), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT9), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n331), .A2(new_n332), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n330), .B(new_n337), .C1(new_n333), .C2(new_n334), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n327), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n306), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n341), .B1(new_n252), .B2(new_n342), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n343), .A2(new_n255), .B1(new_n251), .B2(new_n246), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n257), .A2(G77), .A3(new_n258), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n285), .A2(G244), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n349));
  INV_X1    g0149(.A(G107), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n349), .B1(new_n350), .B2(new_n268), .C1(new_n318), .C2(new_n207), .ZN(new_n351));
  AOI211_X1 g0151(.A(new_n283), .B(new_n348), .C1(new_n351), .C2(new_n266), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(G190), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n353), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n347), .B1(new_n352), .B2(G169), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n339), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT16), .ZN(new_n363));
  INV_X1    g0163(.A(G58), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n208), .ZN(new_n365));
  NOR2_X1   g0165(.A1(G58), .A2(G68), .ZN(new_n366));
  OAI21_X1  g0166(.A(G20), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n249), .A2(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n268), .B2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n208), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AOI211_X1 g0176(.A(KEYINPUT74), .B(new_n208), .C1(new_n372), .C2(new_n373), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n363), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n255), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n374), .A2(new_n369), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n306), .B1(new_n203), .B2(G20), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n257), .B1(new_n246), .B2(new_n306), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n273), .A2(new_n275), .A3(G223), .A4(new_n269), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n273), .A2(new_n275), .A3(G226), .A4(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT75), .A4(new_n387), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n265), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT76), .B1(new_n284), .B2(new_n232), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT76), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n265), .A2(new_n395), .A3(G232), .A4(new_n282), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n283), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(G190), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n396), .ZN(new_n399));
  INV_X1    g0199(.A(new_n283), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(G200), .B1(new_n392), .B2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n382), .A2(new_n384), .A3(new_n398), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n398), .A2(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(new_n384), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n378), .B2(new_n381), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT17), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n362), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n382), .A2(new_n384), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n393), .A2(G179), .A3(new_n397), .ZN(new_n413));
  OAI21_X1  g0213(.A(G169), .B1(new_n392), .B2(new_n401), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n411), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n412), .B1(new_n411), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n403), .A2(new_n404), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n406), .A2(KEYINPUT17), .A3(new_n408), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT77), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n410), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n305), .A2(new_n361), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n203), .A2(G33), .ZN(new_n424));
  AND4_X1   g0224(.A1(new_n221), .A2(new_n245), .A3(new_n254), .A4(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n350), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT25), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n245), .B2(G107), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n425), .A2(G107), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT86), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n273), .A2(new_n275), .A3(new_n204), .A4(G87), .ZN(new_n431));
  AND2_X1   g0231(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n432));
  NOR2_X1   g0232(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n268), .A2(new_n204), .A3(G87), .A4(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G116), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n437), .A2(G20), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT23), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n204), .B2(G107), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n350), .A2(KEYINPUT23), .A3(G20), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n435), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT24), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT24), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n435), .A2(new_n436), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n430), .B1(new_n447), .B2(new_n255), .ZN(new_n448));
  AOI211_X1 g0248(.A(KEYINPUT86), .B(new_n379), .C1(new_n444), .C2(new_n446), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n429), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT87), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(KEYINPUT87), .B(new_n429), .C1(new_n448), .C2(new_n449), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT5), .B(G41), .ZN(new_n454));
  INV_X1    g0254(.A(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(G1), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n454), .A2(new_n265), .A3(G274), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(new_n456), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n265), .ZN(new_n459));
  INV_X1    g0259(.A(G264), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n462));
  INV_X1    g0262(.A(G294), .ZN(new_n463));
  INV_X1    g0263(.A(G250), .ZN(new_n464));
  OAI221_X1 g0264(.A(new_n462), .B1(new_n263), .B2(new_n463), .C1(new_n270), .C2(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n461), .B1(new_n465), .B2(new_n266), .ZN(new_n466));
  INV_X1    g0266(.A(G169), .ZN(new_n467));
  OR3_X1    g0267(.A1(new_n466), .A2(KEYINPUT88), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n466), .A2(G179), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT88), .B1(new_n466), .B2(new_n467), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n452), .A2(new_n453), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT89), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT89), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n452), .A2(new_n471), .A3(new_n474), .A4(new_n453), .ZN(new_n475));
  INV_X1    g0275(.A(new_n450), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n466), .A2(G190), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n477), .C1(new_n354), .C2(new_n466), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  INV_X1    g0281(.A(G116), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n254), .A2(new_n221), .B1(G20), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n204), .C1(G33), .C2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT20), .B1(new_n483), .B2(new_n486), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n245), .A2(G116), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n379), .A2(new_n245), .A3(new_n424), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n492), .B2(new_n482), .ZN(new_n493));
  OAI21_X1  g0293(.A(G169), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n273), .A2(new_n275), .A3(G257), .A4(new_n269), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n273), .A2(new_n275), .A3(G264), .A4(G1698), .ZN(new_n496));
  XOR2_X1   g0296(.A(KEYINPUT81), .B(G303), .Z(new_n497));
  OAI211_X1 g0297(.A(new_n495), .B(new_n496), .C1(new_n497), .C2(new_n268), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n498), .A2(KEYINPUT82), .A3(new_n266), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT82), .B1(new_n498), .B2(new_n266), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n458), .A2(G270), .A3(new_n265), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n457), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n502), .A2(KEYINPUT80), .A3(new_n457), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n494), .B1(new_n501), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT83), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n481), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n498), .A2(new_n266), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT82), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n498), .A2(KEYINPUT82), .A3(new_n266), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n502), .A2(KEYINPUT80), .A3(new_n457), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT80), .B1(new_n502), .B2(new_n457), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n494), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n517), .A2(new_n509), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT84), .B1(new_n510), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n517), .A2(new_n518), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT21), .B1(new_n521), .B2(KEYINPUT83), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT84), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n508), .A2(new_n509), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n489), .ZN(new_n527));
  INV_X1    g0327(.A(new_n493), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n356), .ZN(new_n531));
  INV_X1    g0331(.A(new_n517), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n481), .B2(new_n521), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n529), .B1(new_n517), .B2(G200), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n328), .B2(new_n517), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n246), .A2(new_n485), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n492), .B2(new_n485), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n308), .A2(new_n251), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  AND2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n350), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n540), .B1(new_n546), .B2(G20), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT78), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n372), .A2(new_n373), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G107), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT78), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n204), .B1(new_n544), .B2(new_n545), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n540), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n539), .B1(new_n554), .B2(new_n255), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n273), .A2(new_n275), .A3(G250), .A4(G1698), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(new_n269), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT4), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n484), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n266), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n266), .B1(new_n456), .B2(new_n454), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G257), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n457), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G200), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n555), .B(new_n565), .C1(new_n328), .C2(new_n564), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n467), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n557), .A2(new_n558), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(new_n484), .A4(new_n556), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n266), .B1(G257), .B2(new_n562), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n356), .A3(new_n457), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n547), .A2(KEYINPUT78), .B1(new_n549), .B2(G107), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n379), .B1(new_n573), .B2(new_n553), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n567), .B(new_n572), .C1(new_n574), .C2(new_n539), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n273), .A2(new_n275), .A3(G238), .A4(new_n269), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n437), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n266), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n265), .A2(G274), .A3(new_n456), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT79), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n456), .A2(new_n464), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n581), .A2(new_n582), .B1(new_n265), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n265), .A2(KEYINPUT79), .A3(G274), .A4(new_n456), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n584), .A3(G190), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n204), .B1(new_n267), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n543), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n273), .A2(new_n275), .A3(new_n204), .A4(G68), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n587), .B1(new_n252), .B2(new_n485), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(new_n255), .B1(new_n246), .B2(new_n342), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n425), .A2(G87), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n586), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n456), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n582), .B1(new_n281), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n583), .A2(new_n265), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n599), .A2(new_n585), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n354), .B1(new_n601), .B2(new_n580), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n580), .A2(new_n584), .A3(new_n356), .A4(new_n585), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n594), .A2(new_n255), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n342), .A2(new_n246), .ZN(new_n605));
  INV_X1    g0405(.A(new_n342), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n425), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(G169), .B1(new_n601), .B2(new_n580), .ZN(new_n610));
  OAI22_X1  g0410(.A1(new_n597), .A2(new_n602), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n576), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n526), .A2(new_n535), .A3(new_n537), .A4(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n423), .A2(new_n480), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g0415(.A(new_n615), .B(KEYINPUT90), .Z(G372));
  AOI21_X1  g0416(.A(new_n300), .B1(new_n304), .B2(new_n359), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n410), .A2(new_n421), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n418), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n336), .A2(new_n338), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n327), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n423), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n534), .B1(new_n520), .B2(new_n525), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n471), .A2(new_n450), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n576), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n584), .A2(new_n585), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT91), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n580), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n579), .A2(KEYINPUT91), .A3(new_n266), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT92), .B1(new_n631), .B2(new_n354), .ZN(new_n632));
  INV_X1    g0432(.A(new_n630), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT91), .B1(new_n579), .B2(new_n266), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n601), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT92), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(G200), .ZN(new_n637));
  INV_X1    g0437(.A(new_n597), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n632), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n603), .B(new_n608), .C1(new_n631), .C2(G169), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n478), .A2(new_n626), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n625), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  INV_X1    g0444(.A(new_n575), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT26), .B1(new_n575), .B2(new_n611), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n646), .A2(new_n640), .A3(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n643), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n621), .B1(new_n622), .B2(new_n649), .ZN(new_n650));
  XOR2_X1   g0450(.A(new_n650), .B(KEYINPUT93), .Z(G369));
  NAND2_X1  g0451(.A1(new_n526), .A2(new_n535), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n530), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n623), .A2(new_n537), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n660), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n452), .A2(new_n453), .A3(new_n658), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n479), .A2(new_n666), .B1(new_n472), .B2(new_n659), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n652), .A2(new_n659), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n479), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n624), .A2(new_n658), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(G399));
  INV_X1    g0473(.A(new_n223), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n590), .A2(G116), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G1), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n220), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n623), .A2(new_n473), .A3(new_n475), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n642), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n644), .B1(new_n575), .B2(new_n611), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT94), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n645), .A2(new_n639), .A3(KEYINPUT26), .A4(new_n640), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT94), .B(new_n644), .C1(new_n575), .C2(new_n611), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n640), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT95), .B1(new_n691), .B2(new_n659), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT95), .ZN(new_n693));
  AOI211_X1 g0493(.A(new_n693), .B(new_n658), .C1(new_n682), .C2(new_n690), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT29), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n658), .B1(new_n643), .B2(new_n648), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(KEYINPUT29), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n480), .A2(new_n614), .A3(new_n659), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n601), .A2(new_n580), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n466), .A2(new_n701), .A3(G179), .A4(new_n571), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  OR3_X1    g0503(.A1(new_n702), .A2(new_n703), .A3(new_n517), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n466), .A2(G179), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n517), .A3(new_n564), .A4(new_n635), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n702), .B2(new_n517), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n708), .A2(new_n709), .A3(new_n658), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n709), .B1(new_n708), .B2(new_n658), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n700), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n699), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n680), .B1(new_n718), .B2(G1), .ZN(G364));
  AND2_X1   g0519(.A1(new_n204), .A2(G13), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n203), .B1(new_n720), .B2(G45), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n675), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n665), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(G330), .B2(new_n663), .ZN(new_n725));
  INV_X1    g0525(.A(new_n723), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n221), .B1(G20), .B2(new_n467), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n204), .A2(new_n356), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(G190), .A3(new_n354), .ZN(new_n730));
  INV_X1    g0530(.A(G322), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n204), .A2(G179), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G190), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G329), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n730), .A2(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G283), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n732), .A2(new_n328), .A3(G200), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n732), .A2(G190), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(G303), .ZN(new_n740));
  OAI22_X1  g0540(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n328), .A2(G179), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n204), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n463), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n729), .A2(new_n733), .ZN(new_n745));
  INV_X1    g0545(.A(G311), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n276), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR4_X1   g0547(.A1(new_n736), .A2(new_n741), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n729), .A2(G200), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT98), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n328), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G326), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n751), .A2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  XOR2_X1   g0556(.A(KEYINPUT33), .B(G317), .Z(new_n757));
  OAI221_X1 g0557(.A(new_n748), .B1(new_n753), .B2(new_n754), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(G50), .A2(new_n752), .B1(new_n755), .B2(G68), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n738), .A2(new_n350), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n743), .A2(new_n485), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT32), .ZN(new_n762));
  INV_X1    g0562(.A(new_n734), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(G159), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n760), .B(new_n761), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n268), .B1(new_n730), .B2(new_n364), .ZN(new_n766));
  INV_X1    g0566(.A(new_n745), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(G77), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n764), .ZN(new_n769));
  INV_X1    g0569(.A(new_n739), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n769), .A2(KEYINPUT32), .B1(new_n770), .B2(G87), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n759), .A2(new_n765), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n728), .B1(new_n758), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT97), .Z(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n727), .ZN(new_n777));
  INV_X1    g0577(.A(new_n220), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n455), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n674), .A2(new_n268), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n240), .C2(new_n455), .ZN(new_n781));
  INV_X1    g0581(.A(G355), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(KEYINPUT96), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n223), .A2(new_n268), .A3(new_n784), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n781), .B1(G116), .B2(new_n223), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n726), .B(new_n773), .C1(new_n777), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n776), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n663), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n725), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(G396));
  AOI22_X1  g0591(.A1(G283), .A2(new_n755), .B1(new_n752), .B2(G303), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n730), .A2(new_n463), .B1(new_n745), .B2(new_n482), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n268), .B(new_n793), .C1(G311), .C2(new_n763), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n738), .A2(new_n589), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n795), .B(new_n761), .C1(G107), .C2(new_n770), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n792), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n730), .ZN(new_n798));
  XOR2_X1   g0598(.A(KEYINPUT99), .B(G143), .Z(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n798), .A2(new_n800), .B1(new_n767), .B2(G159), .ZN(new_n801));
  INV_X1    g0601(.A(G137), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n801), .B1(new_n753), .B2(new_n802), .C1(new_n307), .C2(new_n756), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT100), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n268), .B1(new_n734), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT101), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n743), .A2(new_n364), .B1(new_n739), .B2(new_n313), .ZN(new_n809));
  INV_X1    g0609(.A(new_n738), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G68), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n805), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n797), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n727), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n727), .A2(new_n774), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n815), .B1(G77), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n359), .A2(new_n659), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n347), .A2(new_n658), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n355), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n820), .B1(new_n360), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n775), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n723), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n717), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n696), .B(new_n823), .Z(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n726), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n825), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT102), .ZN(G384));
  OR2_X1    g0632(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n221), .A2(new_n204), .A3(new_n482), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT36), .Z(new_n837));
  OAI211_X1 g0637(.A(new_n778), .B(G77), .C1(new_n364), .C2(new_n208), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n313), .A2(G68), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n203), .B(G13), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n374), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(KEYINPUT16), .A3(new_n370), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n363), .B1(new_n374), .B2(new_n369), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(new_n255), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n384), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n415), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n403), .A3(KEYINPUT103), .ZN(new_n848));
  INV_X1    g0648(.A(new_n656), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT103), .B1(new_n847), .B2(new_n403), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n411), .A2(new_n415), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n656), .B(KEYINPUT104), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n411), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .A4(new_n403), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT105), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n859), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n853), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n850), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n422), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n862), .A2(new_n864), .A3(KEYINPUT38), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT40), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n262), .A2(new_n659), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n301), .A2(new_n304), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n304), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n870), .B1(new_n300), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n869), .A2(new_n714), .A3(new_n823), .A4(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n854), .A2(new_n403), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n877), .A2(KEYINPUT105), .A3(new_n857), .A4(new_n856), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n858), .A2(new_n859), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n854), .A2(new_n856), .A3(new_n403), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n878), .A2(new_n879), .B1(KEYINPUT37), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n405), .A2(new_n409), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n856), .B1(new_n882), .B2(new_n418), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n866), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n868), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n885), .A2(new_n714), .A3(new_n823), .A4(new_n875), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(KEYINPUT40), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n716), .B1(new_n876), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n423), .B2(new_n717), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT106), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n876), .A2(new_n887), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n622), .A2(new_n715), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT39), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n885), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n867), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n300), .A2(new_n659), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n418), .A2(new_n855), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n820), .B1(new_n696), .B2(new_n823), .ZN(new_n901));
  INV_X1    g0701(.A(new_n875), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n867), .A2(new_n868), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n695), .A2(new_n423), .A3(new_n698), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n907), .A2(new_n621), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n906), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n893), .A2(new_n909), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT107), .ZN(new_n912));
  OAI221_X1 g0712(.A(new_n910), .B1(new_n203), .B2(new_n720), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n911), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(KEYINPUT107), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n841), .B1(new_n913), .B2(new_n915), .ZN(G367));
  OAI21_X1  g0716(.A(new_n626), .B1(new_n555), .B2(new_n659), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n575), .B2(new_n659), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n670), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT42), .Z(new_n920));
  AOI21_X1  g0720(.A(new_n917), .B1(new_n473), .B2(new_n475), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n659), .B1(new_n921), .B2(new_n645), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n595), .A2(new_n596), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n658), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n641), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n640), .B2(new_n925), .ZN(new_n927));
  OR3_X1    g0727(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT108), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n927), .B(KEYINPUT43), .Z(new_n931));
  AOI22_X1  g0731(.A1(new_n928), .A2(new_n929), .B1(new_n923), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT109), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n668), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n918), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n933), .B1(new_n930), .B2(new_n932), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n935), .B2(new_n938), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n675), .B(KEYINPUT41), .Z(new_n941));
  NOR2_X1   g0741(.A1(new_n672), .A2(new_n918), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT110), .Z(new_n943));
  INV_X1    g0743(.A(KEYINPUT44), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n672), .A2(new_n918), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT45), .Z(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(new_n936), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n936), .ZN(new_n951));
  MUX2_X1   g0751(.A(new_n479), .B(new_n667), .S(new_n669), .Z(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n664), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n718), .A2(new_n953), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n941), .B1(new_n955), .B2(new_n718), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n939), .B(new_n940), .C1(new_n956), .C2(new_n722), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n777), .B1(new_n223), .B2(new_n342), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n780), .A2(new_n229), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n723), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G159), .A2(new_n755), .B1(new_n752), .B2(new_n800), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n745), .A2(new_n313), .B1(new_n734), .B2(new_n802), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n276), .B(new_n962), .C1(G150), .C2(new_n798), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n739), .A2(new_n364), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n738), .A2(new_n251), .ZN(new_n965));
  INV_X1    g0765(.A(new_n743), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n964), .B(new_n965), .C1(G68), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n961), .A2(new_n963), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n770), .A2(G116), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT46), .ZN(new_n970));
  INV_X1    g0770(.A(new_n497), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n268), .B1(new_n798), .B2(new_n971), .ZN(new_n972));
  AOI22_X1  g0772(.A1(G283), .A2(new_n767), .B1(new_n763), .B2(G317), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n966), .A2(G107), .B1(new_n810), .B2(G97), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n463), .A2(new_n756), .B1(new_n753), .B2(new_n746), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n968), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT111), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n960), .B1(new_n979), .B2(new_n727), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n788), .B2(new_n927), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n957), .A2(new_n981), .ZN(G387));
  NAND2_X1  g0782(.A1(new_n340), .A2(new_n313), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT50), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n677), .B(new_n455), .C1(new_n208), .C2(new_n251), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n780), .B1(new_n984), .B2(new_n985), .C1(new_n235), .C2(new_n455), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n674), .A2(new_n677), .A3(new_n276), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n350), .B2(new_n674), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n986), .A2(KEYINPUT112), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n777), .ZN(new_n990));
  AOI21_X1  g0790(.A(KEYINPUT112), .B1(new_n986), .B2(new_n988), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n723), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n743), .A2(new_n342), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n268), .B1(new_n745), .B2(new_n208), .C1(new_n313), .C2(new_n730), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(G97), .C2(new_n810), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n755), .A2(new_n340), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n739), .A2(new_n251), .B1(new_n734), .B2(new_n307), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT113), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n752), .A2(G159), .B1(KEYINPUT113), .B2(new_n997), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n966), .A2(G283), .B1(new_n770), .B2(G294), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G317), .A2(new_n798), .B1(new_n971), .B2(new_n767), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n753), .B2(new_n731), .C1(new_n746), .C2(new_n756), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n1005), .B(KEYINPUT114), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT49), .Z(new_n1009));
  OAI221_X1 g0809(.A(new_n276), .B1(new_n734), .B2(new_n754), .C1(new_n482), .C2(new_n738), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n992), .B1(new_n1011), .B2(new_n727), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n667), .A2(new_n788), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n1012), .A2(new_n1013), .B1(new_n953), .B2(new_n722), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n718), .A2(new_n953), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1016), .A2(new_n675), .A3(new_n954), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1015), .A2(KEYINPUT115), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(G393));
  OAI21_X1  g0819(.A(new_n954), .B1(new_n950), .B2(new_n951), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n955), .A2(new_n675), .A3(new_n1020), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n950), .A2(new_n951), .A3(new_n721), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n777), .B1(new_n485), .B2(new_n223), .ZN(new_n1023));
  NOR3_X1   g0823(.A1(new_n243), .A2(new_n674), .A3(new_n268), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n723), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n752), .A2(G317), .B1(G311), .B2(new_n798), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT52), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n756), .A2(new_n497), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n276), .B1(new_n734), .B2(new_n731), .C1(new_n463), .C2(new_n745), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n760), .B1(G283), .B2(new_n770), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n482), .B2(new_n743), .ZN(new_n1031));
  NOR4_X1   g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(KEYINPUT116), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n752), .A2(G150), .B1(G159), .B2(new_n798), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT51), .Z(new_n1036));
  OAI221_X1 g0836(.A(new_n268), .B1(new_n745), .B2(new_n306), .C1(new_n734), .C2(new_n799), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n795), .B1(G68), .B2(new_n770), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n251), .B2(new_n743), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(G50), .C2(new_n755), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1033), .A2(new_n1034), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1025), .B1(new_n1042), .B2(new_n727), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n788), .B2(new_n918), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1021), .A2(new_n1022), .A3(new_n1044), .ZN(G390));
  NAND3_X1  g0845(.A1(new_n691), .A2(KEYINPUT95), .A3(new_n659), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n689), .B1(new_n642), .B2(new_n681), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n693), .B1(new_n1047), .B2(new_n658), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1048), .A3(new_n819), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n822), .A2(new_n360), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n875), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n885), .A2(new_n898), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n897), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n714), .A2(G330), .A3(new_n823), .A4(new_n875), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1053), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n717), .A2(new_n423), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n907), .A2(new_n621), .A3(new_n1062), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n479), .A2(new_n613), .A3(new_n658), .ZN(new_n1064));
  OAI211_X1 g0864(.A(G330), .B(new_n823), .C1(new_n1064), .C2(new_n712), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n902), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n901), .B1(new_n1066), .B2(new_n1057), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1066), .A2(new_n1057), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1061), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1063), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1071), .A2(new_n675), .A3(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1059), .A2(new_n722), .A3(new_n1060), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n726), .B1(new_n306), .B2(new_n816), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n752), .A2(G283), .B1(G97), .B2(new_n767), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n350), .B2(new_n756), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT117), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n208), .A2(new_n738), .B1(new_n739), .B2(new_n589), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n276), .B1(new_n734), .B2(new_n463), .C1(new_n730), .C2(new_n482), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(G77), .C2(new_n966), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(KEYINPUT54), .B(G143), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n276), .B1(new_n767), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n739), .A2(new_n307), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT53), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n798), .A2(G132), .B1(new_n763), .B2(G125), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n966), .A2(G159), .B1(new_n810), .B2(G50), .ZN(new_n1089));
  AND4_X1   g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G128), .A2(new_n752), .B1(new_n755), .B2(G137), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1079), .A2(new_n1082), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n897), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1076), .B1(new_n728), .B2(new_n1092), .C1(new_n1093), .C2(new_n775), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT118), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1074), .A2(new_n1075), .A3(new_n1095), .ZN(G378));
  INV_X1    g0896(.A(new_n1063), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1073), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT123), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1073), .A2(KEYINPUT123), .A3(new_n1097), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n906), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n331), .A2(new_n656), .ZN(new_n1104));
  AND2_X1   g0904(.A1(new_n336), .A2(new_n338), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1105), .B2(new_n327), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1104), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n339), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1109), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n339), .A2(new_n1107), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n327), .B(new_n1104), .C1(new_n336), .C2(new_n338), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n888), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1110), .A2(new_n1114), .A3(KEYINPUT122), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT122), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n716), .B(new_n1119), .C1(new_n876), .C2(new_n887), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1103), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1119), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n888), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1123), .B(new_n906), .C1(new_n888), .C2(new_n1115), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1121), .A2(new_n1124), .A3(KEYINPUT57), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n676), .B1(new_n1102), .B2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1073), .A2(KEYINPUT123), .A3(new_n1097), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT123), .B1(new_n1073), .B2(new_n1097), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT57), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1126), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1127), .A2(new_n722), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n723), .B1(G50), .B2(new_n817), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT121), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n268), .A2(G41), .ZN(new_n1137));
  AOI211_X1 g0937(.A(G50), .B(new_n1137), .C1(new_n263), .C2(new_n264), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n743), .A2(new_n208), .B1(new_n738), .B2(new_n364), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n798), .A2(G107), .B1(new_n767), .B2(new_n606), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n737), .B2(new_n734), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n752), .C2(G116), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1137), .B1(new_n251), .B2(new_n739), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT119), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(new_n485), .C2(new_n756), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT58), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1138), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n743), .A2(new_n307), .B1(new_n745), .B2(new_n802), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n752), .B2(G125), .ZN(new_n1149));
  INV_X1    g0949(.A(G128), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n730), .A2(new_n1150), .B1(new_n739), .B2(new_n1083), .ZN(new_n1151));
  XOR2_X1   g0951(.A(new_n1151), .B(KEYINPUT120), .Z(new_n1152));
  OAI211_X1 g0952(.A(new_n1149), .B(new_n1152), .C1(new_n806), .C2(new_n756), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n810), .A2(G159), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1147), .B1(new_n1146), .B2(new_n1145), .C1(new_n1154), .C2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1136), .B1(new_n1159), .B2(new_n727), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1122), .B2(new_n775), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1134), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1133), .A2(new_n1163), .ZN(G375));
  AOI21_X1  g0964(.A(new_n726), .B1(new_n208), .B2(new_n816), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G132), .A2(new_n752), .B1(new_n755), .B2(new_n1084), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n745), .A2(new_n307), .B1(new_n734), .B2(new_n1150), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n276), .B(new_n1167), .C1(G137), .C2(new_n798), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n743), .A2(new_n313), .B1(new_n738), .B2(new_n364), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G159), .B2(new_n770), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1166), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G116), .A2(new_n755), .B1(new_n752), .B2(G294), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n745), .A2(new_n350), .B1(new_n734), .B2(new_n740), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n268), .B(new_n1173), .C1(G283), .C2(new_n798), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n965), .B(new_n993), .C1(G97), .C2(new_n770), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1177), .A2(KEYINPUT125), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT125), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n727), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n774), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1165), .B1(new_n1178), .B2(new_n1180), .C1(new_n875), .C2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n1070), .B2(new_n721), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n941), .B(KEYINPUT124), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1072), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1070), .A2(new_n1063), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1183), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(G381));
  INV_X1    g0988(.A(G390), .ZN(new_n1189));
  INV_X1    g0989(.A(G384), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(G393), .A2(G396), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1187), .A4(new_n1191), .ZN(new_n1192));
  OR4_X1    g0992(.A1(G387), .A2(new_n1192), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g0993(.A1(new_n657), .A2(G213), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(G375), .A2(G378), .A3(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT126), .Z(new_n1196));
  NAND3_X1  g0996(.A1(G407), .A2(new_n1196), .A3(G213), .ZN(G409));
  NAND3_X1  g0997(.A1(new_n957), .A2(new_n981), .A3(G390), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(G390), .B1(new_n957), .B2(new_n981), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(G393), .A2(G396), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(new_n1191), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1199), .A2(new_n1200), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(G387), .A2(new_n1189), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1203), .B1(new_n1206), .B2(new_n1198), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT61), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT60), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1072), .A2(new_n1186), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(new_n676), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1186), .B1(new_n1072), .B2(new_n1210), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1183), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(G384), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1194), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(G2897), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1215), .B(new_n1217), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1130), .A2(new_n1184), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G378), .B1(new_n1219), .B2(new_n1163), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1102), .B2(new_n1127), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1125), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n675), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G378), .B(new_n1163), .C1(new_n1221), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT127), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT127), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1133), .A2(new_n1226), .A3(G378), .A4(new_n1163), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1220), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1218), .B1(new_n1228), .B2(new_n1216), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1228), .A2(new_n1216), .A3(new_n1215), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1209), .B(new_n1229), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1220), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1215), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1194), .A3(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(KEYINPUT62), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1208), .B1(new_n1232), .B2(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1229), .A2(new_n1209), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT63), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1230), .A2(KEYINPUT63), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1240), .A2(new_n1241), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1239), .A2(new_n1245), .ZN(G405));
  INV_X1    g1046(.A(G378), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G375), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1233), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(new_n1215), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(new_n1241), .ZN(G402));
endmodule


