

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730;

  NOR2_X1 U376 ( .A1(n649), .A2(n634), .ZN(n578) );
  AND2_X1 U377 ( .A1(n671), .A2(n670), .ZN(n543) );
  AND2_X1 U378 ( .A1(n577), .A2(n576), .ZN(n634) );
  XNOR2_X1 U379 ( .A(n497), .B(KEYINPUT104), .ZN(n645) );
  XNOR2_X1 U380 ( .A(n551), .B(n550), .ZN(n728) );
  AND2_X4 U381 ( .A1(n693), .A2(n597), .ZN(n696) );
  XNOR2_X1 U382 ( .A(n486), .B(KEYINPUT1), .ZN(n667) );
  NOR2_X2 U383 ( .A1(n495), .A2(n506), .ZN(n496) );
  AND2_X1 U384 ( .A1(n506), .A2(n495), .ZN(n497) );
  XNOR2_X2 U385 ( .A(n457), .B(n456), .ZN(n506) );
  XNOR2_X2 U386 ( .A(n589), .B(KEYINPUT45), .ZN(n707) );
  AND2_X1 U387 ( .A1(n423), .A2(n422), .ZN(n509) );
  XNOR2_X1 U388 ( .A(n542), .B(n541), .ZN(n572) );
  NOR2_X1 U389 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U390 ( .A(G143), .B(G113), .ZN(n446) );
  NAND2_X1 U391 ( .A1(n533), .A2(n532), .ZN(n591) );
  NOR2_X1 U392 ( .A1(n631), .A2(n579), .ZN(n580) );
  OR2_X1 U393 ( .A1(n698), .A2(G902), .ZN(n396) );
  OR2_X1 U394 ( .A1(n604), .A2(G902), .ZN(n409) );
  XNOR2_X1 U395 ( .A(n558), .B(n557), .ZN(n568) );
  XNOR2_X1 U396 ( .A(n556), .B(KEYINPUT71), .ZN(n557) );
  INV_X1 U397 ( .A(KEYINPUT22), .ZN(n556) );
  NAND2_X1 U398 ( .A1(n595), .A2(n594), .ZN(n693) );
  INV_X1 U399 ( .A(KEYINPUT64), .ZN(n382) );
  AND2_X1 U400 ( .A1(n543), .A2(n667), .ZN(n571) );
  XNOR2_X1 U401 ( .A(KEYINPUT15), .B(G902), .ZN(n596) );
  XNOR2_X1 U402 ( .A(n388), .B(n387), .ZN(n389) );
  INV_X1 U403 ( .A(G107), .ZN(n387) );
  XNOR2_X1 U404 ( .A(n591), .B(n534), .ZN(n716) );
  AND2_X1 U405 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X2 U406 ( .A(G953), .ZN(n720) );
  OR2_X1 U407 ( .A1(n667), .A2(n566), .ZN(n567) );
  XNOR2_X1 U408 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U409 ( .A(n445), .B(n444), .Z(n354) );
  XOR2_X1 U410 ( .A(n446), .B(KEYINPUT97), .Z(n355) );
  XOR2_X1 U411 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n356) );
  XOR2_X1 U412 ( .A(n604), .B(KEYINPUT62), .Z(n357) );
  OR2_X1 U413 ( .A1(n552), .A2(n670), .ZN(n358) );
  INV_X1 U414 ( .A(KEYINPUT70), .ZN(n399) );
  XNOR2_X1 U415 ( .A(n359), .B(KEYINPUT92), .ZN(n361) );
  XNOR2_X1 U416 ( .A(G128), .B(G137), .ZN(n364) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n376) );
  XNOR2_X1 U418 ( .A(n377), .B(KEYINPUT91), .ZN(n378) );
  XNOR2_X1 U419 ( .A(n383), .B(n459), .ZN(n437) );
  XNOR2_X1 U420 ( .A(n389), .B(n452), .ZN(n392) );
  NOR2_X1 U421 ( .A1(n490), .A2(n525), .ZN(n485) );
  XNOR2_X1 U422 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U423 ( .A(n437), .B(n385), .ZN(n718) );
  XNOR2_X1 U424 ( .A(n718), .B(n386), .ZN(n408) );
  NOR2_X1 U425 ( .A1(n574), .A2(n688), .ZN(n546) );
  XNOR2_X1 U426 ( .A(n398), .B(n397), .ZN(n575) );
  BUF_X1 U427 ( .A(n716), .Z(n719) );
  INV_X1 U428 ( .A(n547), .ZN(n548) );
  INV_X1 U429 ( .A(n702), .ZN(n606) );
  XNOR2_X1 U430 ( .A(n698), .B(n697), .ZN(n699) );
  INV_X1 U431 ( .A(KEYINPUT35), .ZN(n550) );
  INV_X1 U432 ( .A(KEYINPUT121), .ZN(n602) );
  XOR2_X1 U433 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n359) );
  NAND2_X1 U434 ( .A1(G234), .A2(n596), .ZN(n360) );
  AND2_X1 U435 ( .A1(n376), .A2(G221), .ZN(n363) );
  INV_X1 U436 ( .A(KEYINPUT21), .ZN(n362) );
  XNOR2_X1 U437 ( .A(n363), .B(n362), .ZN(n553) );
  INV_X1 U438 ( .A(n553), .ZN(n671) );
  XNOR2_X1 U439 ( .A(n364), .B(KEYINPUT23), .ZN(n366) );
  XNOR2_X1 U440 ( .A(KEYINPUT89), .B(KEYINPUT90), .ZN(n365) );
  XNOR2_X1 U441 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U442 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n368) );
  NAND2_X1 U443 ( .A1(G234), .A2(n720), .ZN(n367) );
  XNOR2_X1 U444 ( .A(n368), .B(n367), .ZN(n462) );
  NAND2_X1 U445 ( .A1(n462), .A2(G221), .ZN(n369) );
  XNOR2_X1 U446 ( .A(n370), .B(n369), .ZN(n375) );
  XNOR2_X1 U447 ( .A(G146), .B(G125), .ZN(n430) );
  XNOR2_X1 U448 ( .A(n430), .B(KEYINPUT10), .ZN(n453) );
  XNOR2_X1 U449 ( .A(G119), .B(G140), .ZN(n372) );
  XNOR2_X1 U450 ( .A(G110), .B(KEYINPUT24), .ZN(n371) );
  XNOR2_X1 U451 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U452 ( .A(n453), .B(n373), .ZN(n374) );
  XNOR2_X1 U453 ( .A(n375), .B(n374), .ZN(n612) );
  INV_X1 U454 ( .A(G902), .ZN(n455) );
  NAND2_X1 U455 ( .A1(n612), .A2(n455), .ZN(n381) );
  AND2_X1 U456 ( .A1(G217), .A2(n376), .ZN(n379) );
  XOR2_X1 U457 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n377) );
  XNOR2_X2 U458 ( .A(n381), .B(n380), .ZN(n670) );
  XNOR2_X1 U459 ( .A(n382), .B(KEYINPUT4), .ZN(n383) );
  XNOR2_X2 U460 ( .A(G143), .B(G128), .ZN(n459) );
  XNOR2_X1 U461 ( .A(G134), .B(G137), .ZN(n384) );
  XNOR2_X1 U462 ( .A(n384), .B(KEYINPUT67), .ZN(n385) );
  XNOR2_X1 U463 ( .A(KEYINPUT65), .B(G101), .ZN(n431) );
  XNOR2_X1 U464 ( .A(n431), .B(G146), .ZN(n386) );
  NAND2_X1 U465 ( .A1(G227), .A2(n720), .ZN(n388) );
  XOR2_X1 U466 ( .A(G131), .B(G140), .Z(n452) );
  XNOR2_X1 U467 ( .A(G110), .B(G104), .ZN(n390) );
  XNOR2_X1 U468 ( .A(n390), .B(KEYINPUT85), .ZN(n426) );
  INV_X1 U469 ( .A(n426), .ZN(n391) );
  XNOR2_X1 U470 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U471 ( .A(n408), .B(n393), .ZN(n698) );
  INV_X1 U472 ( .A(KEYINPUT69), .ZN(n394) );
  XNOR2_X1 U473 ( .A(n394), .B(G469), .ZN(n395) );
  XNOR2_X2 U474 ( .A(n396), .B(n395), .ZN(n486) );
  NAND2_X1 U475 ( .A1(n543), .A2(n486), .ZN(n398) );
  INV_X1 U476 ( .A(KEYINPUT95), .ZN(n397) );
  XNOR2_X1 U477 ( .A(n575), .B(KEYINPUT107), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n399), .B(KEYINPUT3), .ZN(n401) );
  XNOR2_X1 U479 ( .A(G119), .B(G113), .ZN(n400) );
  XNOR2_X1 U480 ( .A(n401), .B(n400), .ZN(n425) );
  NOR2_X1 U481 ( .A1(G953), .A2(G237), .ZN(n449) );
  NAND2_X1 U482 ( .A1(n449), .A2(G210), .ZN(n403) );
  XNOR2_X1 U483 ( .A(G131), .B(G116), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n403), .B(n402), .ZN(n405) );
  XNOR2_X1 U485 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n404) );
  XNOR2_X1 U486 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U487 ( .A(n425), .B(n406), .ZN(n407) );
  XNOR2_X1 U488 ( .A(n408), .B(n407), .ZN(n604) );
  XNOR2_X2 U489 ( .A(n409), .B(G472), .ZN(n673) );
  NOR2_X1 U490 ( .A1(G237), .A2(G902), .ZN(n410) );
  XNOR2_X1 U491 ( .A(n410), .B(KEYINPUT73), .ZN(n439) );
  AND2_X1 U492 ( .A1(n439), .A2(G214), .ZN(n412) );
  INV_X1 U493 ( .A(KEYINPUT86), .ZN(n411) );
  XNOR2_X1 U494 ( .A(n412), .B(n411), .ZN(n484) );
  NAND2_X1 U495 ( .A1(n673), .A2(n484), .ZN(n414) );
  XNOR2_X1 U496 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n413) );
  XNOR2_X1 U497 ( .A(n414), .B(n413), .ZN(n421) );
  XOR2_X1 U498 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n416) );
  NAND2_X1 U499 ( .A1(G237), .A2(G234), .ZN(n415) );
  XNOR2_X1 U500 ( .A(n416), .B(n415), .ZN(n417) );
  NAND2_X1 U501 ( .A1(G952), .A2(n417), .ZN(n686) );
  NOR2_X1 U502 ( .A1(G953), .A2(n686), .ZN(n538) );
  NAND2_X1 U503 ( .A1(G902), .A2(n417), .ZN(n536) );
  OR2_X1 U504 ( .A1(n720), .A2(n536), .ZN(n418) );
  NOR2_X1 U505 ( .A1(G900), .A2(n418), .ZN(n419) );
  OR2_X1 U506 ( .A1(n538), .A2(n419), .ZN(n420) );
  XNOR2_X1 U507 ( .A(n420), .B(KEYINPUT77), .ZN(n473) );
  NOR2_X1 U508 ( .A1(n421), .A2(n473), .ZN(n422) );
  XNOR2_X1 U509 ( .A(G116), .B(G107), .ZN(n424) );
  XNOR2_X1 U510 ( .A(n424), .B(G122), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n425), .B(n461), .ZN(n429) );
  INV_X1 U512 ( .A(KEYINPUT16), .ZN(n427) );
  XNOR2_X1 U513 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U514 ( .A(n429), .B(n428), .ZN(n703) );
  XNOR2_X1 U515 ( .A(n431), .B(n430), .ZN(n435) );
  NAND2_X1 U516 ( .A1(G224), .A2(n720), .ZN(n433) );
  XNOR2_X1 U517 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n432) );
  XNOR2_X1 U518 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U519 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U520 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U521 ( .A(n703), .B(n438), .ZN(n625) );
  NAND2_X1 U522 ( .A1(n625), .A2(n596), .ZN(n441) );
  NAND2_X1 U523 ( .A1(G210), .A2(n439), .ZN(n440) );
  XNOR2_X2 U524 ( .A(n441), .B(n440), .ZN(n490) );
  INV_X1 U525 ( .A(KEYINPUT38), .ZN(n442) );
  XNOR2_X1 U526 ( .A(n490), .B(n442), .ZN(n658) );
  INV_X1 U527 ( .A(n658), .ZN(n443) );
  NAND2_X1 U528 ( .A1(n509), .A2(n443), .ZN(n445) );
  INV_X1 U529 ( .A(KEYINPUT39), .ZN(n444) );
  XNOR2_X1 U530 ( .A(G122), .B(G104), .ZN(n447) );
  XNOR2_X1 U531 ( .A(n356), .B(n447), .ZN(n448) );
  XNOR2_X1 U532 ( .A(n355), .B(n448), .ZN(n451) );
  NAND2_X1 U533 ( .A1(n449), .A2(G214), .ZN(n450) );
  XNOR2_X1 U534 ( .A(n451), .B(n450), .ZN(n454) );
  XNOR2_X1 U535 ( .A(n453), .B(n452), .ZN(n717) );
  XNOR2_X1 U536 ( .A(n454), .B(n717), .ZN(n617) );
  NAND2_X1 U537 ( .A1(n617), .A2(n455), .ZN(n457) );
  XOR2_X1 U538 ( .A(KEYINPUT13), .B(G475), .Z(n456) );
  XOR2_X1 U539 ( .A(KEYINPUT98), .B(G134), .Z(n458) );
  XNOR2_X1 U540 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U541 ( .A(n461), .B(n460), .ZN(n466) );
  XOR2_X1 U542 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n464) );
  NAND2_X1 U543 ( .A1(G217), .A2(n462), .ZN(n463) );
  XNOR2_X1 U544 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U545 ( .A(n466), .B(n465), .ZN(n598) );
  NOR2_X1 U546 ( .A1(n598), .A2(G902), .ZN(n467) );
  XNOR2_X1 U547 ( .A(G478), .B(n467), .ZN(n495) );
  NAND2_X1 U548 ( .A1(n354), .A2(n497), .ZN(n469) );
  INV_X1 U549 ( .A(KEYINPUT40), .ZN(n468) );
  XNOR2_X1 U550 ( .A(n469), .B(n468), .ZN(n611) );
  INV_X1 U551 ( .A(n484), .ZN(n657) );
  NOR2_X1 U552 ( .A1(n658), .A2(n657), .ZN(n470) );
  XNOR2_X1 U553 ( .A(n470), .B(KEYINPUT109), .ZN(n662) );
  INV_X1 U554 ( .A(n495), .ZN(n505) );
  NOR2_X1 U555 ( .A1(n506), .A2(n505), .ZN(n471) );
  XNOR2_X1 U556 ( .A(KEYINPUT101), .B(n471), .ZN(n661) );
  NOR2_X1 U557 ( .A1(n662), .A2(n661), .ZN(n472) );
  XNOR2_X1 U558 ( .A(n472), .B(KEYINPUT41), .ZN(n687) );
  NOR2_X1 U559 ( .A1(n473), .A2(n553), .ZN(n474) );
  XOR2_X1 U560 ( .A(KEYINPUT68), .B(n474), .Z(n475) );
  NOR2_X1 U561 ( .A1(n475), .A2(n670), .ZN(n481) );
  NAND2_X1 U562 ( .A1(n481), .A2(n673), .ZN(n477) );
  INV_X1 U563 ( .A(KEYINPUT28), .ZN(n476) );
  XNOR2_X1 U564 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U565 ( .A1(n478), .A2(n486), .ZN(n493) );
  NOR2_X1 U566 ( .A1(n687), .A2(n493), .ZN(n479) );
  XNOR2_X1 U567 ( .A(n479), .B(KEYINPUT42), .ZN(n730) );
  NOR2_X2 U568 ( .A1(n611), .A2(n730), .ZN(n480) );
  XNOR2_X1 U569 ( .A(n480), .B(KEYINPUT46), .ZN(n522) );
  NAND2_X1 U570 ( .A1(n645), .A2(n481), .ZN(n482) );
  XNOR2_X1 U571 ( .A(n673), .B(KEYINPUT6), .ZN(n570) );
  NOR2_X1 U572 ( .A1(n482), .A2(n570), .ZN(n483) );
  NAND2_X1 U573 ( .A1(n484), .A2(n483), .ZN(n525) );
  XOR2_X1 U574 ( .A(KEYINPUT36), .B(n485), .Z(n488) );
  INV_X1 U575 ( .A(n667), .ZN(n487) );
  NOR2_X1 U576 ( .A1(n488), .A2(n487), .ZN(n652) );
  INV_X1 U577 ( .A(KEYINPUT82), .ZN(n489) );
  XNOR2_X1 U578 ( .A(n652), .B(n489), .ZN(n520) );
  NOR2_X1 U579 ( .A1(n490), .A2(n657), .ZN(n492) );
  XNOR2_X1 U580 ( .A(KEYINPUT74), .B(KEYINPUT19), .ZN(n491) );
  XNOR2_X1 U581 ( .A(n492), .B(n491), .ZN(n540) );
  NOR2_X1 U582 ( .A1(n540), .A2(n493), .ZN(n494) );
  XOR2_X1 U583 ( .A(KEYINPUT76), .B(n494), .Z(n638) );
  XOR2_X1 U584 ( .A(KEYINPUT99), .B(n496), .Z(n648) );
  XNOR2_X1 U585 ( .A(n648), .B(KEYINPUT100), .ZN(n531) );
  NOR2_X2 U586 ( .A1(n497), .A2(n531), .ZN(n663) );
  XOR2_X1 U587 ( .A(KEYINPUT72), .B(n663), .Z(n499) );
  INV_X1 U588 ( .A(KEYINPUT47), .ZN(n498) );
  NAND2_X1 U589 ( .A1(n499), .A2(n498), .ZN(n500) );
  NOR2_X1 U590 ( .A1(n638), .A2(n500), .ZN(n518) );
  AND2_X1 U591 ( .A1(n663), .A2(KEYINPUT78), .ZN(n501) );
  NOR2_X1 U592 ( .A1(n638), .A2(n501), .ZN(n502) );
  NAND2_X1 U593 ( .A1(KEYINPUT72), .A2(n502), .ZN(n503) );
  NAND2_X1 U594 ( .A1(n503), .A2(KEYINPUT47), .ZN(n516) );
  NAND2_X1 U595 ( .A1(n663), .A2(KEYINPUT47), .ZN(n504) );
  INV_X1 U596 ( .A(KEYINPUT78), .ZN(n511) );
  NAND2_X1 U597 ( .A1(n504), .A2(n511), .ZN(n510) );
  NAND2_X1 U598 ( .A1(n506), .A2(n505), .ZN(n507) );
  XOR2_X1 U599 ( .A(KEYINPUT103), .B(n507), .Z(n547) );
  NOR2_X1 U600 ( .A1(n547), .A2(n490), .ZN(n508) );
  NAND2_X1 U601 ( .A1(n509), .A2(n508), .ZN(n642) );
  NAND2_X1 U602 ( .A1(n510), .A2(n642), .ZN(n514) );
  INV_X1 U603 ( .A(n642), .ZN(n512) );
  NAND2_X1 U604 ( .A1(n512), .A2(n511), .ZN(n513) );
  NAND2_X1 U605 ( .A1(n514), .A2(n513), .ZN(n515) );
  NAND2_X1 U606 ( .A1(n516), .A2(n515), .ZN(n517) );
  NOR2_X1 U607 ( .A1(n518), .A2(n517), .ZN(n519) );
  AND2_X1 U608 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U609 ( .A1(n522), .A2(n521), .ZN(n524) );
  INV_X1 U610 ( .A(KEYINPUT48), .ZN(n523) );
  XNOR2_X1 U611 ( .A(n524), .B(n523), .ZN(n533) );
  XNOR2_X1 U612 ( .A(KEYINPUT105), .B(n525), .ZN(n526) );
  NAND2_X1 U613 ( .A1(n526), .A2(n487), .ZN(n527) );
  XOR2_X1 U614 ( .A(n527), .B(KEYINPUT106), .Z(n528) );
  XNOR2_X1 U615 ( .A(n528), .B(KEYINPUT43), .ZN(n530) );
  INV_X1 U616 ( .A(n490), .ZN(n529) );
  NOR2_X1 U617 ( .A1(n530), .A2(n529), .ZN(n655) );
  AND2_X1 U618 ( .A1(n354), .A2(n531), .ZN(n609) );
  NOR2_X1 U619 ( .A1(n655), .A2(n609), .ZN(n532) );
  INV_X1 U620 ( .A(KEYINPUT80), .ZN(n534) );
  INV_X1 U621 ( .A(KEYINPUT2), .ZN(n535) );
  AND2_X1 U622 ( .A1(n716), .A2(n535), .ZN(n590) );
  OR2_X1 U623 ( .A1(n720), .A2(G898), .ZN(n704) );
  NOR2_X1 U624 ( .A1(n536), .A2(n704), .ZN(n537) );
  NOR2_X1 U625 ( .A1(n538), .A2(n537), .ZN(n539) );
  INV_X1 U626 ( .A(KEYINPUT0), .ZN(n541) );
  XNOR2_X1 U627 ( .A(KEYINPUT88), .B(n572), .ZN(n574) );
  INV_X1 U628 ( .A(n570), .ZN(n544) );
  NAND2_X1 U629 ( .A1(n571), .A2(n544), .ZN(n545) );
  XOR2_X1 U630 ( .A(KEYINPUT33), .B(n545), .Z(n688) );
  XNOR2_X1 U631 ( .A(n546), .B(KEYINPUT34), .ZN(n549) );
  NAND2_X1 U632 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT75), .ZN(n552) );
  OR2_X1 U634 ( .A1(n487), .A2(n358), .ZN(n559) );
  INV_X1 U635 ( .A(n661), .ZN(n555) );
  NOR2_X1 U636 ( .A1(n572), .A2(n553), .ZN(n554) );
  NAND2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n558) );
  NOR2_X1 U638 ( .A1(n559), .A2(n568), .ZN(n560) );
  XNOR2_X1 U639 ( .A(n560), .B(KEYINPUT32), .ZN(n729) );
  NOR2_X1 U640 ( .A1(n673), .A2(n670), .ZN(n561) );
  NAND2_X1 U641 ( .A1(n487), .A2(n561), .ZN(n562) );
  NOR2_X1 U642 ( .A1(n568), .A2(n562), .ZN(n610) );
  NOR2_X1 U643 ( .A1(n729), .A2(n610), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n728), .A2(n583), .ZN(n563) );
  XNOR2_X1 U645 ( .A(n563), .B(KEYINPUT44), .ZN(n565) );
  INV_X1 U646 ( .A(KEYINPUT83), .ZN(n564) );
  NAND2_X1 U647 ( .A1(n565), .A2(n564), .ZN(n588) );
  INV_X1 U648 ( .A(n670), .ZN(n566) );
  NOR2_X1 U649 ( .A1(n568), .A2(n567), .ZN(n569) );
  AND2_X1 U650 ( .A1(n570), .A2(n569), .ZN(n631) );
  NAND2_X1 U651 ( .A1(n571), .A2(n673), .ZN(n677) );
  NOR2_X1 U652 ( .A1(n572), .A2(n677), .ZN(n573) );
  XOR2_X1 U653 ( .A(KEYINPUT31), .B(n573), .Z(n649) );
  INV_X1 U654 ( .A(n574), .ZN(n577) );
  NOR2_X1 U655 ( .A1(n575), .A2(n673), .ZN(n576) );
  NOR2_X1 U656 ( .A1(n663), .A2(n578), .ZN(n579) );
  XNOR2_X1 U657 ( .A(n580), .B(KEYINPUT102), .ZN(n582) );
  NAND2_X1 U658 ( .A1(KEYINPUT83), .A2(n728), .ZN(n581) );
  AND2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U660 ( .A1(KEYINPUT44), .A2(n583), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n584), .A2(KEYINPUT83), .ZN(n585) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n707), .ZN(n595) );
  INV_X1 U664 ( .A(n591), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n707), .A2(n592), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n593), .A2(KEYINPUT2), .ZN(n594) );
  INV_X1 U667 ( .A(n596), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n696), .A2(G478), .ZN(n599) );
  XNOR2_X1 U669 ( .A(n599), .B(n598), .ZN(n601) );
  INV_X1 U670 ( .A(G952), .ZN(n600) );
  AND2_X1 U671 ( .A1(n600), .A2(G953), .ZN(n702) );
  NOR2_X2 U672 ( .A1(n601), .A2(n702), .ZN(n603) );
  XNOR2_X1 U673 ( .A(n603), .B(n602), .ZN(G63) );
  NAND2_X1 U674 ( .A1(n696), .A2(G472), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n605), .B(n357), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U677 ( .A(n608), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U678 ( .A(G134), .B(n609), .Z(G36) );
  XOR2_X1 U679 ( .A(n610), .B(G110), .Z(G12) );
  XOR2_X1 U680 ( .A(n611), .B(G131), .Z(G33) );
  NAND2_X1 U681 ( .A1(n696), .A2(G217), .ZN(n614) );
  XOR2_X1 U682 ( .A(KEYINPUT122), .B(n612), .Z(n613) );
  XNOR2_X1 U683 ( .A(n614), .B(n613), .ZN(n615) );
  NOR2_X1 U684 ( .A1(n615), .A2(n702), .ZN(G66) );
  NAND2_X1 U685 ( .A1(n696), .A2(G475), .ZN(n619) );
  XNOR2_X1 U686 ( .A(KEYINPUT120), .B(KEYINPUT59), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X2 U689 ( .A1(n620), .A2(n702), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n621), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U691 ( .A1(n696), .A2(G210), .ZN(n627) );
  XOR2_X1 U692 ( .A(KEYINPUT84), .B(KEYINPUT79), .Z(n623) );
  XNOR2_X1 U693 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n622) );
  XNOR2_X1 U694 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U696 ( .A(n627), .B(n626), .ZN(n628) );
  NOR2_X2 U697 ( .A1(n628), .A2(n702), .ZN(n630) );
  XOR2_X1 U698 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G51) );
  XOR2_X1 U700 ( .A(G101), .B(n631), .Z(G3) );
  NAND2_X1 U701 ( .A1(n634), .A2(n645), .ZN(n632) );
  XNOR2_X1 U702 ( .A(n632), .B(KEYINPUT110), .ZN(n633) );
  XNOR2_X1 U703 ( .A(G104), .B(n633), .ZN(G6) );
  XOR2_X1 U704 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n636) );
  NAND2_X1 U705 ( .A1(n634), .A2(n648), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U707 ( .A(G107), .B(n637), .ZN(G9) );
  XOR2_X1 U708 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n640) );
  INV_X1 U709 ( .A(n638), .ZN(n643) );
  NAND2_X1 U710 ( .A1(n648), .A2(n643), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(n641) );
  XOR2_X1 U712 ( .A(G128), .B(n641), .Z(G30) );
  XNOR2_X1 U713 ( .A(G143), .B(n642), .ZN(G45) );
  NAND2_X1 U714 ( .A1(n643), .A2(n645), .ZN(n644) );
  XNOR2_X1 U715 ( .A(n644), .B(G146), .ZN(G48) );
  NAND2_X1 U716 ( .A1(n645), .A2(n649), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n646), .B(KEYINPUT112), .ZN(n647) );
  XNOR2_X1 U718 ( .A(G113), .B(n647), .ZN(G15) );
  XOR2_X1 U719 ( .A(G116), .B(KEYINPUT113), .Z(n651) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(G18) );
  XNOR2_X1 U722 ( .A(n652), .B(KEYINPUT114), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(KEYINPUT37), .ZN(n654) );
  XNOR2_X1 U724 ( .A(G125), .B(n654), .ZN(G27) );
  XNOR2_X1 U725 ( .A(G140), .B(n655), .ZN(n656) );
  XNOR2_X1 U726 ( .A(n656), .B(KEYINPUT115), .ZN(G42) );
  NAND2_X1 U727 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U728 ( .A(KEYINPUT118), .B(n659), .Z(n660) );
  NOR2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n666), .A2(n688), .ZN(n683) );
  NOR2_X1 U733 ( .A1(n667), .A2(n543), .ZN(n669) );
  XOR2_X1 U734 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n668) );
  XNOR2_X1 U735 ( .A(n669), .B(n668), .ZN(n676) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT49), .B(n672), .Z(n674) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n680) );
  XOR2_X1 U741 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n679) );
  XNOR2_X1 U742 ( .A(n680), .B(n679), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n681), .A2(n687), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n691) );
  NOR2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U748 ( .A(n689), .B(KEYINPUT119), .Z(n690) );
  OR2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U750 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U751 ( .A1(n694), .A2(G953), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n695), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U753 ( .A1(n696), .A2(G469), .ZN(n700) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n697) );
  NOR2_X1 U755 ( .A1(n702), .A2(n701), .ZN(G54) );
  XNOR2_X1 U756 ( .A(n703), .B(G101), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n706), .B(KEYINPUT125), .ZN(n715) );
  NAND2_X1 U759 ( .A1(n707), .A2(n720), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n708), .B(KEYINPUT124), .ZN(n713) );
  XOR2_X1 U761 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n710) );
  NAND2_X1 U762 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U763 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U764 ( .A1(n711), .A2(G898), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(G69) );
  XOR2_X1 U767 ( .A(n718), .B(n717), .Z(n722) );
  XNOR2_X1 U768 ( .A(n719), .B(n722), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n721), .A2(n720), .ZN(n727) );
  XOR2_X1 U770 ( .A(G227), .B(n722), .Z(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(G900), .ZN(n724) );
  XNOR2_X1 U772 ( .A(KEYINPUT126), .B(n724), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n725), .A2(G953), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n727), .A2(n726), .ZN(G72) );
  XNOR2_X1 U775 ( .A(n728), .B(G122), .ZN(G24) );
  XOR2_X1 U776 ( .A(G119), .B(n729), .Z(G21) );
  XOR2_X1 U777 ( .A(G137), .B(n730), .Z(G39) );
endmodule

