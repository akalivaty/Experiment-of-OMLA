//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT95), .ZN(new_n204));
  AOI21_X1  g003(.A(G8gat), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n205), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210));
  XOR2_X1   g009(.A(G57gat), .B(G64gat), .Z(new_n211));
  XNOR2_X1  g010(.A(G71gat), .B(G78gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT98), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT98), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n211), .A2(new_n218), .A3(new_n212), .A4(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(new_n215), .ZN(new_n221));
  NOR2_X1   g020(.A1(G71gat), .A2(G78gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT97), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(new_n213), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n221), .B(new_n224), .C1(new_n223), .C2(new_n213), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n227), .A2(KEYINPUT100), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(KEYINPUT100), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G231gat), .A2(G233gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT99), .ZN(new_n232));
  XOR2_X1   g031(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n233));
  XOR2_X1   g032(.A(new_n232), .B(new_n233), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n234), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n229), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n226), .A2(new_n210), .ZN(new_n239));
  XOR2_X1   g038(.A(G127gat), .B(G155gat), .Z(new_n240));
  XNOR2_X1  g039(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(G183gat), .B(G211gat), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n235), .A3(new_n237), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n248));
  NAND3_X1  g047(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n249), .ZN(new_n251));
  NAND2_X1  g050(.A1(G99gat), .A2(G106gat), .ZN(new_n252));
  INV_X1    g051(.A(G85gat), .ZN(new_n253));
  INV_X1    g052(.A(G92gat), .ZN(new_n254));
  AOI22_X1  g053(.A1(KEYINPUT8), .A2(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n250), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(G99gat), .B(G106gat), .Z(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n250), .A2(new_n259), .A3(new_n251), .A4(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n226), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT10), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n258), .A2(new_n220), .A3(new_n225), .A4(new_n260), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n261), .ZN(new_n266));
  AND2_X1   g065(.A1(new_n220), .A2(new_n225), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT10), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G230gat), .A2(G233gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT104), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(KEYINPUT104), .A3(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n262), .A2(new_n264), .ZN(new_n275));
  INV_X1    g074(.A(new_n270), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n273), .A2(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G120gat), .B(G148gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279));
  XOR2_X1   g078(.A(new_n278), .B(new_n279), .Z(new_n280));
  OR2_X1    g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n282), .A2(KEYINPUT92), .ZN(new_n283));
  OR3_X1    g082(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(KEYINPUT92), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT93), .B(G36gat), .Z(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G29gat), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G43gat), .B(G50gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT15), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n284), .A2(new_n282), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT94), .B(KEYINPUT15), .Z(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(new_n294), .B2(new_n290), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n289), .A2(new_n291), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(G232gat), .A2(G233gat), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n266), .A2(new_n296), .B1(KEYINPUT41), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(KEYINPUT17), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n296), .A2(KEYINPUT17), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n301), .B2(new_n266), .ZN(new_n302));
  XNOR2_X1  g101(.A(G190gat), .B(G218gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT103), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n297), .A2(KEYINPUT41), .ZN(new_n306));
  XNOR2_X1  g105(.A(G134gat), .B(G162gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n304), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n309), .B(new_n298), .C1(new_n301), .C2(new_n266), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n305), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n305), .B2(new_n310), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n280), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n275), .B2(new_n276), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n271), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n247), .A2(new_n281), .A3(new_n313), .A4(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT96), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT25), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT66), .A2(KEYINPUT25), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  INV_X1    g123(.A(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(KEYINPUT24), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT24), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(G183gat), .A3(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n330), .B2(KEYINPUT23), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n339), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n323), .B1(new_n336), .B2(new_n341), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n343));
  AND4_X1   g142(.A1(new_n323), .A2(new_n343), .A3(new_n341), .A4(new_n328), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n322), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT1), .ZN(new_n346));
  INV_X1    g145(.A(G113gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(G120gat), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G127gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT70), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT70), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G127gat), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n353), .A2(new_n355), .A3(G134gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT69), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(new_n352), .B2(G134gat), .ZN(new_n358));
  INV_X1    g157(.A(G134gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n351), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT71), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n364), .B(new_n351), .C1(new_n356), .C2(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n349), .A2(G113gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n347), .A2(G120gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G127gat), .B(G134gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n346), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT72), .A4(new_n346), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT27), .B(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G190gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT68), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT68), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n382), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT27), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G183gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n387));
  AOI21_X1  g186(.A(G190gat), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n387), .B2(new_n377), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n378), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n332), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n392), .A2(KEYINPUT26), .A3(new_n330), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n330), .A2(KEYINPUT26), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n327), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n345), .A2(new_n376), .A3(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n363), .A2(new_n365), .B1(new_n373), .B2(new_n374), .ZN(new_n399));
  INV_X1    g198(.A(new_n323), .ZN(new_n400));
  INV_X1    g199(.A(new_n341), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n328), .A2(new_n332), .A3(new_n334), .A4(new_n331), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n343), .A2(new_n341), .A3(new_n323), .A4(new_n328), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n321), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n396), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n384), .B2(new_n390), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n399), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT64), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n398), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT32), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n417), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n411), .B(KEYINPUT32), .C1(new_n413), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n398), .A2(new_n408), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n409), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n410), .A2(KEYINPUT34), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n423), .A2(KEYINPUT34), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G197gat), .B(G204gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT22), .ZN(new_n429));
  INV_X1    g228(.A(G211gat), .ZN(new_n430));
  INV_X1    g229(.A(G218gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g232(.A(G211gat), .B(G218gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n428), .A3(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OR2_X1    g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(G141gat), .A2(G148gat), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G155gat), .A2(G162gat), .ZN(new_n442));
  INV_X1    g241(.A(G155gat), .ZN(new_n443));
  INV_X1    g242(.A(G162gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(KEYINPUT2), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n441), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT3), .ZN(new_n448));
  OR2_X1    g247(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n449));
  NAND2_X1  g248(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n439), .A2(new_n449), .A3(new_n440), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n442), .A2(KEYINPUT76), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n445), .ZN(new_n454));
  NOR2_X1   g253(.A1(G155gat), .A2(G162gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT76), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n447), .B(new_n448), .C1(new_n452), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT78), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT76), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n460), .A2(G155gat), .A3(G162gat), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n445), .B2(new_n453), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n462), .A2(new_n451), .B1(new_n446), .B2(new_n441), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(new_n448), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT29), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n438), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT3), .B1(new_n438), .B2(new_n467), .ZN(new_n469));
  OAI211_X1 g268(.A(G228gat), .B(G233gat), .C1(new_n469), .C2(new_n463), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT82), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n436), .A2(new_n437), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n448), .B1(new_n473), .B2(KEYINPUT29), .ZN(new_n474));
  INV_X1    g273(.A(new_n463), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT29), .B1(new_n459), .B2(new_n465), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n476), .B(new_n477), .C1(new_n438), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n474), .A2(KEYINPUT81), .A3(new_n475), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT81), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n469), .B2(new_n463), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n472), .B1(new_n484), .B2(new_n468), .ZN(new_n485));
  INV_X1    g284(.A(G22gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT83), .ZN(new_n487));
  XNOR2_X1  g286(.A(G78gat), .B(G106gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT31), .B(G50gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  MUX2_X1   g289(.A(new_n486), .B(new_n487), .S(new_n490), .Z(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n480), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n480), .B2(new_n485), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n418), .A2(new_n425), .A3(new_n420), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n427), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n427), .A2(new_n495), .A3(KEYINPUT89), .A4(new_n496), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT79), .B1(new_n399), .B2(new_n463), .ZN(new_n502));
  INV_X1    g301(.A(new_n365), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n353), .A2(new_n355), .A3(G134gat), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n504), .A2(new_n358), .A3(new_n360), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n364), .B1(new_n505), .B2(new_n351), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n463), .B(new_n375), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT79), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT4), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n507), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n466), .A2(new_n376), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g316(.A1(G225gat), .A2(G233gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n466), .A2(new_n376), .A3(new_n515), .ZN(new_n521));
  INV_X1    g320(.A(new_n518), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n366), .A2(KEYINPUT79), .A3(new_n463), .A4(new_n375), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT4), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT80), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT4), .ZN(new_n528));
  OAI22_X1  g327(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n511), .ZN(new_n529));
  AOI211_X1 g328(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n524), .C2(new_n525), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n523), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n524), .B(new_n525), .C1(new_n463), .C2(new_n399), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n517), .B1(new_n532), .B2(new_n522), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n520), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G1gat), .B(G29gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT0), .ZN(new_n536));
  XNOR2_X1  g335(.A(G57gat), .B(G85gat), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(new_n537), .Z(new_n538));
  AOI21_X1  g337(.A(KEYINPUT6), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  INV_X1    g339(.A(new_n533), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n511), .A2(new_n528), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n528), .B1(new_n502), .B2(new_n509), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT80), .ZN(new_n544));
  INV_X1    g343(.A(new_n530), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n541), .B1(new_n546), .B2(new_n523), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n540), .B1(new_n547), .B2(new_n520), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n539), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(KEYINPUT6), .B(new_n540), .C1(new_n547), .C2(new_n520), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G226gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT73), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n345), .A2(new_n554), .A3(new_n397), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n467), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(new_n405), .B2(new_n407), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n438), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n555), .A2(new_n558), .A3(new_n473), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT74), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n473), .B1(new_n555), .B2(new_n558), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G8gat), .B(G36gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G64gat), .B(G92gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n567), .B(new_n568), .Z(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT75), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AOI211_X1 g372(.A(KEYINPUT74), .B(new_n473), .C1(new_n555), .C2(new_n558), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n555), .A2(new_n558), .A3(new_n473), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(new_n563), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n576), .B2(KEYINPUT74), .ZN(new_n577));
  INV_X1    g376(.A(new_n569), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n562), .B2(new_n565), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT30), .B1(new_n580), .B2(KEYINPUT75), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n501), .A2(new_n551), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n520), .ZN(new_n585));
  INV_X1    g384(.A(new_n523), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n544), .B2(new_n545), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n538), .B(new_n585), .C1(new_n587), .C2(new_n541), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n538), .B(KEYINPUT84), .Z(new_n591));
  NOR2_X1   g390(.A1(new_n534), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n550), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT88), .B(KEYINPUT35), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n582), .A2(new_n497), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n584), .A2(KEYINPUT35), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT87), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n576), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n599), .A2(KEYINPUT38), .A3(new_n569), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT86), .B1(new_n566), .B2(new_n598), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT86), .ZN(new_n602));
  AOI211_X1 g401(.A(new_n602), .B(KEYINPUT37), .C1(new_n562), .C2(new_n565), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n600), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n570), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n597), .B1(new_n593), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n602), .B1(new_n577), .B2(KEYINPUT37), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n566), .A2(KEYINPUT86), .A3(new_n598), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n580), .B1(new_n609), .B2(new_n600), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n588), .B(new_n589), .C1(new_n534), .C2(new_n591), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n610), .A2(KEYINPUT87), .A3(new_n550), .A4(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT38), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n569), .B1(new_n577), .B2(KEYINPUT37), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n606), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n532), .A2(new_n522), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n528), .B1(new_n524), .B2(new_n525), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n619), .A2(new_n521), .A3(new_n512), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n618), .B(KEYINPUT39), .C1(new_n620), .C2(new_n518), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n622), .B(new_n522), .C1(new_n514), .C2(new_n521), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n623), .A3(new_n591), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT85), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT40), .ZN(new_n626));
  INV_X1    g425(.A(new_n592), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT40), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(KEYINPUT85), .A3(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n626), .A2(new_n582), .A3(new_n627), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n495), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n496), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n425), .B1(new_n420), .B2(new_n418), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT36), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT36), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n634), .B2(new_n635), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n582), .B1(new_n549), .B2(new_n550), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n640), .B1(new_n641), .B2(new_n495), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n596), .B1(new_n633), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n209), .B1(new_n299), .B2(new_n300), .ZN(new_n645));
  INV_X1    g444(.A(new_n296), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(new_n209), .ZN(new_n647));
  NAND2_X1  g446(.A1(G229gat), .A2(G233gat), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT18), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n645), .A2(new_n647), .A3(KEYINPUT18), .A4(new_n648), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n646), .B(new_n209), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n648), .B(KEYINPUT13), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT90), .B(G197gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT11), .B(G169gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT91), .B(KEYINPUT12), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n651), .A2(new_n665), .A3(new_n652), .A4(new_n655), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n318), .B1(new_n644), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n584), .A2(KEYINPUT35), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n595), .A2(new_n593), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n611), .A2(new_n550), .A3(new_n570), .A4(new_n604), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n615), .B1(new_n673), .B2(new_n597), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n631), .B1(new_n674), .B2(new_n612), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n675), .B2(new_n642), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n676), .A2(KEYINPUT96), .A3(new_n667), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n317), .B1(new_n669), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n551), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g480(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G8gat), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n678), .A2(new_n582), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(G8gat), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n678), .B2(new_n582), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n678), .A2(new_n582), .A3(new_n683), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(G1325gat));
  INV_X1    g490(.A(new_n678), .ZN(new_n692));
  INV_X1    g491(.A(new_n636), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n692), .A2(G15gat), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n692), .B2(new_n640), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(G1326gat));
  INV_X1    g495(.A(new_n495), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n281), .A2(new_n316), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n701), .A2(new_n247), .ZN(new_n702));
  INV_X1    g501(.A(new_n313), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n669), .B2(new_n677), .ZN(new_n705));
  INV_X1    g504(.A(G29gat), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n679), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n642), .B1(new_n617), .B2(new_n632), .ZN(new_n710));
  OAI211_X1 g509(.A(KEYINPUT44), .B(new_n703), .C1(new_n710), .C2(new_n596), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n676), .B2(new_n703), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n702), .A2(new_n667), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT106), .Z(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n679), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G29gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n707), .A2(new_n708), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n709), .A2(new_n718), .A3(new_n719), .ZN(G1328gat));
  NOR2_X1   g519(.A1(new_n583), .A2(new_n287), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n644), .B2(new_n313), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n724), .A2(new_n582), .A3(new_n711), .A4(new_n716), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n722), .A2(KEYINPUT46), .B1(new_n287), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n722), .B2(KEYINPUT46), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n705), .A2(KEYINPUT107), .A3(new_n729), .A4(new_n721), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n726), .A2(new_n728), .A3(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT47), .ZN(new_n733));
  INV_X1    g532(.A(new_n640), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n724), .A2(new_n734), .A3(new_n711), .A4(new_n716), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n732), .A2(KEYINPUT47), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n669), .A2(new_n677), .ZN(new_n739));
  INV_X1    g538(.A(new_n704), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n693), .A2(G43gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  AND4_X1   g541(.A1(new_n733), .A2(new_n736), .A3(new_n738), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n737), .B1(new_n705), .B2(new_n741), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n733), .B1(new_n744), .B2(new_n736), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n745), .ZN(G1330gat));
  INV_X1    g545(.A(G50gat), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n724), .A2(new_n697), .A3(new_n711), .A4(new_n716), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(KEYINPUT109), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n714), .A2(new_n750), .A3(new_n697), .A4(new_n716), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n495), .A2(G50gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n705), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n705), .A2(new_n754), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n748), .A2(G50gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(G1331gat));
  INV_X1    g559(.A(new_n701), .ZN(new_n761));
  INV_X1    g560(.A(new_n247), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n761), .A2(new_n762), .A3(new_n667), .A4(new_n703), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n676), .A2(new_n679), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  OAI21_X1  g564(.A(new_n763), .B1(new_n710), .B2(new_n596), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n676), .A2(KEYINPUT110), .A3(new_n763), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n770), .A2(new_n583), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT111), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT49), .B(G64gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n768), .A2(new_n582), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n772), .B1(new_n771), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(G1333gat));
  AND2_X1   g576(.A1(new_n768), .A2(new_n769), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(G71gat), .A3(new_n734), .ZN(new_n779));
  INV_X1    g578(.A(G71gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n766), .B2(new_n693), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n779), .A2(KEYINPUT50), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT50), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n778), .A2(new_n697), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n247), .A2(new_n667), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n701), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n714), .A2(new_n679), .A3(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n703), .B(new_n787), .C1(new_n710), .C2(new_n596), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n676), .A2(KEYINPUT51), .A3(new_n703), .A4(new_n787), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n701), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n679), .A2(new_n253), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n789), .A2(new_n253), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  NOR3_X1   g596(.A1(new_n761), .A2(new_n583), .A3(G92gat), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n794), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n724), .A2(new_n582), .A3(new_n711), .A4(new_n788), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G92gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n798), .B(KEYINPUT112), .Z(new_n804));
  AOI22_X1  g603(.A1(G92gat), .A2(new_n800), .B1(new_n794), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(G1337gat));
  AND3_X1   g605(.A1(new_n714), .A2(new_n734), .A3(new_n788), .ZN(new_n807));
  INV_X1    g606(.A(G99gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n636), .A2(new_n808), .ZN(new_n809));
  OAI22_X1  g608(.A1(new_n807), .A2(new_n808), .B1(new_n795), .B2(new_n809), .ZN(G1338gat));
  NAND4_X1  g609(.A1(new_n724), .A2(new_n697), .A3(new_n711), .A4(new_n788), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(G106gat), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n495), .A2(G106gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n795), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n812), .B(new_n816), .C1(new_n795), .C2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n273), .A2(new_n819), .A3(new_n274), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n269), .B2(new_n270), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n265), .A2(new_n276), .A3(new_n268), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n820), .A2(KEYINPUT55), .A3(new_n314), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n316), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(new_n827), .A3(new_n316), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n820), .A2(new_n314), .A3(new_n823), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n826), .A2(new_n667), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n653), .A2(new_n654), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n648), .B1(new_n645), .B2(new_n647), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n661), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n701), .A2(new_n666), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n703), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n666), .A2(new_n835), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n313), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n826), .A2(new_n828), .A3(new_n839), .A4(new_n831), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n762), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n317), .A2(KEYINPUT113), .A3(new_n667), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT113), .B1(new_n317), .B2(new_n667), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n551), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n501), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n582), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(G113gat), .B1(new_n849), .B2(new_n667), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n697), .B1(new_n842), .B2(new_n845), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n551), .A2(new_n582), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(new_n636), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n668), .A2(new_n347), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(G1340gat));
  AOI21_X1  g654(.A(G120gat), .B1(new_n849), .B2(new_n701), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n761), .A2(new_n349), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1341gat));
  NAND2_X1  g657(.A1(new_n849), .A2(new_n247), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n353), .A2(new_n355), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n762), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n860), .A2(new_n862), .B1(new_n853), .B2(new_n863), .ZN(G1342gat));
  NAND2_X1  g663(.A1(new_n853), .A2(new_n703), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G134gat), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n313), .A2(G134gat), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT56), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n849), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n866), .A2(new_n869), .A3(new_n874), .A4(new_n871), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n852), .A2(new_n640), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n831), .A2(new_n667), .A3(new_n316), .A4(new_n824), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n836), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n313), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n247), .B1(new_n880), .B2(new_n840), .ZN(new_n881));
  INV_X1    g680(.A(new_n845), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n697), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n883), .B2(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n495), .B1(new_n842), .B2(new_n845), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(G141gat), .B1(new_n888), .B2(new_n668), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n640), .A2(new_n697), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n582), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n846), .A2(new_n891), .ZN(new_n892));
  OR3_X1    g691(.A1(new_n892), .A2(G141gat), .A3(new_n668), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n889), .B(new_n893), .C1(new_n896), .C2(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1344gat));
  NOR2_X1   g699(.A1(new_n495), .A2(KEYINPUT57), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n317), .A2(new_n667), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT118), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n901), .B1(new_n881), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n877), .A2(new_n761), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n904), .B(new_n905), .C1(new_n885), .C2(new_n886), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(G148gat), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT59), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(G148gat), .C1(new_n888), .C2(new_n761), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  OR3_X1    g712(.A1(new_n892), .A2(G148gat), .A3(new_n761), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n888), .B2(new_n762), .ZN(new_n916));
  INV_X1    g715(.A(new_n892), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n443), .A3(new_n247), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1346gat));
  NOR3_X1   g718(.A1(new_n888), .A2(new_n444), .A3(new_n313), .ZN(new_n920));
  AOI21_X1  g719(.A(G162gat), .B1(new_n917), .B2(new_n703), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1347gat));
  AOI21_X1  g721(.A(new_n679), .B1(new_n842), .B2(new_n845), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n847), .A2(new_n583), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(G169gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n667), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n679), .A2(new_n583), .A3(new_n693), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n851), .A2(new_n667), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT120), .A3(G169gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT120), .B1(new_n929), .B2(G169gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT121), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n934), .B(new_n927), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n925), .A2(new_n937), .A3(new_n701), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n851), .A2(new_n928), .ZN(new_n939));
  OAI21_X1  g738(.A(G176gat), .B1(new_n939), .B2(new_n761), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1349gat));
  AND2_X1   g740(.A1(new_n247), .A2(new_n377), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n924), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT122), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n923), .A2(new_n945), .A3(new_n924), .A4(new_n942), .ZN(new_n946));
  AOI22_X1  g745(.A1(new_n944), .A2(new_n946), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n948), .B1(new_n939), .B2(new_n762), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n851), .A2(KEYINPUT123), .A3(new_n247), .A4(new_n928), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(G183gat), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g750(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n947), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n952), .B1(new_n947), .B2(new_n951), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n939), .B2(new_n313), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n925), .A2(new_n325), .A3(new_n703), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1351gat));
  NOR2_X1   g758(.A1(new_n890), .A2(new_n583), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n923), .A2(new_n960), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n961), .A2(G197gat), .A3(new_n668), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT125), .Z(new_n963));
  NOR3_X1   g762(.A1(new_n734), .A2(new_n679), .A3(new_n583), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n904), .B(new_n964), .C1(new_n885), .C2(new_n886), .ZN(new_n965));
  OAI21_X1  g764(.A(G197gat), .B1(new_n965), .B2(new_n668), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n963), .A2(new_n966), .ZN(G1352gat));
  NOR3_X1   g766(.A1(new_n961), .A2(G204gat), .A3(new_n761), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT62), .ZN(new_n969));
  OAI21_X1  g768(.A(G204gat), .B1(new_n965), .B2(new_n761), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(G1353gat));
  INV_X1    g770(.A(new_n965), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(new_n247), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n974));
  OAI211_X1 g773(.A(KEYINPUT63), .B(G211gat), .C1(new_n965), .C2(new_n762), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n247), .A2(new_n430), .ZN(new_n977));
  OAI22_X1  g776(.A1(new_n974), .A2(new_n976), .B1(new_n961), .B2(new_n977), .ZN(G1354gat));
  NOR2_X1   g777(.A1(new_n313), .A2(new_n431), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n923), .A2(new_n703), .A3(new_n960), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n982));
  AND3_X1   g781(.A1(new_n981), .A2(new_n982), .A3(new_n431), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n982), .B1(new_n981), .B2(new_n431), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI211_X1 g786(.A(new_n980), .B(KEYINPUT127), .C1(new_n984), .C2(new_n983), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(G1355gat));
endmodule


