

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584;

  XNOR2_X1 U326 ( .A(n397), .B(n296), .ZN(n564) );
  NOR2_X1 U327 ( .A1(n583), .A2(n578), .ZN(n502) );
  NOR2_X1 U328 ( .A1(n497), .A2(n528), .ZN(n514) );
  AND2_X1 U329 ( .A1(n560), .A2(n559), .ZN(n565) );
  XOR2_X1 U330 ( .A(n479), .B(KEYINPUT41), .Z(n531) );
  INV_X1 U331 ( .A(n548), .ZN(n559) );
  NAND2_X1 U332 ( .A1(n543), .A2(n372), .ZN(n349) );
  XNOR2_X1 U333 ( .A(n513), .B(KEYINPUT48), .ZN(n541) );
  NAND2_X1 U334 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U335 ( .A(n510), .B(n509), .ZN(n511) );
  AND2_X1 U336 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U337 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n294) );
  XOR2_X1 U338 ( .A(KEYINPUT45), .B(n502), .Z(n295) );
  XOR2_X1 U339 ( .A(n396), .B(n395), .Z(n296) );
  XOR2_X1 U340 ( .A(n390), .B(n389), .Z(n297) );
  XOR2_X1 U341 ( .A(n584), .B(KEYINPUT62), .Z(n298) );
  XNOR2_X1 U342 ( .A(G36GAT), .B(G190GAT), .ZN(n338) );
  XNOR2_X1 U343 ( .A(KEYINPUT116), .B(KEYINPUT47), .ZN(n509) );
  XNOR2_X1 U344 ( .A(n338), .B(KEYINPUT79), .ZN(n386) );
  NOR2_X1 U345 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U346 ( .A(n564), .B(KEYINPUT103), .ZN(n462) );
  XNOR2_X1 U347 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U348 ( .A(n433), .B(n432), .ZN(n479) );
  XNOR2_X1 U349 ( .A(n570), .B(KEYINPUT125), .ZN(n582) );
  XOR2_X1 U350 ( .A(G211GAT), .B(KEYINPUT88), .Z(n300) );
  XNOR2_X1 U351 ( .A(KEYINPUT22), .B(KEYINPUT89), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n317) );
  XOR2_X1 U353 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n302) );
  NAND2_X1 U354 ( .A1(G228GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U356 ( .A(n303), .B(KEYINPUT23), .Z(n309) );
  XOR2_X1 U357 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n305) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(G162GAT), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n331) );
  XOR2_X1 U360 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n307) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(G218GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n345) );
  XNOR2_X1 U363 ( .A(n331), .B(n345), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U365 ( .A(G155GAT), .B(G204GAT), .Z(n311) );
  XOR2_X1 U366 ( .A(G50GAT), .B(KEYINPUT75), .Z(n385) );
  XOR2_X1 U367 ( .A(G106GAT), .B(G78GAT), .Z(n428) );
  XNOR2_X1 U368 ( .A(n385), .B(n428), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U370 ( .A(n313), .B(n312), .Z(n315) );
  XNOR2_X1 U371 ( .A(G22GAT), .B(G148GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U373 ( .A(n317), .B(n316), .Z(n546) );
  XOR2_X1 U374 ( .A(n546), .B(KEYINPUT28), .Z(n497) );
  XOR2_X1 U375 ( .A(KEYINPUT93), .B(KEYINPUT91), .Z(n319) );
  XNOR2_X1 U376 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n335) );
  XOR2_X1 U378 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n321) );
  XNOR2_X1 U379 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U381 ( .A(n322), .B(G57GAT), .Z(n324) );
  XOR2_X1 U382 ( .A(G120GAT), .B(G148GAT), .Z(n429) );
  XNOR2_X1 U383 ( .A(n429), .B(G85GAT), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n329) );
  XNOR2_X1 U385 ( .A(G1GAT), .B(G127GAT), .ZN(n325) );
  XNOR2_X1 U386 ( .A(n325), .B(G155GAT), .ZN(n400) );
  XOR2_X1 U387 ( .A(G113GAT), .B(KEYINPUT0), .Z(n353) );
  XOR2_X1 U388 ( .A(n400), .B(n353), .Z(n327) );
  NAND2_X1 U389 ( .A1(G225GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U390 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U391 ( .A(n329), .B(n328), .Z(n333) );
  XNOR2_X1 U392 ( .A(G29GAT), .B(G134GAT), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n330), .B(KEYINPUT78), .ZN(n393) );
  XNOR2_X1 U394 ( .A(n331), .B(n393), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U396 ( .A(n335), .B(n334), .Z(n376) );
  XNOR2_X1 U397 ( .A(KEYINPUT95), .B(n376), .ZN(n543) );
  XOR2_X1 U398 ( .A(G64GAT), .B(G92GAT), .Z(n337) );
  XNOR2_X1 U399 ( .A(G176GAT), .B(G204GAT), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n337), .B(n336), .ZN(n419) );
  XOR2_X1 U401 ( .A(KEYINPUT96), .B(n386), .Z(n340) );
  NAND2_X1 U402 ( .A1(G226GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U404 ( .A(G8GAT), .B(G183GAT), .Z(n341) );
  XOR2_X1 U405 ( .A(G211GAT), .B(n341), .Z(n399) );
  XOR2_X1 U406 ( .A(n342), .B(n399), .Z(n347) );
  XOR2_X1 U407 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n344) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n352), .B(n345), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n419), .B(n348), .ZN(n540) );
  XNOR2_X1 U413 ( .A(KEYINPUT27), .B(n540), .ZN(n372) );
  XOR2_X1 U414 ( .A(KEYINPUT97), .B(n349), .Z(n528) );
  XNOR2_X1 U415 ( .A(KEYINPUT98), .B(n514), .ZN(n367) );
  XOR2_X1 U416 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n351) );
  XNOR2_X1 U417 ( .A(G134GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n366) );
  XOR2_X1 U419 ( .A(n353), .B(n352), .Z(n355) );
  XNOR2_X1 U420 ( .A(G43GAT), .B(G99GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U422 ( .A(G71GAT), .B(G120GAT), .Z(n357) );
  NAND2_X1 U423 ( .A1(G227GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U425 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U426 ( .A(G127GAT), .B(G176GAT), .Z(n361) );
  XNOR2_X1 U427 ( .A(KEYINPUT85), .B(G183GAT), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U429 ( .A(G15GAT), .B(n362), .ZN(n363) );
  XNOR2_X1 U430 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n548) );
  NAND2_X1 U432 ( .A1(n367), .A2(n548), .ZN(n379) );
  NAND2_X1 U433 ( .A1(n540), .A2(n559), .ZN(n368) );
  NAND2_X1 U434 ( .A1(n368), .A2(n546), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n369), .B(KEYINPUT99), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n370), .B(KEYINPUT25), .ZN(n374) );
  NOR2_X1 U437 ( .A1(n546), .A2(n559), .ZN(n371) );
  XNOR2_X1 U438 ( .A(n371), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U439 ( .A1(n372), .A2(n568), .ZN(n373) );
  NAND2_X1 U440 ( .A1(n374), .A2(n373), .ZN(n375) );
  XNOR2_X1 U441 ( .A(KEYINPUT100), .B(n375), .ZN(n377) );
  NAND2_X1 U442 ( .A1(n377), .A2(n376), .ZN(n378) );
  NAND2_X1 U443 ( .A1(n379), .A2(n378), .ZN(n463) );
  XOR2_X1 U444 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n381) );
  XNOR2_X1 U445 ( .A(KEYINPUT76), .B(KEYINPUT11), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U447 ( .A(n382), .B(KEYINPUT77), .Z(n384) );
  XOR2_X1 U448 ( .A(G99GAT), .B(G85GAT), .Z(n427) );
  XNOR2_X1 U449 ( .A(G218GAT), .B(n427), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n390) );
  XOR2_X1 U451 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U452 ( .A1(G232GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U454 ( .A(G43GAT), .B(KEYINPUT7), .Z(n392) );
  XNOR2_X1 U455 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n440) );
  XNOR2_X1 U457 ( .A(n440), .B(n393), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n297), .B(n394), .ZN(n397) );
  XOR2_X1 U459 ( .A(KEYINPUT9), .B(G92GAT), .Z(n396) );
  XNOR2_X1 U460 ( .A(G162GAT), .B(G106GAT), .ZN(n395) );
  XNOR2_X1 U461 ( .A(G71GAT), .B(G57GAT), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n294), .B(n398), .ZN(n418) );
  XOR2_X1 U463 ( .A(n418), .B(n399), .Z(n413) );
  XOR2_X1 U464 ( .A(G64GAT), .B(n400), .Z(n402) );
  XOR2_X1 U465 ( .A(G15GAT), .B(G22GAT), .Z(n437) );
  XNOR2_X1 U466 ( .A(n437), .B(G78GAT), .ZN(n401) );
  XNOR2_X1 U467 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U468 ( .A(KEYINPUT83), .B(KEYINPUT15), .Z(n404) );
  NAND2_X1 U469 ( .A1(G231GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U470 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U471 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U472 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n408) );
  XNOR2_X1 U473 ( .A(KEYINPUT81), .B(KEYINPUT14), .ZN(n407) );
  XNOR2_X1 U474 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n409), .B(KEYINPUT82), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U477 ( .A(n413), .B(n412), .Z(n535) );
  INV_X1 U478 ( .A(n535), .ZN(n578) );
  NOR2_X1 U479 ( .A1(n564), .A2(n578), .ZN(n415) );
  XNOR2_X1 U480 ( .A(KEYINPUT16), .B(KEYINPUT84), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n416) );
  NAND2_X1 U482 ( .A1(n463), .A2(n416), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n417), .B(KEYINPUT101), .ZN(n480) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n424) );
  XOR2_X1 U485 ( .A(KEYINPUT32), .B(KEYINPUT73), .Z(n421) );
  NAND2_X1 U486 ( .A1(G230GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U487 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U488 ( .A(n422), .B(KEYINPUT31), .Z(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n426) );
  INV_X1 U490 ( .A(KEYINPUT33), .ZN(n425) );
  XNOR2_X1 U491 ( .A(n426), .B(n425), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n429), .B(KEYINPUT72), .ZN(n430) );
  XOR2_X1 U494 ( .A(G141GAT), .B(G113GAT), .Z(n435) );
  XNOR2_X1 U495 ( .A(G50GAT), .B(G29GAT), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U497 ( .A(n436), .B(G36GAT), .Z(n439) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n444) );
  XOR2_X1 U500 ( .A(n440), .B(KEYINPUT68), .Z(n442) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U503 ( .A(n444), .B(n443), .Z(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT30), .B(G1GAT), .Z(n446) );
  XNOR2_X1 U505 ( .A(G197GAT), .B(G8GAT), .ZN(n445) );
  XNOR2_X1 U506 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U507 ( .A(KEYINPUT70), .B(KEYINPUT66), .Z(n448) );
  XNOR2_X1 U508 ( .A(KEYINPUT29), .B(KEYINPUT67), .ZN(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U511 ( .A(n452), .B(n451), .Z(n529) );
  INV_X1 U512 ( .A(n529), .ZN(n571) );
  NOR2_X1 U513 ( .A1(n479), .A2(n571), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(KEYINPUT74), .ZN(n468) );
  AND2_X1 U515 ( .A1(n480), .A2(n468), .ZN(n459) );
  NAND2_X1 U516 ( .A1(n459), .A2(n543), .ZN(n454) );
  XNOR2_X1 U517 ( .A(KEYINPUT34), .B(n454), .ZN(n455) );
  XNOR2_X1 U518 ( .A(G1GAT), .B(n455), .ZN(G1324GAT) );
  NAND2_X1 U519 ( .A1(n540), .A2(n459), .ZN(n456) );
  XNOR2_X1 U520 ( .A(n456), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U521 ( .A(G15GAT), .B(KEYINPUT35), .Z(n458) );
  NAND2_X1 U522 ( .A1(n459), .A2(n559), .ZN(n457) );
  XNOR2_X1 U523 ( .A(n458), .B(n457), .ZN(G1326GAT) );
  NAND2_X1 U524 ( .A1(n459), .A2(n497), .ZN(n460) );
  XNOR2_X1 U525 ( .A(n460), .B(KEYINPUT102), .ZN(n461) );
  XNOR2_X1 U526 ( .A(G22GAT), .B(n461), .ZN(G1327GAT) );
  XOR2_X1 U527 ( .A(G29GAT), .B(KEYINPUT39), .Z(n471) );
  XNOR2_X1 U528 ( .A(n462), .B(KEYINPUT36), .ZN(n583) );
  NAND2_X1 U529 ( .A1(n578), .A2(n463), .ZN(n464) );
  XNOR2_X1 U530 ( .A(KEYINPUT104), .B(n464), .ZN(n465) );
  NOR2_X1 U531 ( .A1(n583), .A2(n465), .ZN(n467) );
  XNOR2_X1 U532 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n466) );
  XNOR2_X1 U533 ( .A(n467), .B(n466), .ZN(n491) );
  NAND2_X1 U534 ( .A1(n468), .A2(n491), .ZN(n469) );
  XOR2_X1 U535 ( .A(KEYINPUT38), .B(n469), .Z(n476) );
  NAND2_X1 U536 ( .A1(n476), .A2(n543), .ZN(n470) );
  XNOR2_X1 U537 ( .A(n471), .B(n470), .ZN(G1328GAT) );
  NAND2_X1 U538 ( .A1(n476), .A2(n540), .ZN(n472) );
  XNOR2_X1 U539 ( .A(n472), .B(KEYINPUT106), .ZN(n473) );
  XNOR2_X1 U540 ( .A(G36GAT), .B(n473), .ZN(G1329GAT) );
  NAND2_X1 U541 ( .A1(n476), .A2(n559), .ZN(n474) );
  XNOR2_X1 U542 ( .A(n474), .B(KEYINPUT40), .ZN(n475) );
  XNOR2_X1 U543 ( .A(G43GAT), .B(n475), .ZN(G1330GAT) );
  XOR2_X1 U544 ( .A(G50GAT), .B(KEYINPUT107), .Z(n478) );
  NAND2_X1 U545 ( .A1(n497), .A2(n476), .ZN(n477) );
  XNOR2_X1 U546 ( .A(n478), .B(n477), .ZN(G1331GAT) );
  INV_X1 U547 ( .A(n531), .ZN(n553) );
  NOR2_X1 U548 ( .A1(n529), .A2(n553), .ZN(n490) );
  NAND2_X1 U549 ( .A1(n490), .A2(n480), .ZN(n481) );
  XOR2_X1 U550 ( .A(KEYINPUT108), .B(n481), .Z(n487) );
  NAND2_X1 U551 ( .A1(n487), .A2(n543), .ZN(n482) );
  XNOR2_X1 U552 ( .A(n482), .B(KEYINPUT42), .ZN(n483) );
  XNOR2_X1 U553 ( .A(G57GAT), .B(n483), .ZN(G1332GAT) );
  XOR2_X1 U554 ( .A(G64GAT), .B(KEYINPUT109), .Z(n485) );
  NAND2_X1 U555 ( .A1(n487), .A2(n540), .ZN(n484) );
  XNOR2_X1 U556 ( .A(n485), .B(n484), .ZN(G1333GAT) );
  NAND2_X1 U557 ( .A1(n487), .A2(n559), .ZN(n486) );
  XNOR2_X1 U558 ( .A(n486), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U559 ( .A(G78GAT), .B(KEYINPUT43), .Z(n489) );
  NAND2_X1 U560 ( .A1(n497), .A2(n487), .ZN(n488) );
  XNOR2_X1 U561 ( .A(n489), .B(n488), .ZN(G1335GAT) );
  AND2_X1 U562 ( .A1(n491), .A2(n490), .ZN(n498) );
  NAND2_X1 U563 ( .A1(n543), .A2(n498), .ZN(n492) );
  XNOR2_X1 U564 ( .A(n492), .B(KEYINPUT110), .ZN(n493) );
  XNOR2_X1 U565 ( .A(G85GAT), .B(n493), .ZN(G1336GAT) );
  XOR2_X1 U566 ( .A(G92GAT), .B(KEYINPUT111), .Z(n495) );
  NAND2_X1 U567 ( .A1(n498), .A2(n540), .ZN(n494) );
  XNOR2_X1 U568 ( .A(n495), .B(n494), .ZN(G1337GAT) );
  NAND2_X1 U569 ( .A1(n498), .A2(n559), .ZN(n496) );
  XNOR2_X1 U570 ( .A(n496), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n500) );
  NAND2_X1 U572 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U573 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U574 ( .A(G106GAT), .B(n501), .Z(G1339GAT) );
  NOR2_X1 U575 ( .A1(n479), .A2(n295), .ZN(n503) );
  NAND2_X1 U576 ( .A1(n503), .A2(n571), .ZN(n512) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(n535), .Z(n561) );
  AND2_X1 U578 ( .A1(n529), .A2(n531), .ZN(n505) );
  XNOR2_X1 U579 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n504) );
  XNOR2_X1 U580 ( .A(n505), .B(n504), .ZN(n506) );
  NOR2_X1 U581 ( .A1(n561), .A2(n506), .ZN(n507) );
  XNOR2_X1 U582 ( .A(n507), .B(KEYINPUT115), .ZN(n508) );
  NOR2_X1 U583 ( .A1(n564), .A2(n508), .ZN(n510) );
  NAND2_X1 U584 ( .A1(n541), .A2(n514), .ZN(n515) );
  NOR2_X1 U585 ( .A1(n548), .A2(n515), .ZN(n516) );
  XOR2_X1 U586 ( .A(KEYINPUT117), .B(n516), .Z(n523) );
  NAND2_X1 U587 ( .A1(n529), .A2(n523), .ZN(n517) );
  XNOR2_X1 U588 ( .A(n517), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n519) );
  NAND2_X1 U590 ( .A1(n523), .A2(n531), .ZN(n518) );
  XNOR2_X1 U591 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U592 ( .A(G120GAT), .B(n520), .ZN(G1341GAT) );
  NAND2_X1 U593 ( .A1(n523), .A2(n561), .ZN(n521) );
  XNOR2_X1 U594 ( .A(n521), .B(KEYINPUT50), .ZN(n522) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n522), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n525) );
  NAND2_X1 U597 ( .A1(n523), .A2(n564), .ZN(n524) );
  XNOR2_X1 U598 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U599 ( .A(G134GAT), .B(n526), .Z(G1343GAT) );
  NAND2_X1 U600 ( .A1(n541), .A2(n568), .ZN(n527) );
  NOR2_X1 U601 ( .A1(n528), .A2(n527), .ZN(n538) );
  NAND2_X1 U602 ( .A1(n529), .A2(n538), .ZN(n530) );
  XNOR2_X1 U603 ( .A(n530), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n533) );
  NAND2_X1 U605 ( .A1(n538), .A2(n531), .ZN(n532) );
  XNOR2_X1 U606 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(n534), .ZN(G1345GAT) );
  XNOR2_X1 U608 ( .A(G155GAT), .B(KEYINPUT120), .ZN(n537) );
  NAND2_X1 U609 ( .A1(n535), .A2(n538), .ZN(n536) );
  XNOR2_X1 U610 ( .A(n537), .B(n536), .ZN(G1346GAT) );
  NAND2_X1 U611 ( .A1(n538), .A2(n564), .ZN(n539) );
  XNOR2_X1 U612 ( .A(n539), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U613 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U614 ( .A(n542), .B(KEYINPUT54), .ZN(n544) );
  XNOR2_X1 U615 ( .A(n545), .B(KEYINPUT64), .ZN(n569) );
  NAND2_X1 U616 ( .A1(n546), .A2(n569), .ZN(n547) );
  XNOR2_X2 U617 ( .A(n547), .B(KEYINPUT55), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n571), .A2(n548), .ZN(n549) );
  AND2_X1 U619 ( .A1(n560), .A2(n549), .ZN(n550) );
  XNOR2_X1 U620 ( .A(G169GAT), .B(n550), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n551), .B(KEYINPUT121), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n552) );
  NOR2_X1 U623 ( .A1(n553), .A2(n552), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n555) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U626 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U627 ( .A(KEYINPUT56), .B(n556), .ZN(n557) );
  XNOR2_X1 U628 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n565), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT124), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G190GAT), .ZN(G1351GAT) );
  NOR2_X1 U635 ( .A1(n571), .A2(n582), .ZN(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U640 ( .A(n582), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n575), .A2(n479), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  INV_X1 U643 ( .A(KEYINPUT126), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n578), .A2(n582), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n298), .ZN(G1355GAT) );
endmodule

