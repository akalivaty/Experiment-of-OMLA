//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1155;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT68), .B(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT70), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n464), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n468), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n467), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n477), .B(new_n480), .C1(G124), .C2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(new_n464), .A3(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT72), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n487), .A2(new_n464), .A3(G138), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n467), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n464), .C1(new_n484), .C2(new_n485), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n489), .A2(new_n492), .B1(KEYINPUT4), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OR2_X1    g070(.A1(KEYINPUT71), .A2(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT71), .A2(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n464), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n481), .A2(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n494), .A2(new_n500), .ZN(G164));
  OR2_X1    g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n509), .B2(new_n510), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n507), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G89), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(new_n513), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT74), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(new_n506), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n527), .B2(new_n508), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT73), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n524), .A2(new_n532), .ZN(G168));
  AND2_X1   g108(.A1(new_n529), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n535), .A2(new_n506), .B1(new_n536), .B2(new_n513), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n511), .A2(new_n512), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n502), .A2(new_n503), .B1(new_n527), .B2(new_n508), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(G81), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n529), .A2(G43), .B1(new_n543), .B2(KEYINPUT75), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT76), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n528), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT77), .B(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n540), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(G91), .B2(new_n545), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  OAI21_X1  g139(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT78), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n545), .A2(G87), .B1(new_n528), .B2(G49), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(G288));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  INV_X1    g144(.A(G48), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n513), .A2(new_n569), .B1(new_n515), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(G61), .B1(new_n511), .B2(new_n512), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n506), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AND2_X1   g151(.A1(new_n529), .A2(G47), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n578), .A2(new_n506), .B1(new_n579), .B2(new_n513), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G290));
  AOI22_X1  g157(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n506), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n545), .A2(G92), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(KEYINPUT10), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n529), .A2(G54), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n591), .B2(G171), .ZN(G284));
  OAI21_X1  g168(.A(new_n592), .B1(new_n591), .B2(G171), .ZN(G321));
  NAND2_X1  g169(.A1(G299), .A2(new_n591), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(G168), .B2(new_n591), .ZN(G297));
  OAI21_X1  g171(.A(new_n595), .B1(G168), .B2(new_n591), .ZN(G280));
  INV_X1    g172(.A(new_n590), .ZN(new_n598));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n547), .A2(new_n548), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(new_n591), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n590), .A2(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n591), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n467), .A2(new_n465), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n478), .A2(G135), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT79), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G111), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n612), .A2(new_n613), .B1(new_n615), .B2(G2105), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n482), .A2(G123), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT81), .Z(new_n619));
  INV_X1    g194(.A(G2096), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n609), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT82), .Z(G156));
  INV_X1    g199(.A(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT85), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n630), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n635), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n659), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n657), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n664), .B(new_n666), .C1(new_n657), .C2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  INV_X1    g248(.A(G29), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n674), .A2(G25), .ZN(new_n675));
  OAI21_X1  g250(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g252(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n678));
  OAI221_X1 g253(.A(G2104), .B1(G107), .B2(new_n464), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  AOI22_X1  g255(.A1(G119), .A2(new_n482), .B1(new_n478), .B2(G131), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n675), .B1(new_n682), .B2(new_n674), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT90), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT35), .B(G1991), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(KEYINPUT90), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n686), .B1(new_n684), .B2(new_n687), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G24), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n581), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1986), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n688), .A2(new_n689), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n690), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1971), .ZN(new_n697));
  NOR2_X1   g272(.A1(G6), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n575), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(G288), .A2(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n690), .A2(G23), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(new_n707), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n711), .ZN(new_n713));
  OAI21_X1  g288(.A(KEYINPUT93), .B1(new_n713), .B2(new_n708), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n715));
  NAND4_X1  g290(.A1(new_n702), .A2(new_n712), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n694), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT94), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n694), .A2(KEYINPUT94), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n702), .A2(new_n712), .A3(new_n714), .ZN(new_n722));
  INV_X1    g297(.A(new_n715), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT36), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n721), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n725), .B1(KEYINPUT95), .B2(KEYINPUT36), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n721), .A2(new_n728), .A3(new_n724), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT97), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI22_X1  g308(.A1(G129), .A2(new_n482), .B1(new_n478), .B2(G141), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT101), .B(KEYINPUT26), .Z(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n465), .A2(G105), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n734), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  MUX2_X1   g314(.A(G32), .B(new_n739), .S(G29), .Z(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT27), .B(G1996), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT102), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT103), .ZN(new_n744));
  INV_X1    g319(.A(G34), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(KEYINPUT24), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(KEYINPUT24), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n674), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G160), .B2(new_n674), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT100), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n744), .B1(G2084), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n690), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n690), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT104), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G168), .A2(new_n690), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n690), .B2(G21), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n752), .B(new_n757), .C1(G1966), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n598), .B2(G16), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n478), .A2(G140), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n482), .A2(G128), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n464), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G29), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n674), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n690), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n549), .B2(new_n690), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n775), .B1(G1341), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n765), .B(new_n778), .C1(G1341), .C2(new_n777), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n674), .A2(G35), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G162), .B2(new_n674), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT29), .B(G2090), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G164), .A2(new_n674), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G27), .B2(new_n674), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n785), .B1(new_n788), .B2(G2078), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n690), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n760), .B2(G1966), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n787), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT30), .B(G28), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n797), .A2(new_n674), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n618), .B2(new_n674), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n802));
  NAND2_X1  g377(.A1(G103), .A2(G2104), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n478), .A2(G139), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(new_n464), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G29), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G33), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT99), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n801), .B1(new_n815), .B2(G2072), .ZN(new_n816));
  INV_X1    g391(.A(G2072), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n742), .A2(new_n740), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G2084), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n816), .B(new_n818), .C1(new_n819), .C2(new_n750), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n789), .A2(new_n794), .A3(new_n796), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n761), .A2(new_n781), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n780), .B2(new_n779), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n733), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n732), .B1(new_n730), .B2(new_n731), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(G311));
  INV_X1    g401(.A(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n827), .A2(new_n733), .A3(new_n823), .ZN(G150));
  NAND2_X1  g403(.A1(new_n598), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n529), .A2(G55), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT105), .B(G93), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n832), .A2(new_n506), .B1(new_n513), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n549), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n831), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n601), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n830), .B(new_n839), .Z(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n835), .A2(new_n842), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  NAND2_X1  g422(.A1(new_n489), .A2(new_n492), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT106), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n494), .A2(KEYINPUT106), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n500), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n770), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n739), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n809), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n855), .A2(new_n739), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n739), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(new_n810), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n680), .A2(new_n681), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n607), .ZN(new_n863));
  OR2_X1    g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n864), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n865), .B1(new_n481), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(G142), .B2(new_n478), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n863), .B(new_n868), .Z(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n861), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n861), .A2(KEYINPUT107), .A3(new_n870), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT107), .B1(new_n861), .B2(new_n870), .ZN(new_n877));
  AOI211_X1 g452(.A(new_n872), .B(new_n869), .C1(new_n857), .C2(new_n860), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT108), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n861), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n869), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n876), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G162), .B(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n618), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n880), .B2(new_n869), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n877), .B2(new_n878), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n885), .A2(KEYINPUT40), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT40), .B1(new_n885), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(G395));
  NAND2_X1  g468(.A1(new_n837), .A2(new_n591), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n581), .B(G303), .ZN(new_n895));
  XNOR2_X1  g470(.A(G288), .B(new_n575), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n897), .A2(KEYINPUT42), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n897), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n900), .B2(KEYINPUT42), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n590), .B(G299), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n839), .B(new_n603), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n903), .B2(new_n908), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n901), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n894), .B1(new_n911), .B2(new_n591), .ZN(G295));
  OAI21_X1  g487(.A(new_n894), .B1(new_n911), .B2(new_n591), .ZN(G331));
  AOI21_X1  g488(.A(G301), .B1(new_n836), .B2(new_n838), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n836), .A2(new_n838), .A3(G301), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(G168), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G286), .B1(new_n918), .B2(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n903), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n904), .A2(new_n917), .A3(new_n919), .A4(new_n906), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n897), .B(KEYINPUT109), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(KEYINPUT110), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n900), .B1(new_n921), .B2(new_n922), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(G37), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT43), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n900), .A2(new_n921), .A3(new_n922), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n926), .A2(KEYINPUT43), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n926), .A2(KEYINPUT111), .A3(new_n935), .A4(new_n932), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n927), .B2(new_n930), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n934), .B1(new_n942), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g518(.A(G299), .B(KEYINPUT57), .Z(new_n944));
  XNOR2_X1  g519(.A(KEYINPUT118), .B(G1956), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n946));
  INV_X1    g521(.A(new_n500), .ZN(new_n947));
  AOI221_X4 g522(.A(new_n851), .B1(new_n493), .B2(KEYINPUT4), .C1(new_n489), .C2(new_n492), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT106), .B1(new_n848), .B2(new_n849), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(G160), .A2(G40), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n494), .B2(new_n500), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(KEYINPUT50), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n945), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n950), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n953), .B1(new_n959), .B2(new_n955), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(G2072), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n958), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n944), .B1(new_n957), .B2(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n957), .A2(new_n944), .A3(new_n963), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n590), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n946), .B1(new_n854), .B2(G1384), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n955), .A2(new_n946), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n953), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n950), .A2(new_n954), .A3(new_n951), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n970), .A2(G1348), .B1(G2067), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n964), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n958), .A2(new_n974), .A3(new_n960), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT58), .B(G1341), .Z(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n549), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT120), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT59), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n601), .B1(new_n975), .B2(new_n977), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT120), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n979), .A2(KEYINPUT120), .A3(new_n981), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT61), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n965), .B2(new_n964), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n957), .A2(new_n963), .ZN(new_n989));
  INV_X1    g564(.A(new_n944), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n957), .A2(new_n944), .A3(new_n963), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(KEYINPUT61), .A3(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n985), .A2(new_n986), .A3(new_n988), .A4(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n971), .A2(G2067), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT50), .B1(new_n950), .B2(new_n951), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n954), .B1(new_n996), .B2(new_n968), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n995), .B1(new_n997), .B2(new_n764), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(KEYINPUT60), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT60), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n598), .B1(new_n972), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(KEYINPUT60), .A3(new_n590), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n973), .B1(new_n994), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n1005));
  INV_X1    g580(.A(G8), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G168), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1007), .B2(KEYINPUT122), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n819), .B(new_n954), .C1(new_n996), .C2(new_n968), .ZN(new_n1010));
  INV_X1    g585(.A(G1966), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n950), .B2(new_n951), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n954), .B1(new_n955), .B2(new_n959), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1007), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1009), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1006), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1019), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT121), .ZN(new_n1021));
  AND4_X1   g596(.A1(new_n1021), .A2(new_n1015), .A3(G8), .A4(G286), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(new_n1019), .B2(G286), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1018), .A2(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT113), .B(G2090), .Z(new_n1026));
  NAND2_X1  g601(.A1(new_n954), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n967), .B2(new_n969), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1971), .B1(new_n958), .B2(new_n960), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1025), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n958), .A2(new_n960), .ZN(new_n1031));
  INV_X1    g606(.A(G1971), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n954), .B(new_n1026), .C1(new_n996), .C2(new_n968), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(KEYINPUT114), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G303), .A2(G8), .ZN(new_n1036));
  XNOR2_X1  g611(.A(new_n1036), .B(KEYINPUT55), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1030), .A2(new_n1035), .A3(G8), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1026), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n952), .A2(new_n956), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(G8), .B1(new_n1041), .B2(new_n1029), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1037), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n566), .A2(G1976), .A3(new_n567), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n971), .A2(G8), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1981), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n545), .A2(G86), .B1(new_n528), .B2(G48), .ZN(new_n1049));
  INV_X1    g624(.A(new_n574), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n571), .A2(new_n574), .A3(G1981), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT49), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1051), .A2(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1053), .B(new_n1054), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n971), .A2(new_n1057), .A3(G8), .A4(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT115), .B(G1976), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n971), .A2(new_n1044), .A3(G8), .A4(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1047), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1039), .A2(new_n1043), .A3(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(G171), .B(KEYINPUT54), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n997), .A2(new_n756), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT124), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1031), .B2(G2078), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n959), .B1(new_n854), .B2(G1384), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n953), .A2(new_n1069), .A3(G2078), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n958), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1067), .A2(KEYINPUT124), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1013), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(new_n1071), .A3(new_n795), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT123), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1077), .A2(new_n1071), .A3(new_n1080), .A4(new_n795), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(KEYINPUT53), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1066), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(new_n1067), .A3(new_n1070), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1065), .B1(new_n1076), .B2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1004), .A2(new_n1024), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1024), .A2(KEYINPUT62), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1016), .A2(new_n1017), .A3(new_n1009), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1008), .B1(new_n1019), .B2(new_n1007), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(new_n1091), .C1(new_n1023), .C2(new_n1022), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1082), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n1065), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1087), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(G288), .A2(G1976), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1059), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g673(.A(G8), .B(new_n971), .C1(new_n1098), .C2(new_n1052), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1047), .B2(new_n1063), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1046), .A2(KEYINPUT117), .A3(new_n1062), .A4(new_n1059), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1099), .B1(new_n1103), .B2(new_n1039), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1019), .A2(G168), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1065), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1030), .A2(new_n1035), .A3(G8), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1037), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1106), .A2(new_n1105), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1109), .A2(new_n1110), .A3(new_n1111), .A4(new_n1039), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1104), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1086), .A2(new_n1096), .A3(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1071), .A2(new_n953), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n770), .B(G2067), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT112), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n739), .B(new_n974), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n862), .A2(new_n686), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n682), .A2(new_n685), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n581), .B(G1986), .Z(new_n1122));
  OAI21_X1  g697(.A(new_n1115), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1114), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1115), .A2(new_n974), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT46), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT125), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1115), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n739), .B1(KEYINPUT46), .B2(new_n974), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1117), .A2(new_n1131), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1128), .A2(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT47), .ZN(new_n1134));
  OR3_X1    g709(.A1(new_n1130), .A2(G1986), .A3(G290), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(KEYINPUT48), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1121), .A2(new_n1115), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(KEYINPUT48), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1141), .A2(new_n1120), .B1(G2067), .B2(new_n770), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1115), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1134), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1124), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(KEYINPUT126), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1124), .A2(new_n1147), .A3(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g724(.A(new_n889), .B1(new_n882), .B2(new_n884), .ZN(new_n1151));
  NOR4_X1   g725(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1152));
  INV_X1    g726(.A(new_n1152), .ZN(new_n1153));
  NOR3_X1   g727(.A1(new_n942), .A2(new_n1151), .A3(new_n1153), .ZN(G308));
  NAND2_X1  g728(.A1(new_n885), .A2(new_n890), .ZN(new_n1155));
  OAI211_X1 g729(.A(new_n1155), .B(new_n1152), .C1(new_n941), .C2(new_n940), .ZN(G225));
endmodule


