//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(KEYINPUT16), .A3(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT95), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(G8gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n205), .B(new_n207), .C1(new_n204), .C2(new_n203), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(G8gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT96), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  INV_X1    g012(.A(G50gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT93), .A3(G43gat), .ZN(new_n215));
  XOR2_X1   g014(.A(G43gat), .B(G50gat), .Z(new_n216));
  OAI211_X1 g015(.A(new_n213), .B(new_n215), .C1(new_n216), .C2(KEYINPUT93), .ZN(new_n217));
  NOR2_X1   g016(.A1(G29gat), .A2(G36gat), .ZN(new_n218));
  XOR2_X1   g017(.A(new_n218), .B(KEYINPUT14), .Z(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT92), .B(G36gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G29gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n217), .A2(new_n219), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT94), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT91), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n223), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n219), .A2(new_n227), .ZN(new_n230));
  OAI211_X1 g029(.A(KEYINPUT15), .B(new_n220), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT97), .B1(new_n212), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n210), .B(KEYINPUT96), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT97), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(new_n231), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n210), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n240), .B1(new_n239), .B2(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n202), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n238), .B1(new_n234), .B2(new_n236), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n243), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n238), .A2(KEYINPUT18), .A3(new_n243), .A4(new_n241), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n245), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT90), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(G197gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT11), .B(G169gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(KEYINPUT12), .Z(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n256), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(KEYINPUT90), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G183gat), .B(G190gat), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT24), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n263));
  INV_X1    g062(.A(G169gat), .ZN(new_n264));
  INV_X1    g063(.A(G176gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT23), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT24), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(new_n265), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n264), .A2(new_n265), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT23), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n262), .A2(new_n268), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT25), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT27), .B(G183gat), .ZN(new_n278));
  INV_X1    g077(.A(G190gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n272), .B1(new_n273), .B2(KEYINPUT26), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n285), .A3(new_n267), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n278), .A2(new_n281), .A3(new_n279), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n283), .A2(new_n287), .A3(new_n269), .A4(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT25), .ZN(new_n290));
  OR2_X1    g089(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n291), .A2(KEYINPUT23), .A3(new_n265), .A4(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n275), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n270), .B1(new_n261), .B2(KEYINPUT24), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G127gat), .B(G134gat), .Z(new_n298));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n299), .A2(new_n300), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G120gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G113gat), .ZN(new_n307));
  XOR2_X1   g106(.A(KEYINPUT68), .B(G113gat), .Z(new_n308));
  OAI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(new_n306), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n298), .A2(KEYINPUT1), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G227gat), .ZN(new_n314));
  INV_X1    g113(.A(G233gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n276), .A2(KEYINPUT25), .B1(new_n294), .B2(new_n295), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n305), .A2(new_n311), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n289), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT32), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT33), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G15gat), .B(G43gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G71gat), .B(G99gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n323), .A3(new_n327), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT33), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n320), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n316), .B1(new_n313), .B2(new_n319), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT34), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI211_X1 g135(.A(KEYINPUT34), .B(new_n316), .C1(new_n313), .C2(new_n319), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n336), .A2(new_n337), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n328), .A3(new_n332), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(KEYINPUT70), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT70), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n333), .A2(new_n338), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT36), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT71), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n347), .A3(new_n341), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT36), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n340), .A2(new_n328), .A3(KEYINPUT71), .A4(new_n332), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G226gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(new_n315), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n297), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n354), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n357), .B1(new_n317), .B2(new_n289), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT72), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n362));
  OR2_X1    g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n361), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT74), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n297), .A2(new_n354), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n358), .A2(KEYINPUT73), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n356), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n368), .B(new_n372), .C1(new_n377), .C2(new_n367), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT30), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT76), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n356), .A2(new_n366), .A3(new_n358), .ZN(new_n381));
  INV_X1    g180(.A(new_n356), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n373), .A2(new_n374), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT73), .B1(new_n297), .B2(new_n354), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n381), .B1(new_n385), .B2(new_n366), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT30), .A4(new_n372), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n380), .A2(new_n388), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n372), .B(KEYINPUT75), .Z(new_n390));
  OAI21_X1  g189(.A(KEYINPUT30), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n378), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n394));
  INV_X1    g193(.A(G141gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(G148gat), .ZN(new_n396));
  INV_X1    g195(.A(G148gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G141gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT2), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G155gat), .B(G162gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(KEYINPUT78), .B(G155gat), .Z(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(G162gat), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n400), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n396), .A2(new_n398), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n395), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n402), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT80), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n407), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n396), .A2(new_n398), .A3(new_n408), .ZN(new_n414));
  INV_X1    g213(.A(G162gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G155gat), .ZN(new_n416));
  INV_X1    g215(.A(G155gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G162gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n410), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g219(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT78), .B(G155gat), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT2), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT80), .B1(new_n420), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n394), .B(new_n404), .C1(new_n413), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT82), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n412), .B1(new_n407), .B2(new_n411), .ZN(new_n429));
  INV_X1    g228(.A(new_n419), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n425), .A2(new_n430), .A3(KEYINPUT80), .A4(new_n409), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n429), .A2(new_n431), .B1(new_n403), .B2(new_n401), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n394), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n404), .B1(new_n413), .B2(new_n426), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(KEYINPUT81), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT3), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n440), .A3(new_n318), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n432), .A2(new_n312), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT4), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT5), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n438), .A2(new_n318), .A3(new_n439), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n443), .ZN(new_n448));
  INV_X1    g247(.A(new_n442), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n441), .A2(new_n444), .A3(new_n446), .A4(new_n442), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT0), .ZN(new_n455));
  XNOR2_X1  g254(.A(G57gat), .B(G85gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(new_n457), .A3(new_n452), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT83), .B(KEYINPUT6), .Z(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n457), .B1(new_n451), .B2(new_n452), .ZN(new_n463));
  INV_X1    g262(.A(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n393), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G78gat), .B(G106gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G50gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G22gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(new_n469), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n367), .B1(new_n435), .B2(new_n355), .ZN(new_n475));
  INV_X1    g274(.A(G228gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n315), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT3), .B1(new_n367), .B2(new_n355), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n438), .A2(new_n439), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n478), .A2(new_n432), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  OAI221_X1 g281(.A(new_n474), .B1(new_n475), .B2(new_n480), .C1(new_n482), .C2(new_n477), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n435), .A2(new_n355), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n366), .ZN(new_n485));
  INV_X1    g284(.A(new_n481), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n477), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n475), .A2(new_n480), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n473), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n352), .B1(new_n466), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT85), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT85), .B1(new_n389), .B2(new_n392), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n442), .B1(new_n441), .B2(new_n444), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT39), .B1(new_n448), .B2(new_n449), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT39), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n458), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n501), .B1(new_n500), .B2(new_n503), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n386), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n372), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n386), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT38), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n385), .A2(new_n367), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n512), .B1(new_n359), .B2(new_n366), .ZN(new_n516));
  AOI211_X1 g315(.A(KEYINPUT38), .B(new_n390), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n517), .A2(new_n509), .B1(new_n386), .B2(new_n372), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n518), .A3(new_n465), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n460), .A2(new_n461), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n496), .A2(new_n522), .A3(new_n497), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n490), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n492), .B1(new_n507), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n348), .A2(new_n350), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT35), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n491), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n495), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n465), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n490), .B1(new_n344), .B2(new_n342), .ZN(new_n531));
  INV_X1    g330(.A(new_n393), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n465), .B1(new_n521), .B2(new_n463), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n529), .A2(new_n530), .B1(KEYINPUT35), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT89), .B1(new_n525), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n349), .B1(new_n342), .B2(new_n344), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n533), .A2(new_n532), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n539), .B1(new_n490), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n494), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n389), .A2(new_n392), .A3(KEYINPUT85), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n496), .B(new_n497), .C1(new_n504), .C2(new_n505), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n548));
  NOR3_X1   g347(.A1(new_n547), .A2(new_n548), .A3(new_n521), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n491), .B1(new_n549), .B2(new_n519), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n541), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n552));
  INV_X1    g351(.A(new_n528), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n553), .A3(new_n544), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n534), .A2(KEYINPUT35), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n260), .B1(new_n536), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n533), .ZN(new_n559));
  NAND2_X1  g358(.A1(G85gat), .A2(G92gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(G92gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G99gat), .B(G106gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  AND2_X1   g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n236), .A2(new_n568), .B1(KEYINPUT41), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n232), .B2(KEYINPUT17), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n236), .A2(new_n239), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n577));
  XNOR2_X1  g376(.A(G134gat), .B(G162gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n583));
  INV_X1    g382(.A(G64gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(G57gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT100), .Z(new_n586));
  INV_X1    g385(.A(G57gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(G64gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT99), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  INV_X1    g391(.A(G71gat), .ZN(new_n593));
  INV_X1    g392(.A(G78gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n588), .A2(new_n585), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n597), .A2(new_n595), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n591), .B(KEYINPUT98), .ZN(new_n599));
  OAI22_X1  g398(.A1(new_n590), .A2(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n212), .B1(new_n583), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n583), .ZN(new_n602));
  XNOR2_X1  g401(.A(G127gat), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT101), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n605), .A2(new_n611), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n582), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n571), .A2(new_n600), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT103), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n619), .A3(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n600), .B(new_n568), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT102), .B(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(G230gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n315), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G120gat), .B(G148gat), .Z(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  OAI211_X1 g433(.A(new_n629), .B(new_n634), .C1(new_n628), .C2(new_n622), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n627), .B1(new_n621), .B2(new_n624), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n628), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n615), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n558), .A2(new_n559), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g442(.A1(new_n558), .A2(new_n641), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT16), .B(G8gat), .Z(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n495), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(G8gat), .B1(new_n644), .B2(new_n544), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  MUX2_X1   g448(.A(new_n647), .B(new_n649), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g449(.A(new_n526), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n644), .A2(G15gat), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(G15gat), .B1(new_n644), .B2(new_n352), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(G1326gat));
  OR3_X1    g453(.A1(new_n644), .A2(KEYINPUT106), .A3(new_n491), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT106), .B1(new_n644), .B2(new_n491), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  NOR2_X1   g458(.A1(new_n614), .A2(new_n640), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n582), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n558), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G29gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n559), .A2(new_n664), .ZN(new_n665));
  OR3_X1    g464(.A1(new_n663), .A2(KEYINPUT107), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT107), .B1(new_n663), .B2(new_n665), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(KEYINPUT45), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n260), .A2(new_n661), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n536), .A2(new_n557), .ZN(new_n671));
  INV_X1    g470(.A(new_n582), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n525), .A2(new_n535), .A3(KEYINPUT108), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT108), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n551), .B2(new_n556), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n669), .B1(new_n673), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n533), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT45), .B1(new_n666), .B2(new_n667), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n682), .A2(new_n683), .ZN(G1328gat));
  NOR3_X1   g483(.A1(new_n663), .A2(new_n222), .A3(new_n544), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n222), .B1(new_n680), .B2(new_n544), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1329gat));
  OAI21_X1  g487(.A(G43gat), .B1(new_n680), .B2(new_n352), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n663), .A2(G43gat), .A3(new_n651), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1330gat));
  OAI21_X1  g492(.A(G50gat), .B1(new_n680), .B2(new_n491), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n558), .A2(new_n214), .A3(new_n490), .A4(new_n662), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT48), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1331gat));
  NOR2_X1   g497(.A1(new_n674), .A2(new_n676), .ZN(new_n699));
  INV_X1    g498(.A(new_n260), .ZN(new_n700));
  INV_X1    g499(.A(new_n640), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n700), .A2(new_n615), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n533), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT110), .B(G57gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1332gat));
  OR2_X1    g505(.A1(new_n703), .A2(KEYINPUT111), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(KEYINPUT111), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n495), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT49), .B(G64gat), .Z(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n709), .B2(new_n711), .ZN(G1333gat));
  NAND4_X1  g511(.A1(new_n707), .A2(G71gat), .A3(new_n539), .A4(new_n708), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n593), .B1(new_n703), .B2(new_n651), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n713), .B2(new_n714), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1334gat));
  NAND3_X1  g517(.A1(new_n707), .A2(new_n490), .A3(new_n708), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g519(.A1(new_n673), .A2(new_n679), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n700), .A2(new_n614), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n640), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n721), .A2(new_n533), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n525), .A2(new_n535), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n672), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT51), .B1(new_n725), .B2(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n559), .A2(new_n563), .A3(new_n640), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n724), .A2(new_n563), .B1(new_n731), .B2(new_n732), .ZN(G1336gat));
  INV_X1    g532(.A(new_n723), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n495), .B(new_n734), .C1(new_n673), .C2(new_n679), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G92gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n544), .A2(new_n701), .A3(G92gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n736), .B(new_n737), .C1(new_n731), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n727), .B1(new_n741), .B2(KEYINPUT51), .ZN(new_n742));
  OAI211_X1 g541(.A(KEYINPUT113), .B(new_n728), .C1(new_n725), .C2(new_n726), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n736), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT114), .B1(new_n746), .B2(KEYINPUT52), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n744), .B1(new_n735), .B2(G92gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n748), .A2(new_n749), .A3(new_n737), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n740), .B1(new_n747), .B2(new_n750), .ZN(G1337gat));
  NOR3_X1   g550(.A1(new_n721), .A2(new_n352), .A3(new_n723), .ZN(new_n752));
  INV_X1    g551(.A(G99gat), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n651), .A2(new_n701), .A3(G99gat), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT115), .Z(new_n755));
  OAI22_X1  g554(.A1(new_n752), .A2(new_n753), .B1(new_n731), .B2(new_n755), .ZN(G1338gat));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n490), .B(new_n734), .C1(new_n673), .C2(new_n679), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G106gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n743), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n701), .A2(new_n491), .A3(G106gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n758), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n729), .A2(new_n730), .A3(new_n762), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n758), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(G106gat), .B2(new_n759), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n757), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n766), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n759), .A2(G106gat), .B1(new_n761), .B2(new_n762), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n770), .B(KEYINPUT116), .C1(new_n771), .C2(new_n758), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n768), .A2(new_n772), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n246), .A2(new_n247), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n243), .B1(new_n238), .B2(new_n241), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n774), .B(new_n255), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n233), .A2(new_n237), .B1(new_n212), .B2(new_n232), .ZN(new_n778));
  INV_X1    g577(.A(new_n247), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n242), .A2(new_n244), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n255), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT117), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n245), .A2(new_n248), .A3(new_n249), .A4(new_n258), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n777), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n621), .A2(new_n627), .A3(new_n624), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n629), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n634), .B1(new_n637), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n788), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n635), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n784), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n614), .B1(new_n794), .B2(new_n672), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n777), .A2(new_n782), .A3(new_n783), .A4(new_n640), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n582), .B(new_n796), .C1(new_n260), .C2(new_n793), .ZN(new_n797));
  AOI22_X1  g596(.A1(new_n795), .A2(new_n797), .B1(new_n260), .B2(new_n641), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n495), .A2(new_n533), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n651), .A2(new_n490), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(G113gat), .B1(new_n803), .B2(new_n260), .ZN(new_n804));
  INV_X1    g603(.A(new_n531), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n798), .A2(new_n805), .A3(new_n800), .ZN(new_n806));
  INV_X1    g605(.A(new_n308), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n806), .A2(new_n700), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n804), .A2(new_n808), .ZN(G1340gat));
  NOR3_X1   g608(.A1(new_n803), .A2(new_n306), .A3(new_n701), .ZN(new_n810));
  AOI21_X1  g609(.A(G120gat), .B1(new_n806), .B2(new_n640), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(new_n811), .ZN(G1341gat));
  INV_X1    g611(.A(new_n614), .ZN(new_n813));
  OAI21_X1  g612(.A(G127gat), .B1(new_n803), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(G127gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n806), .A2(new_n815), .A3(new_n614), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1342gat));
  INV_X1    g616(.A(G134gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n806), .A2(new_n818), .A3(new_n672), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n819), .A2(KEYINPUT56), .ZN(new_n820));
  OAI21_X1  g619(.A(G134gat), .B1(new_n803), .B2(new_n582), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(KEYINPUT56), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(G1343gat));
  NOR2_X1   g622(.A1(new_n800), .A2(new_n539), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n672), .B1(new_n784), .B2(new_n793), .ZN(new_n825));
  INV_X1    g624(.A(new_n259), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n258), .B1(new_n250), .B2(KEYINPUT90), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n826), .A2(new_n793), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n796), .A2(new_n582), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n825), .B(new_n813), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n641), .A2(new_n260), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(new_n832), .B2(new_n490), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  AOI211_X1 g633(.A(new_n834), .B(new_n491), .C1(new_n830), .C2(new_n831), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n700), .B(new_n824), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n824), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n834), .B1(new_n798), .B2(new_n491), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n832), .A2(KEYINPUT57), .A3(new_n490), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(KEYINPUT118), .A3(new_n700), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n838), .A2(new_n843), .A3(G141gat), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n539), .A2(new_n491), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n801), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n700), .A2(new_n395), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n844), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n836), .A2(G141gat), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n847), .A2(new_n848), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT58), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n395), .B1(new_n836), .B2(new_n837), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n849), .B1(new_n858), .B2(new_n843), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n845), .B1(new_n853), .B2(new_n854), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT119), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n857), .A2(new_n861), .ZN(G1344gat));
  AOI21_X1  g661(.A(new_n397), .B1(new_n842), .B2(new_n640), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT59), .ZN(new_n865));
  INV_X1    g664(.A(new_n847), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n397), .A3(new_n640), .ZN(new_n867));
  XOR2_X1   g666(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n868));
  OAI211_X1 g667(.A(new_n865), .B(new_n867), .C1(new_n863), .C2(new_n868), .ZN(G1345gat));
  NAND3_X1  g668(.A1(new_n866), .A2(new_n424), .A3(new_n614), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n842), .A2(new_n614), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n424), .ZN(G1346gat));
  NAND3_X1  g671(.A1(new_n866), .A2(new_n423), .A3(new_n672), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n842), .A2(new_n874), .A3(new_n672), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n406), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n842), .B2(new_n672), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n873), .B1(new_n876), .B2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n544), .A2(new_n559), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n798), .A2(new_n805), .A3(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n881), .A2(new_n700), .A3(new_n291), .A4(new_n292), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n832), .A2(new_n802), .A3(new_n879), .ZN(new_n883));
  OAI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n260), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1348gat));
  INV_X1    g684(.A(new_n883), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(G176gat), .A3(new_n640), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n887), .A2(KEYINPUT122), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n887), .A2(KEYINPUT122), .ZN(new_n889));
  AOI21_X1  g688(.A(G176gat), .B1(new_n881), .B2(new_n640), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(G1349gat));
  NAND3_X1  g690(.A1(new_n881), .A2(new_n278), .A3(new_n614), .ZN(new_n892));
  OAI21_X1  g691(.A(G183gat), .B1(new_n883), .B2(new_n813), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n894));
  AOI22_X1  g693(.A1(new_n892), .A2(new_n893), .B1(KEYINPUT123), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(KEYINPUT123), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n895), .B(new_n896), .ZN(G1350gat));
  NAND2_X1  g696(.A1(new_n886), .A2(new_n672), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G190gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT124), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n901), .A3(G190gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n881), .A2(new_n279), .A3(new_n672), .ZN(new_n906));
  XNOR2_X1  g705(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n905), .B(new_n906), .C1(new_n903), .C2(new_n907), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n840), .A2(new_n841), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n880), .A2(new_n539), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(G197gat), .A3(new_n700), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n832), .A2(new_n490), .A3(new_n910), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT126), .ZN(new_n915));
  AOI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n700), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n913), .A2(new_n916), .ZN(G1352gat));
  NOR3_X1   g716(.A1(new_n914), .A2(G204gat), .A3(new_n701), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(KEYINPUT127), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(KEYINPUT127), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n920), .B(new_n921), .Z(new_n922));
  OAI21_X1  g721(.A(G204gat), .B1(new_n911), .B2(new_n701), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1353gat));
  INV_X1    g723(.A(G211gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n915), .A2(new_n925), .A3(new_n614), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n912), .A2(new_n614), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1354gat));
  INV_X1    g729(.A(G218gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n931), .A3(new_n672), .ZN(new_n932));
  OAI21_X1  g731(.A(G218gat), .B1(new_n911), .B2(new_n582), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1355gat));
endmodule


