//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  NAND2_X1  g000(.A1(KEYINPUT0), .A2(G128), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT0), .B(G128), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n189), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n202), .A2(new_n205), .A3(new_n208), .A4(new_n203), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(KEYINPUT66), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n206), .A2(new_n211), .A3(G131), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n210), .A2(KEYINPUT67), .A3(new_n212), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n199), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n192), .B(G146), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G128), .ZN(new_n221));
  OAI221_X1 g035(.A(new_n219), .B1(G128), .B2(new_n191), .C1(new_n194), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n203), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n201), .A2(G137), .ZN(new_n224));
  OAI21_X1  g038(.A(G131), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(new_n209), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n217), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G116), .ZN(new_n230));
  INV_X1    g044(.A(G116), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G119), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n210), .A2(KEYINPUT67), .A3(new_n212), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT67), .B1(new_n210), .B2(new_n212), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n198), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n226), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n228), .A2(new_n238), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT28), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n215), .A2(new_n216), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n227), .B1(new_n247), .B2(new_n198), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(new_n238), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n217), .A2(new_n237), .A3(new_n227), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT28), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(G101), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G210), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n253), .B(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n246), .A2(new_n251), .A3(KEYINPUT29), .A4(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT72), .B(G902), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(KEYINPUT73), .A3(new_n259), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n198), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n213), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n227), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n237), .B1(new_n267), .B2(KEYINPUT30), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n241), .A2(KEYINPUT30), .A3(new_n226), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n241), .A2(new_n271), .A3(KEYINPUT30), .A4(new_n226), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n273), .A2(new_n250), .A3(new_n256), .ZN(new_n274));
  INV_X1    g088(.A(new_n256), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n267), .A2(new_n238), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT28), .B1(new_n250), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n275), .B1(new_n246), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n262), .B(new_n263), .C1(KEYINPUT29), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G472), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n283));
  INV_X1    g097(.A(new_n268), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n271), .B1(new_n248), .B2(KEYINPUT30), .ZN(new_n285));
  INV_X1    g099(.A(new_n272), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n248), .A2(new_n238), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n256), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT31), .B1(new_n273), .B2(new_n290), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n256), .B1(new_n246), .B2(new_n277), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n283), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n295), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT70), .A3(new_n292), .A4(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G472), .A2(G902), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n300), .B(KEYINPUT71), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n282), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(KEYINPUT32), .B(new_n301), .C1(new_n296), .C2(new_n298), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n281), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n198), .A2(G125), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n222), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G953), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G224), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(G224), .A3(new_n313), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT7), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n312), .A2(new_n317), .A3(new_n314), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G104), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(new_n322), .B2(G107), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n324));
  INV_X1    g138(.A(G107), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G104), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n322), .A2(G107), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G101), .ZN(new_n329));
  INV_X1    g143(.A(G101), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n323), .A2(new_n326), .A3(new_n330), .A4(new_n327), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(KEYINPUT4), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n328), .A2(new_n333), .A3(G101), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n237), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n327), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n322), .A2(G107), .ZN(new_n337));
  OAI21_X1  g151(.A(G101), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n331), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n230), .A2(new_n232), .A3(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(G113), .B1(new_n230), .B2(KEYINPUT5), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n235), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n335), .B1(new_n339), .B2(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(G110), .B(G122), .Z(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n342), .B(KEYINPUT83), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(KEYINPUT82), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n340), .A2(KEYINPUT82), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n235), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT84), .ZN(new_n352));
  INV_X1    g166(.A(new_n339), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n354), .A3(new_n235), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n345), .A2(KEYINPUT8), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n345), .A2(KEYINPUT8), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n358), .B(new_n359), .C1(new_n343), .C2(new_n353), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n346), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(G902), .B1(new_n321), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n315), .A2(new_n316), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n344), .A2(new_n345), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT6), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n366), .B(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n346), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n365), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n307), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n371), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n363), .A3(new_n306), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G214), .B1(G237), .B2(G902), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n376), .B(KEYINPUT80), .Z(new_n377));
  NOR2_X1   g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(G110), .B(G140), .ZN(new_n380));
  INV_X1    g194(.A(G227), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G953), .ZN(new_n382));
  XOR2_X1   g196(.A(new_n380), .B(new_n382), .Z(new_n383));
  XNOR2_X1  g197(.A(new_n353), .B(new_n222), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT12), .B1(new_n247), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n384), .A2(KEYINPUT12), .A3(new_n266), .ZN(new_n386));
  OR2_X1    g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n353), .A2(new_n222), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n353), .A2(new_n222), .A3(KEYINPUT10), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n332), .A2(new_n198), .A3(new_n334), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n247), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n383), .B1(new_n387), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n383), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n393), .A2(new_n394), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G469), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n393), .A2(new_n394), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(new_n398), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n385), .A2(new_n386), .ZN(new_n404));
  OAI22_X1  g218(.A1(new_n403), .A2(new_n383), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G469), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n259), .ZN(new_n407));
  NAND2_X1  g221(.A1(G469), .A2(G902), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT9), .B(G234), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G221), .B1(new_n411), .B2(G902), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G475), .ZN(new_n414));
  INV_X1    g228(.A(G902), .ZN(new_n415));
  INV_X1    g229(.A(G140), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G125), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n309), .A2(G140), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT76), .A4(KEYINPUT16), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT16), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n417), .B2(KEYINPUT16), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n190), .B(new_n419), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n420), .B(new_n422), .C1(KEYINPUT16), .C2(new_n417), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n190), .B1(new_n426), .B2(new_n419), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT89), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G146), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT89), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n254), .A2(G214), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n434), .A2(G143), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(G131), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT17), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n254), .A2(G214), .B1(new_n434), .B2(G143), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n436), .B(new_n208), .C1(new_n435), .C2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n428), .A2(new_n432), .A3(new_n442), .A4(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT18), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n436), .B(new_n448), .C1(new_n435), .C2(new_n444), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT87), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n449), .A3(KEYINPUT87), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT77), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n417), .A2(new_n418), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n455), .B1(new_n417), .B2(new_n418), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n190), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n417), .A2(new_n418), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n459), .B(new_n460), .C1(new_n190), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(KEYINPUT77), .ZN(new_n464));
  AOI21_X1  g278(.A(G146), .B1(new_n464), .B2(new_n456), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n462), .A2(new_n190), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT86), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n441), .A2(KEYINPUT18), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n454), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G113), .B(G122), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(new_n322), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n447), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n427), .B1(new_n440), .B2(new_n445), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT19), .ZN(new_n475));
  OR3_X1    g289(.A1(new_n462), .A2(KEYINPUT88), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT88), .B1(new_n462), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n457), .B2(new_n458), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n476), .A2(new_n190), .A3(new_n477), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n472), .B1(new_n470), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n414), .B(new_n415), .C1(new_n473), .C2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n472), .B1(new_n447), .B2(new_n470), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n415), .B1(new_n473), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G475), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n447), .A2(new_n470), .A3(new_n472), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n463), .A2(new_n467), .B1(new_n441), .B2(KEYINPUT18), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n489), .A2(new_n454), .B1(new_n474), .B2(new_n479), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n488), .B1(new_n472), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n491), .A2(KEYINPUT20), .A3(new_n414), .A4(new_n415), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n484), .A2(new_n487), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n410), .A2(G217), .A3(new_n313), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n231), .A2(G122), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT14), .ZN(new_n496));
  INV_X1    g310(.A(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G116), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n497), .A2(G116), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n496), .A2(KEYINPUT91), .A3(new_n498), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G107), .ZN(new_n507));
  XNOR2_X1  g321(.A(G128), .B(G143), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n201), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n495), .A2(new_n498), .A3(new_n325), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(KEYINPUT13), .ZN(new_n512));
  OR3_X1    g326(.A1(new_n218), .A2(KEYINPUT13), .A3(G143), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(G134), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT90), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n495), .A2(new_n498), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G107), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n517), .A2(new_n510), .B1(new_n201), .B2(new_n508), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n512), .A2(new_n519), .A3(new_n513), .A4(G134), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n515), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n494), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n524));
  INV_X1    g338(.A(new_n494), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n521), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(KEYINPUT92), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n528), .B(new_n494), .C1(new_n511), .C2(new_n522), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n259), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT15), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n530), .B(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n493), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G952), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n535), .A2(KEYINPUT93), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(KEYINPUT93), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n313), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(G234), .B2(G237), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n313), .B(new_n259), .C1(G234), .C2(G237), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT21), .B(G898), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT94), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n534), .A2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n379), .A2(new_n413), .A3(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G110), .Z(new_n547));
  NAND2_X1  g361(.A1(new_n229), .A2(G128), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n229), .A2(KEYINPUT74), .A3(G128), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n550), .A2(new_n551), .B1(G119), .B2(new_n218), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n553), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n547), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT23), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(G119), .B2(new_n218), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n229), .A2(KEYINPUT23), .A3(G128), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n548), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(G110), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n430), .A4(new_n459), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n555), .A2(new_n556), .A3(new_n547), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(G110), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n565), .B(new_n566), .C1(new_n427), .C2(new_n425), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n430), .B(new_n459), .C1(new_n557), .C2(new_n562), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(new_n567), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n313), .A2(G221), .A3(G234), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT22), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G137), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n564), .A2(new_n567), .A3(new_n570), .A4(new_n574), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n259), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT25), .ZN(new_n579));
  INV_X1    g393(.A(G217), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n259), .B2(G234), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n576), .A2(new_n582), .A3(new_n259), .A4(new_n577), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n576), .A2(new_n577), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n581), .A2(G902), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n586), .B(KEYINPUT79), .Z(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n305), .A2(new_n546), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT95), .B(G101), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G3));
  NAND2_X1  g407(.A1(new_n299), .A2(new_n302), .ZN(new_n594));
  INV_X1    g408(.A(G472), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n258), .B1(new_n296), .B2(new_n298), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n378), .A2(new_n544), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n413), .A2(new_n589), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n493), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n527), .A2(new_n603), .A3(new_n529), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n523), .A2(KEYINPUT33), .A3(new_n526), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n604), .A2(G478), .A3(new_n259), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n530), .A2(new_n531), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n602), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n601), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT34), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND2_X1  g427(.A1(new_n602), .A2(new_n533), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n601), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  INV_X1    g433(.A(new_n597), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n575), .A2(KEYINPUT36), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n571), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n571), .A2(new_n621), .ZN(new_n623));
  AND2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n587), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n622), .A2(new_n587), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT98), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n626), .A2(new_n584), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n620), .A2(new_n546), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT37), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(G110), .Z(G12));
  NOR2_X1   g446(.A1(new_n379), .A2(new_n413), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT99), .B(G900), .Z(new_n634));
  NAND2_X1  g448(.A1(new_n540), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n539), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n614), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n305), .A2(new_n633), .A3(new_n629), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  INV_X1    g455(.A(new_n413), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n637), .B(KEYINPUT39), .Z(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT40), .Z(new_n646));
  NAND2_X1  g460(.A1(new_n372), .A2(new_n374), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT38), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n249), .A2(new_n250), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n415), .B1(new_n651), .B2(new_n256), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n275), .B1(new_n287), .B2(new_n289), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n654), .B1(new_n303), .B2(new_n304), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OR2_X1    g470(.A1(new_n656), .A2(KEYINPUT100), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(KEYINPUT100), .ZN(new_n658));
  INV_X1    g472(.A(new_n629), .ZN(new_n659));
  INV_X1    g473(.A(new_n377), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n493), .A2(new_n533), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT101), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n649), .A2(new_n657), .A3(new_n658), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G143), .ZN(G45));
  NAND2_X1  g479(.A1(new_n609), .A2(new_n637), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n305), .A2(new_n633), .A3(new_n629), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G146), .ZN(G48));
  NOR2_X1   g483(.A1(new_n598), .A2(new_n610), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n405), .A2(new_n259), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G469), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n412), .A3(new_n407), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n305), .A2(new_n590), .A3(new_n670), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  AND2_X1   g495(.A1(new_n305), .A2(new_n590), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n598), .A2(new_n614), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n682), .A2(new_n683), .A3(new_n678), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n305), .A2(new_n590), .A3(new_n684), .A4(new_n678), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT103), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT104), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n231), .ZN(G18));
  NOR3_X1   g504(.A1(new_n379), .A2(new_n545), .A3(new_n673), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n305), .A2(new_n691), .A3(new_n629), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT105), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  NAND2_X1  g508(.A1(new_n299), .A2(new_n259), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n256), .B1(new_n246), .B2(new_n251), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n294), .A2(new_n696), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n695), .A2(G472), .B1(new_n302), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n543), .B1(new_n675), .B2(new_n677), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n589), .B(KEYINPUT106), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n661), .A2(new_n647), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(KEYINPUT107), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n661), .A2(new_n703), .A3(new_n647), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND2_X1  g521(.A1(new_n697), .A2(new_n302), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n629), .B(new_n708), .C1(new_n596), .C2(new_n595), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n666), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n379), .A2(new_n673), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G125), .ZN(G27));
  NOR2_X1   g527(.A1(new_n647), .A2(new_n377), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n413), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n305), .A2(new_n590), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n305), .A2(new_n700), .A3(new_n667), .A4(new_n716), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n717), .A2(new_n718), .B1(new_n719), .B2(KEYINPUT42), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G131), .ZN(G33));
  NAND4_X1  g535(.A1(new_n305), .A2(new_n590), .A3(new_n639), .A4(new_n716), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G134), .ZN(G36));
  INV_X1    g537(.A(new_n412), .ZN(new_n724));
  INV_X1    g538(.A(new_n407), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n400), .A2(KEYINPUT45), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n396), .B2(new_n399), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(G469), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n408), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT46), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n725), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n408), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n724), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n734), .A2(new_n735), .A3(new_n644), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n735), .B1(new_n734), .B2(new_n644), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n608), .A2(new_n493), .A3(KEYINPUT43), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n493), .A2(KEYINPUT109), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n606), .A2(new_n607), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n484), .A2(new_n487), .A3(new_n743), .A4(new_n492), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n740), .B1(new_n745), .B2(KEYINPUT43), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n659), .B1(new_n746), .B2(KEYINPUT110), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n597), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(KEYINPUT43), .ZN(new_n750));
  INV_X1    g564(.A(new_n740), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT44), .A4(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n747), .A2(new_n754), .A3(new_n597), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT111), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n715), .B1(new_n756), .B2(new_n757), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n755), .A2(new_n758), .A3(new_n759), .A4(KEYINPUT112), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n739), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT113), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  XOR2_X1   g580(.A(new_n734), .B(KEYINPUT47), .Z(new_n767));
  NAND2_X1  g581(.A1(new_n714), .A2(new_n589), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n767), .A2(new_n305), .A3(new_n666), .A4(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n416), .ZN(G42));
  NAND2_X1  g584(.A1(new_n657), .A2(new_n658), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n672), .A2(new_n407), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(KEYINPUT49), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n660), .B1(new_n772), .B2(KEYINPUT49), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n648), .A2(new_n773), .A3(new_n774), .A4(new_n745), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n771), .A2(new_n412), .A3(new_n700), .A4(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n640), .A2(new_n668), .A3(new_n712), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n626), .A2(new_n584), .A3(new_n628), .A4(new_n637), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n702), .B2(new_n704), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n655), .A2(new_n642), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT118), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n655), .A2(new_n779), .A3(new_n782), .A4(new_n642), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n777), .A2(new_n784), .A3(KEYINPUT52), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(new_n777), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n609), .A2(KEYINPUT114), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n609), .A2(KEYINPUT114), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n614), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n599), .A2(new_n600), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n591), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n792), .B1(new_n685), .B2(new_n687), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n305), .A2(new_n590), .A3(new_n716), .A4(new_n718), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n714), .A2(new_n534), .A3(new_n637), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n797));
  OR2_X1    g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n413), .B1(new_n796), .B2(new_n797), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n305), .A2(new_n798), .A3(new_n629), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n794), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  AND4_X1   g615(.A1(new_n630), .A2(new_n679), .A3(new_n706), .A4(new_n692), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n698), .A2(new_n629), .A3(new_n667), .A4(new_n716), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n710), .A2(KEYINPUT116), .A3(new_n716), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n805), .A2(new_n722), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n793), .A2(new_n801), .A3(new_n802), .A4(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT53), .B1(new_n787), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n792), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n688), .A2(new_n810), .A3(new_n802), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n807), .A2(new_n720), .A3(new_n800), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n781), .A2(new_n783), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n640), .A2(new_n668), .A3(new_n712), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n777), .A2(new_n784), .A3(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT53), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n813), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT54), .B1(new_n809), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(KEYINPUT117), .A3(new_n820), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n809), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n813), .A2(new_n819), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n825), .B2(new_n823), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n826), .B2(KEYINPUT54), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n752), .A2(new_n636), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n698), .A2(new_n700), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n648), .A2(new_n660), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n831), .A2(new_n674), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n709), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n715), .A2(new_n673), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n829), .A2(new_n836), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n833), .A2(KEYINPUT50), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n636), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n771), .A2(new_n590), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n602), .A2(new_n608), .ZN(new_n841));
  OAI221_X1 g655(.A(new_n838), .B1(KEYINPUT50), .B2(new_n833), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n831), .A2(new_n714), .ZN(new_n843));
  INV_X1    g657(.A(new_n772), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n724), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT119), .Z(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n767), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(KEYINPUT51), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n767), .B2(new_n845), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n842), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n538), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n840), .B2(new_n610), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n305), .A2(new_n700), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n837), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n857));
  XOR2_X1   g671(.A(new_n856), .B(new_n857), .Z(new_n858));
  NOR4_X1   g672(.A1(new_n849), .A2(new_n852), .A3(new_n854), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n831), .A2(new_n711), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n827), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(G952), .A2(G953), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n776), .B1(new_n861), .B2(new_n862), .ZN(G75));
  NAND4_X1  g677(.A1(new_n809), .A2(new_n821), .A3(new_n258), .A4(new_n307), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT55), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n369), .A2(new_n370), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(new_n365), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT121), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(new_n872), .A3(new_n865), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n867), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n867), .B2(new_n873), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n313), .A2(G952), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G51));
  INV_X1    g691(.A(new_n822), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n809), .A2(new_n821), .A3(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n809), .A2(new_n821), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(KEYINPUT122), .A3(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n408), .B(KEYINPUT57), .Z(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n405), .ZN(new_n887));
  OR3_X1    g701(.A1(new_n882), .A2(new_n259), .A3(new_n729), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n876), .B1(new_n887), .B2(new_n888), .ZN(G54));
  NAND4_X1  g703(.A1(new_n809), .A2(new_n821), .A3(KEYINPUT58), .A4(new_n258), .ZN(new_n890));
  INV_X1    g704(.A(new_n491), .ZN(new_n891));
  OR3_X1    g705(.A1(new_n890), .A2(new_n414), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n876), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n890), .B2(new_n414), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G60));
  NAND2_X1  g709(.A1(new_n604), .A2(new_n605), .ZN(new_n896));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n827), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n896), .ZN(new_n900));
  INV_X1    g714(.A(new_n898), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n881), .A2(new_n884), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n899), .A2(new_n893), .A3(new_n902), .ZN(G63));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT60), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n809), .A2(new_n821), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT123), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n809), .A2(new_n821), .A3(KEYINPUT123), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n624), .ZN(new_n911));
  INV_X1    g725(.A(new_n585), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n893), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n911), .A2(KEYINPUT61), .A3(new_n893), .A4(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(G66));
  NAND2_X1  g732(.A1(new_n811), .A2(new_n313), .ZN(new_n919));
  INV_X1    g733(.A(G224), .ZN(new_n920));
  OAI21_X1  g734(.A(G953), .B1(new_n542), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n369), .B(new_n370), .C1(G898), .C2(new_n313), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G69));
  INV_X1    g738(.A(G900), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(G953), .ZN(new_n926));
  INV_X1    g740(.A(new_n720), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n738), .A2(new_n705), .A3(new_n855), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n777), .A3(new_n722), .ZN(new_n929));
  NOR4_X1   g743(.A1(new_n764), .A2(new_n927), .A3(new_n929), .A4(new_n769), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n926), .B1(new_n930), .B2(G953), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT125), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n285), .A2(new_n286), .B1(KEYINPUT30), .B2(new_n267), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n936), .B(new_n926), .C1(new_n930), .C2(G953), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n381), .B2(new_n925), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n764), .A2(new_n769), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n717), .A2(new_n644), .A3(new_n790), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT62), .B1(new_n664), .B2(new_n777), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n664), .A2(KEYINPUT62), .A3(new_n777), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n943), .B(new_n944), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n313), .ZN(new_n948));
  INV_X1    g762(.A(new_n935), .ZN(new_n949));
  AOI22_X1  g763(.A1(new_n948), .A2(new_n949), .B1(new_n941), .B2(new_n940), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n938), .A2(new_n942), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n942), .B1(new_n938), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(G72));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n947), .B2(new_n811), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n653), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n930), .A2(new_n793), .A3(new_n802), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n955), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n274), .B(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n653), .A2(new_n274), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n826), .A2(new_n955), .A3(new_n962), .ZN(new_n963));
  AND4_X1   g777(.A1(new_n893), .A2(new_n957), .A3(new_n961), .A4(new_n963), .ZN(G57));
endmodule


