

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n338, n339, n340, n341, n342, n343, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747;

  NOR2_X1 U360 ( .A1(n626), .A2(n715), .ZN(n627) );
  NOR2_X1 U361 ( .A1(n632), .A2(n715), .ZN(n635) );
  NOR2_X1 U362 ( .A1(n562), .A2(n395), .ZN(n370) );
  XNOR2_X1 U363 ( .A(n510), .B(n509), .ZN(n686) );
  INV_X1 U364 ( .A(n489), .ZN(n340) );
  XNOR2_X1 U365 ( .A(n339), .B(n338), .ZN(n502) );
  XNOR2_X1 U366 ( .A(n482), .B(n392), .ZN(n732) );
  XNOR2_X1 U367 ( .A(n500), .B(n501), .ZN(n338) );
  INV_X1 U368 ( .A(n372), .ZN(n339) );
  BUF_X1 U369 ( .A(G143), .Z(n342) );
  XNOR2_X1 U370 ( .A(G134), .B(G107), .ZN(n466) );
  XNOR2_X1 U371 ( .A(G119), .B(G110), .ZN(n499) );
  XNOR2_X1 U372 ( .A(n483), .B(G125), .ZN(n452) );
  AND2_X2 U373 ( .A1(n535), .A2(n547), .ZN(n576) );
  XNOR2_X2 U374 ( .A(n453), .B(KEYINPUT10), .ZN(n733) );
  NOR2_X2 U375 ( .A1(n561), .A2(n562), .ZN(n365) );
  XNOR2_X2 U376 ( .A(n525), .B(n524), .ZN(n595) );
  XNOR2_X2 U377 ( .A(n341), .B(n340), .ZN(n490) );
  OR2_X2 U378 ( .A1(n616), .A2(G902), .ZN(n341) );
  XNOR2_X2 U379 ( .A(n732), .B(n483), .ZN(n497) );
  AND2_X2 U380 ( .A1(n527), .A2(n369), .ZN(n528) );
  NAND2_X1 U381 ( .A1(n343), .A2(n568), .ZN(n583) );
  XNOR2_X1 U382 ( .A(n558), .B(KEYINPUT72), .ZN(n343) );
  AND2_X2 U383 ( .A1(n681), .A2(n682), .ZN(n602) );
  NOR2_X1 U384 ( .A1(G953), .A2(G237), .ZN(n447) );
  NAND2_X2 U385 ( .A1(n415), .A2(n412), .ZN(n563) );
  XNOR2_X2 U386 ( .A(n517), .B(KEYINPUT33), .ZN(n368) );
  BUF_X1 U387 ( .A(n548), .Z(n601) );
  NOR2_X2 U388 ( .A1(n598), .A2(n550), .ZN(n570) );
  NAND2_X2 U389 ( .A1(n547), .A2(n682), .ZN(n598) );
  NOR2_X2 U390 ( .A1(n686), .A2(n685), .ZN(n682) );
  XNOR2_X2 U391 ( .A(n573), .B(n572), .ZN(n742) );
  NAND2_X2 U392 ( .A1(n591), .A2(n663), .ZN(n734) );
  XNOR2_X2 U393 ( .A(n366), .B(n367), .ZN(n539) );
  AND2_X2 U394 ( .A1(n639), .A2(n458), .ZN(n366) );
  INV_X2 U395 ( .A(G143), .ZN(n420) );
  NOR2_X2 U396 ( .A1(n379), .A2(n376), .ZN(n359) );
  XNOR2_X1 U397 ( .A(n666), .B(KEYINPUT2), .ZN(n379) );
  XNOR2_X1 U398 ( .A(n556), .B(KEYINPUT107), .ZN(n744) );
  XNOR2_X1 U399 ( .A(G110), .B(G107), .ZN(n410) );
  NOR2_X1 U400 ( .A1(n557), .A2(n744), .ZN(n558) );
  XNOR2_X1 U401 ( .A(n571), .B(KEYINPUT39), .ZN(n590) );
  XNOR2_X1 U402 ( .A(n554), .B(n553), .ZN(n555) );
  NOR2_X1 U403 ( .A1(KEYINPUT47), .A2(n543), .ZN(n544) );
  NOR2_X1 U404 ( .A1(n675), .A2(n676), .ZN(n575) );
  NAND2_X1 U405 ( .A1(n673), .A2(n672), .ZN(n676) );
  AND2_X1 U406 ( .A1(n540), .A2(n559), .ZN(n677) );
  NOR2_X1 U407 ( .A1(n712), .A2(G902), .ZN(n510) );
  XNOR2_X1 U408 ( .A(n505), .B(n504), .ZN(n712) );
  XNOR2_X1 U409 ( .A(n502), .B(n371), .ZN(n505) );
  XNOR2_X1 U410 ( .A(G140), .B(n452), .ZN(n453) );
  XNOR2_X1 U411 ( .A(n411), .B(n410), .ZN(n486) );
  XNOR2_X1 U412 ( .A(n409), .B(n426), .ZN(n495) );
  XNOR2_X1 U413 ( .A(KEYINPUT3), .B(G119), .ZN(n409) );
  XNOR2_X1 U414 ( .A(G104), .B(G101), .ZN(n411) );
  INV_X2 U415 ( .A(G146), .ZN(n483) );
  INV_X1 U416 ( .A(n373), .ZN(n345) );
  NOR2_X1 U417 ( .A1(n598), .A2(n550), .ZN(n346) );
  INV_X1 U418 ( .A(n511), .ZN(n347) );
  BUF_X1 U419 ( .A(n461), .Z(n348) );
  NOR2_X2 U420 ( .A1(n621), .A2(n614), .ZN(n360) );
  XNOR2_X2 U421 ( .A(n360), .B(n361), .ZN(n551) );
  INV_X1 U422 ( .A(KEYINPUT86), .ZN(n566) );
  INV_X1 U423 ( .A(KEYINPUT30), .ZN(n401) );
  NOR2_X1 U424 ( .A1(n473), .A2(KEYINPUT82), .ZN(n408) );
  INV_X1 U425 ( .A(KEYINPUT84), .ZN(n386) );
  INV_X1 U426 ( .A(G113), .ZN(n426) );
  XNOR2_X1 U427 ( .A(G122), .B(G116), .ZN(n464) );
  XNOR2_X1 U428 ( .A(n481), .B(n393), .ZN(n392) );
  INV_X1 U429 ( .A(G131), .ZN(n393) );
  NOR2_X1 U430 ( .A1(n437), .A2(KEYINPUT88), .ZN(n413) );
  NAND2_X1 U431 ( .A1(n437), .A2(KEYINPUT88), .ZN(n416) );
  NAND2_X1 U432 ( .A1(n396), .A2(n394), .ZN(n550) );
  AND2_X1 U433 ( .A1(n399), .A2(n397), .ZN(n396) );
  NAND2_X1 U434 ( .A1(n395), .A2(KEYINPUT30), .ZN(n394) );
  XNOR2_X1 U435 ( .A(n497), .B(n389), .ZN(n629) );
  XNOR2_X1 U436 ( .A(n391), .B(n390), .ZN(n389) );
  XNOR2_X1 U437 ( .A(n495), .B(n493), .ZN(n390) );
  XNOR2_X1 U438 ( .A(n496), .B(n494), .ZN(n391) );
  XNOR2_X1 U439 ( .A(n499), .B(KEYINPUT94), .ZN(n372) );
  XNOR2_X1 U440 ( .A(G128), .B(G137), .ZN(n501) );
  XNOR2_X1 U441 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n462) );
  XNOR2_X1 U442 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U443 ( .A(n456), .B(n457), .ZN(n639) );
  AND2_X1 U444 ( .A1(n439), .A2(G953), .ZN(n715) );
  NAND2_X1 U445 ( .A1(n385), .A2(n384), .ZN(n383) );
  AND2_X1 U446 ( .A1(n672), .A2(n401), .ZN(n400) );
  NOR2_X1 U447 ( .A1(n549), .A2(n398), .ZN(n397) );
  NOR2_X1 U448 ( .A1(n672), .A2(n401), .ZN(n398) );
  XOR2_X1 U449 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n493) );
  NAND2_X1 U450 ( .A1(n403), .A2(n407), .ZN(n402) );
  INV_X1 U451 ( .A(n408), .ZN(n403) );
  XNOR2_X1 U452 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n422) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n438) );
  INV_X1 U454 ( .A(KEYINPUT19), .ZN(n356) );
  XNOR2_X1 U455 ( .A(n486), .B(n495), .ZN(n429) );
  XNOR2_X1 U456 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n427) );
  XNOR2_X1 U457 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n465) );
  XOR2_X1 U458 ( .A(G104), .B(G113), .Z(n448) );
  XNOR2_X1 U459 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U460 ( .A(n497), .B(n487), .ZN(n616) );
  INV_X1 U461 ( .A(G953), .ZN(n670) );
  AND2_X1 U462 ( .A1(n576), .A2(n537), .ZN(n653) );
  XNOR2_X1 U463 ( .A(n608), .B(KEYINPUT103), .ZN(n746) );
  XNOR2_X1 U464 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U465 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X1 U466 ( .A1(n539), .A2(n522), .ZN(n349) );
  BUF_X1 U467 ( .A(n551), .Z(n552) );
  AND2_X1 U468 ( .A1(n480), .A2(n526), .ZN(n350) );
  AND2_X1 U469 ( .A1(n681), .A2(n347), .ZN(n351) );
  XOR2_X1 U470 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n352) );
  AND2_X1 U471 ( .A1(n663), .A2(n407), .ZN(n353) );
  XOR2_X1 U472 ( .A(n478), .B(n477), .Z(n354) );
  NAND2_X1 U473 ( .A1(n563), .A2(KEYINPUT19), .ZN(n357) );
  NAND2_X1 U474 ( .A1(n355), .A2(n356), .ZN(n358) );
  NAND2_X1 U475 ( .A1(n357), .A2(n358), .ZN(n536) );
  INV_X1 U476 ( .A(n563), .ZN(n355) );
  NOR2_X1 U477 ( .A1(n379), .A2(n376), .ZN(n707) );
  XOR2_X1 U478 ( .A(n434), .B(KEYINPUT80), .Z(n361) );
  NOR2_X1 U479 ( .A1(n514), .A2(n513), .ZN(n362) );
  NOR2_X1 U480 ( .A1(n514), .A2(n513), .ZN(n592) );
  NAND2_X1 U481 ( .A1(n414), .A2(n413), .ZN(n412) );
  AND2_X1 U482 ( .A1(n405), .A2(n406), .ZN(n363) );
  BUF_X1 U483 ( .A(n527), .Z(n480) );
  XNOR2_X1 U484 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X2 U485 ( .A(n547), .B(KEYINPUT1), .ZN(n681) );
  XNOR2_X1 U486 ( .A(n479), .B(n354), .ZN(n527) );
  AND2_X1 U487 ( .A1(n541), .A2(n537), .ZN(n364) );
  XNOR2_X1 U488 ( .A(n365), .B(KEYINPUT105), .ZN(n585) );
  XOR2_X1 U489 ( .A(n460), .B(n459), .Z(n367) );
  XNOR2_X2 U490 ( .A(n490), .B(G469), .ZN(n547) );
  XNOR2_X2 U491 ( .A(n552), .B(KEYINPUT38), .ZN(n673) );
  INV_X1 U492 ( .A(n733), .ZN(n371) );
  XNOR2_X1 U493 ( .A(n733), .B(n419), .ZN(n456) );
  AND2_X1 U494 ( .A1(n526), .A2(n351), .ZN(n369) );
  NAND2_X1 U495 ( .A1(n548), .A2(n400), .ZN(n399) );
  NAND2_X1 U496 ( .A1(n377), .A2(n363), .ZN(n376) );
  NAND2_X1 U497 ( .A1(n374), .A2(n388), .ZN(n387) );
  NAND2_X1 U498 ( .A1(n716), .A2(n408), .ZN(n405) );
  XNOR2_X1 U499 ( .A(n482), .B(n452), .ZN(n425) );
  XNOR2_X1 U500 ( .A(n370), .B(KEYINPUT28), .ZN(n535) );
  XNOR2_X1 U501 ( .A(n425), .B(n424), .ZN(n430) );
  NOR2_X2 U502 ( .A1(n716), .A2(n734), .ZN(n666) );
  XNOR2_X2 U503 ( .A(n613), .B(n612), .ZN(n716) );
  NAND2_X1 U504 ( .A1(n378), .A2(n373), .ZN(n377) );
  INV_X1 U505 ( .A(n716), .ZN(n373) );
  NAND2_X1 U506 ( .A1(n382), .A2(n383), .ZN(n374) );
  NAND2_X1 U507 ( .A1(n375), .A2(n381), .ZN(n380) );
  INV_X1 U508 ( .A(n583), .ZN(n375) );
  NOR2_X2 U509 ( .A1(n619), .A2(n715), .ZN(n620) );
  NOR2_X2 U510 ( .A1(n642), .A2(n715), .ZN(n643) );
  OR2_X2 U511 ( .A1(n539), .A2(n538), .ZN(n559) );
  NAND2_X1 U512 ( .A1(n404), .A2(n402), .ZN(n406) );
  NOR2_X1 U513 ( .A1(n734), .A2(n614), .ZN(n378) );
  NAND2_X1 U514 ( .A1(n380), .A2(n584), .ZN(n382) );
  INV_X1 U515 ( .A(n582), .ZN(n381) );
  INV_X1 U516 ( .A(n583), .ZN(n384) );
  NOR2_X1 U517 ( .A1(n582), .A2(n584), .ZN(n385) );
  XNOR2_X2 U518 ( .A(n387), .B(n386), .ZN(n591) );
  INV_X1 U519 ( .A(n664), .ZN(n388) );
  XNOR2_X2 U520 ( .A(n461), .B(KEYINPUT4), .ZN(n482) );
  INV_X1 U521 ( .A(n548), .ZN(n395) );
  XNOR2_X2 U522 ( .A(n498), .B(G472), .ZN(n548) );
  NAND2_X1 U523 ( .A1(n591), .A2(n353), .ZN(n404) );
  NAND2_X1 U524 ( .A1(n473), .A2(KEYINPUT82), .ZN(n407) );
  INV_X1 U525 ( .A(n551), .ZN(n414) );
  AND2_X2 U526 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U527 ( .A1(n551), .A2(KEYINPUT88), .ZN(n417) );
  NOR2_X2 U528 ( .A1(n661), .A2(n660), .ZN(n567) );
  BUF_X1 U529 ( .A(n359), .Z(n711) );
  OR2_X1 U530 ( .A1(G902), .A2(n708), .ZN(n418) );
  XOR2_X1 U531 ( .A(n455), .B(n454), .Z(n419) );
  INV_X1 U532 ( .A(n743), .ZN(n579) );
  XNOR2_X1 U533 ( .A(KEYINPUT85), .B(KEYINPUT48), .ZN(n584) );
  INV_X1 U534 ( .A(KEYINPUT45), .ZN(n612) );
  NAND2_X1 U535 ( .A1(n686), .A2(n534), .ZN(n562) );
  BUF_X1 U536 ( .A(n593), .Z(n529) );
  XNOR2_X1 U537 ( .A(G110), .B(KEYINPUT114), .ZN(n515) );
  XNOR2_X2 U538 ( .A(n420), .B(G128), .ZN(n461) );
  NAND2_X1 U539 ( .A1(n670), .A2(G224), .ZN(n421) );
  XNOR2_X1 U540 ( .A(n421), .B(KEYINPUT78), .ZN(n423) );
  XNOR2_X1 U541 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U542 ( .A(n464), .B(n427), .ZN(n428) );
  XNOR2_X1 U543 ( .A(n429), .B(n428), .ZN(n724) );
  XNOR2_X1 U544 ( .A(n430), .B(n724), .ZN(n621) );
  XNOR2_X1 U545 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n431) );
  XNOR2_X1 U546 ( .A(n431), .B(G902), .ZN(n473) );
  INV_X1 U547 ( .A(n473), .ZN(n614) );
  NOR2_X1 U548 ( .A1(G237), .A2(G902), .ZN(n432) );
  XNOR2_X1 U549 ( .A(n432), .B(KEYINPUT74), .ZN(n436) );
  INV_X1 U550 ( .A(G210), .ZN(n433) );
  OR2_X1 U551 ( .A1(n436), .A2(n433), .ZN(n434) );
  INV_X1 U552 ( .A(G214), .ZN(n435) );
  OR2_X1 U553 ( .A1(n436), .A2(n435), .ZN(n672) );
  INV_X1 U554 ( .A(n672), .ZN(n437) );
  INV_X1 U555 ( .A(G952), .ZN(n439) );
  XOR2_X1 U556 ( .A(n438), .B(KEYINPUT14), .Z(n441) );
  NOR2_X1 U557 ( .A1(n439), .A2(n441), .ZN(n699) );
  AND2_X1 U558 ( .A1(n670), .A2(n699), .ZN(n533) );
  INV_X1 U559 ( .A(G898), .ZN(n725) );
  NAND2_X1 U560 ( .A1(G953), .A2(G902), .ZN(n440) );
  NOR2_X1 U561 ( .A1(n441), .A2(n440), .ZN(n530) );
  AND2_X1 U562 ( .A1(n725), .A2(n530), .ZN(n442) );
  NOR2_X1 U563 ( .A1(n533), .A2(n442), .ZN(n443) );
  XNOR2_X1 U564 ( .A(n443), .B(KEYINPUT93), .ZN(n444) );
  NAND2_X1 U565 ( .A1(n536), .A2(n444), .ZN(n446) );
  XNOR2_X1 U566 ( .A(KEYINPUT66), .B(KEYINPUT0), .ZN(n445) );
  XNOR2_X1 U567 ( .A(n446), .B(n445), .ZN(n518) );
  XNOR2_X1 U568 ( .A(n342), .B(G131), .ZN(n451) );
  XOR2_X1 U569 ( .A(KEYINPUT77), .B(n447), .Z(n491) );
  NAND2_X1 U570 ( .A1(G214), .A2(n491), .ZN(n449) );
  XNOR2_X1 U571 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U572 ( .A(n451), .B(n450), .ZN(n457) );
  XOR2_X1 U573 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n455) );
  XNOR2_X1 U574 ( .A(G122), .B(KEYINPUT12), .ZN(n454) );
  INV_X1 U575 ( .A(G902), .ZN(n458) );
  XOR2_X1 U576 ( .A(KEYINPUT13), .B(KEYINPUT100), .Z(n460) );
  XNOR2_X1 U577 ( .A(KEYINPUT99), .B(G475), .ZN(n459) );
  XNOR2_X1 U578 ( .A(KEYINPUT102), .B(G478), .ZN(n472) );
  XNOR2_X1 U579 ( .A(n348), .B(KEYINPUT101), .ZN(n471) );
  NAND2_X1 U580 ( .A1(n670), .A2(G234), .ZN(n463) );
  XNOR2_X1 U581 ( .A(n463), .B(n462), .ZN(n503) );
  NAND2_X1 U582 ( .A1(n503), .A2(G217), .ZN(n469) );
  XNOR2_X1 U583 ( .A(n465), .B(n464), .ZN(n467) );
  XNOR2_X1 U584 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U585 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U586 ( .A(n471), .B(n470), .ZN(n708) );
  XNOR2_X1 U587 ( .A(n472), .B(n418), .ZN(n538) );
  INV_X1 U588 ( .A(n538), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n539), .A2(n522), .ZN(n675) );
  NAND2_X1 U590 ( .A1(G234), .A2(n473), .ZN(n474) );
  XNOR2_X1 U591 ( .A(n474), .B(KEYINPUT20), .ZN(n506) );
  NAND2_X1 U592 ( .A1(G221), .A2(n506), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n475), .B(KEYINPUT21), .ZN(n685) );
  OR2_X1 U594 ( .A1(n675), .A2(n685), .ZN(n476) );
  NOR2_X2 U595 ( .A1(n518), .A2(n476), .ZN(n479) );
  XNOR2_X1 U596 ( .A(KEYINPUT70), .B(KEYINPUT22), .ZN(n478) );
  INV_X1 U597 ( .A(KEYINPUT64), .ZN(n477) );
  INV_X1 U598 ( .A(n480), .ZN(n514) );
  XNOR2_X1 U599 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n489) );
  XNOR2_X1 U600 ( .A(G134), .B(G137), .ZN(n481) );
  NAND2_X1 U601 ( .A1(G227), .A2(n670), .ZN(n484) );
  XNOR2_X1 U602 ( .A(n484), .B(G140), .ZN(n485) );
  XNOR2_X1 U603 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U604 ( .A(n681), .ZN(n660) );
  NAND2_X1 U605 ( .A1(n491), .A2(G210), .ZN(n496) );
  XNOR2_X1 U606 ( .A(G101), .B(G116), .ZN(n492) );
  XNOR2_X1 U607 ( .A(n352), .B(n492), .ZN(n494) );
  OR2_X2 U608 ( .A1(n629), .A2(G902), .ZN(n498) );
  XOR2_X1 U609 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n500) );
  NAND2_X1 U610 ( .A1(G221), .A2(n503), .ZN(n504) );
  NAND2_X1 U611 ( .A1(n506), .A2(G217), .ZN(n508) );
  INV_X1 U612 ( .A(KEYINPUT25), .ZN(n507) );
  INV_X1 U613 ( .A(n686), .ZN(n511) );
  NOR2_X1 U614 ( .A1(n601), .A2(n511), .ZN(n512) );
  NAND2_X1 U615 ( .A1(n660), .A2(n512), .ZN(n513) );
  XOR2_X1 U616 ( .A(n515), .B(n362), .Z(G12) );
  INV_X1 U617 ( .A(KEYINPUT6), .ZN(n516) );
  XNOR2_X1 U618 ( .A(n548), .B(n516), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n602), .A2(n560), .ZN(n517) );
  BUF_X1 U620 ( .A(n518), .Z(n519) );
  INV_X1 U621 ( .A(n519), .ZN(n603) );
  NAND2_X1 U622 ( .A1(n368), .A2(n603), .ZN(n521) );
  XNOR2_X1 U623 ( .A(KEYINPUT79), .B(KEYINPUT34), .ZN(n520) );
  XNOR2_X1 U624 ( .A(n521), .B(n520), .ZN(n523) );
  NAND2_X1 U625 ( .A1(n523), .A2(n349), .ZN(n525) );
  XOR2_X1 U626 ( .A(KEYINPUT83), .B(KEYINPUT35), .Z(n524) );
  XOR2_X1 U627 ( .A(n595), .B(G122), .Z(G24) );
  INV_X1 U628 ( .A(n560), .ZN(n526) );
  XNOR2_X1 U629 ( .A(n528), .B(KEYINPUT32), .ZN(n593) );
  XOR2_X1 U630 ( .A(n529), .B(G119), .Z(G21) );
  XOR2_X1 U631 ( .A(n530), .B(KEYINPUT104), .Z(n531) );
  NOR2_X1 U632 ( .A1(G900), .A2(n531), .ZN(n532) );
  NOR2_X1 U633 ( .A1(n533), .A2(n532), .ZN(n549) );
  NOR2_X1 U634 ( .A1(n685), .A2(n549), .ZN(n534) );
  BUF_X1 U635 ( .A(n536), .Z(n537) );
  AND2_X1 U636 ( .A1(n539), .A2(n538), .ZN(n657) );
  INV_X1 U637 ( .A(n657), .ZN(n540) );
  NOR2_X1 U638 ( .A1(n677), .A2(KEYINPUT73), .ZN(n541) );
  NAND2_X1 U639 ( .A1(n364), .A2(n576), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n542), .A2(KEYINPUT47), .ZN(n546) );
  XOR2_X1 U641 ( .A(KEYINPUT73), .B(n677), .Z(n543) );
  NAND2_X1 U642 ( .A1(n544), .A2(n653), .ZN(n545) );
  NAND2_X1 U643 ( .A1(n546), .A2(n545), .ZN(n557) );
  NAND2_X1 U644 ( .A1(n570), .A2(n414), .ZN(n554) );
  INV_X1 U645 ( .A(KEYINPUT106), .ZN(n553) );
  NAND2_X1 U646 ( .A1(n555), .A2(n349), .ZN(n556) );
  INV_X2 U647 ( .A(n559), .ZN(n655) );
  NAND2_X1 U648 ( .A1(n655), .A2(n560), .ZN(n561) );
  NOR2_X1 U649 ( .A1(n585), .A2(n563), .ZN(n565) );
  INV_X1 U650 ( .A(KEYINPUT36), .ZN(n564) );
  XNOR2_X1 U651 ( .A(n565), .B(n564), .ZN(n661) );
  XNOR2_X1 U652 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U653 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n573) );
  NAND2_X1 U654 ( .A1(n346), .A2(n673), .ZN(n571) );
  NAND2_X1 U655 ( .A1(n655), .A2(n590), .ZN(n572) );
  INV_X1 U656 ( .A(n742), .ZN(n580) );
  XOR2_X1 U657 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n578) );
  XNOR2_X1 U658 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n574) );
  XNOR2_X1 U659 ( .A(n575), .B(n574), .ZN(n694) );
  NAND2_X1 U660 ( .A1(n576), .A2(n694), .ZN(n577) );
  XNOR2_X1 U661 ( .A(n577), .B(n578), .ZN(n743) );
  NAND2_X1 U662 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U663 ( .A(n581), .B(KEYINPUT46), .ZN(n582) );
  INV_X1 U664 ( .A(n585), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n586), .A2(n672), .ZN(n587) );
  NOR2_X1 U666 ( .A1(n681), .A2(n587), .ZN(n588) );
  XNOR2_X1 U667 ( .A(n588), .B(KEYINPUT43), .ZN(n589) );
  NOR2_X1 U668 ( .A1(n589), .A2(n414), .ZN(n664) );
  NAND2_X1 U669 ( .A1(n590), .A2(n657), .ZN(n663) );
  NOR2_X1 U670 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n594), .B(KEYINPUT87), .ZN(n596) );
  NOR2_X2 U672 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT44), .ZN(n611) );
  OR2_X1 U674 ( .A1(n598), .A2(n601), .ZN(n599) );
  NOR2_X1 U675 ( .A1(n519), .A2(n599), .ZN(n600) );
  XNOR2_X1 U676 ( .A(n600), .B(KEYINPUT96), .ZN(n645) );
  AND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n692) );
  NAND2_X1 U678 ( .A1(n692), .A2(n603), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n604), .B(KEYINPUT31), .ZN(n658) );
  NOR2_X1 U680 ( .A1(n645), .A2(n658), .ZN(n605) );
  XOR2_X1 U681 ( .A(KEYINPUT97), .B(n605), .Z(n606) );
  NOR2_X1 U682 ( .A1(n606), .A2(n677), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n347), .A2(n681), .ZN(n607) );
  NAND2_X1 U684 ( .A1(n350), .A2(n607), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n609), .A2(n746), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n707), .A2(G469), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n615) );
  XNOR2_X1 U689 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U690 ( .A(n620), .B(KEYINPUT120), .ZN(G54) );
  NAND2_X1 U691 ( .A1(n359), .A2(G210), .ZN(n625) );
  BUF_X1 U692 ( .A(n621), .Z(n623) );
  XOR2_X1 U693 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n622) );
  XNOR2_X1 U694 ( .A(n625), .B(n624), .ZN(n626) );
  XNOR2_X1 U695 ( .A(n627), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U696 ( .A1(n359), .A2(G472), .ZN(n631) );
  XOR2_X1 U697 ( .A(KEYINPUT89), .B(KEYINPUT62), .Z(n628) );
  XNOR2_X1 U698 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U699 ( .A(KEYINPUT111), .B(KEYINPUT63), .ZN(n633) );
  XOR2_X1 U700 ( .A(n633), .B(KEYINPUT91), .Z(n634) );
  XNOR2_X1 U701 ( .A(n635), .B(n634), .ZN(G57) );
  NAND2_X1 U702 ( .A1(n707), .A2(G475), .ZN(n641) );
  XNOR2_X1 U703 ( .A(KEYINPUT90), .B(KEYINPUT121), .ZN(n637) );
  XNOR2_X1 U704 ( .A(KEYINPUT59), .B(KEYINPUT65), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U706 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U707 ( .A(n643), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U708 ( .A1(n645), .A2(n655), .ZN(n644) );
  XNOR2_X1 U709 ( .A(n644), .B(G104), .ZN(G6) );
  XOR2_X1 U710 ( .A(KEYINPUT113), .B(KEYINPUT26), .Z(n647) );
  NAND2_X1 U711 ( .A1(n657), .A2(n645), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(n649) );
  XOR2_X1 U713 ( .A(G107), .B(KEYINPUT27), .Z(n648) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(G9) );
  XOR2_X1 U715 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n651) );
  NAND2_X1 U716 ( .A1(n653), .A2(n657), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U718 ( .A(G128), .B(n652), .Z(G30) );
  NAND2_X1 U719 ( .A1(n653), .A2(n655), .ZN(n654) );
  XNOR2_X1 U720 ( .A(n654), .B(G146), .ZN(G48) );
  NAND2_X1 U721 ( .A1(n658), .A2(n655), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n656), .B(G113), .ZN(G15) );
  NAND2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U724 ( .A(n659), .B(G116), .ZN(G18) );
  XNOR2_X1 U725 ( .A(n567), .B(G125), .ZN(n662) );
  XNOR2_X1 U726 ( .A(n662), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U727 ( .A(G134), .B(n663), .ZN(G36) );
  XNOR2_X1 U728 ( .A(n664), .B(G140), .ZN(n665) );
  XNOR2_X1 U729 ( .A(n665), .B(KEYINPUT117), .ZN(G42) );
  NOR2_X1 U730 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n667) );
  XNOR2_X1 U731 ( .A(n666), .B(n667), .ZN(n669) );
  NAND2_X1 U732 ( .A1(KEYINPUT2), .A2(KEYINPUT81), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n671), .A2(n670), .ZN(n705) );
  NAND2_X1 U735 ( .A1(n368), .A2(n694), .ZN(n702) );
  NOR2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U737 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  OR2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U740 ( .A1(n368), .A2(n680), .ZN(n697) );
  OR2_X1 U741 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U742 ( .A(n683), .B(KEYINPUT50), .ZN(n684) );
  NAND2_X1 U743 ( .A1(n684), .A2(n395), .ZN(n689) );
  NAND2_X1 U744 ( .A1(n347), .A2(n685), .ZN(n687) );
  XNOR2_X1 U745 ( .A(KEYINPUT49), .B(n687), .ZN(n688) );
  NOR2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U747 ( .A(n690), .B(KEYINPUT118), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U749 ( .A(KEYINPUT51), .B(n693), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U751 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U752 ( .A(KEYINPUT52), .B(n698), .ZN(n700) );
  NAND2_X1 U753 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U754 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U755 ( .A(KEYINPUT119), .B(n703), .Z(n704) );
  NOR2_X1 U756 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U757 ( .A(KEYINPUT53), .B(n706), .ZN(G75) );
  NAND2_X1 U758 ( .A1(n711), .A2(G478), .ZN(n709) );
  XNOR2_X1 U759 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U760 ( .A1(n715), .A2(n710), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n711), .A2(G217), .ZN(n713) );
  XNOR2_X1 U762 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n715), .A2(n714), .ZN(G66) );
  NOR2_X1 U764 ( .A1(n345), .A2(G953), .ZN(n717) );
  XNOR2_X1 U765 ( .A(n717), .B(KEYINPUT124), .ZN(n723) );
  NAND2_X1 U766 ( .A1(G224), .A2(G953), .ZN(n718) );
  XNOR2_X1 U767 ( .A(n718), .B(KEYINPUT61), .ZN(n719) );
  XNOR2_X1 U768 ( .A(KEYINPUT122), .B(n719), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n720), .A2(G898), .ZN(n721) );
  XNOR2_X1 U770 ( .A(KEYINPUT123), .B(n721), .ZN(n722) );
  NOR2_X1 U771 ( .A1(n723), .A2(n722), .ZN(n729) );
  INV_X1 U772 ( .A(n724), .ZN(n727) );
  NAND2_X1 U773 ( .A1(n725), .A2(G953), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U775 ( .A(n729), .B(n728), .ZN(n731) );
  XOR2_X1 U776 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n730) );
  XNOR2_X1 U777 ( .A(n731), .B(n730), .ZN(G69) );
  XNOR2_X1 U778 ( .A(n733), .B(n732), .ZN(n737) );
  XOR2_X1 U779 ( .A(n737), .B(n734), .Z(n735) );
  NOR2_X1 U780 ( .A1(G953), .A2(n735), .ZN(n736) );
  XNOR2_X1 U781 ( .A(n736), .B(KEYINPUT127), .ZN(n741) );
  XNOR2_X1 U782 ( .A(G227), .B(n737), .ZN(n738) );
  NAND2_X1 U783 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U784 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U785 ( .A1(n741), .A2(n740), .ZN(G72) );
  XOR2_X1 U786 ( .A(n742), .B(G131), .Z(G33) );
  XOR2_X1 U787 ( .A(G137), .B(n743), .Z(G39) );
  XOR2_X1 U788 ( .A(n342), .B(n744), .Z(n745) );
  XNOR2_X1 U789 ( .A(KEYINPUT116), .B(n745), .ZN(G45) );
  XOR2_X1 U790 ( .A(G101), .B(n746), .Z(n747) );
  XNOR2_X1 U791 ( .A(KEYINPUT112), .B(n747), .ZN(G3) );
endmodule

