//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n632,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT68), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G125), .C1(new_n467), .C2(new_n468), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n471), .B1(new_n477), .B2(G2105), .ZN(G160));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n464), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  MUX2_X1   g057(.A(G100), .B(G112), .S(G2105), .Z(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(G136), .B2(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g064(.A(G138), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n486), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n469), .B2(new_n490), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT69), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n499), .A2(new_n500), .A3(G126), .A4(G2105), .ZN(new_n501));
  MUX2_X1   g076(.A(G102), .B(G114), .S(G2105), .Z(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2104), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n498), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n496), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI211_X1 g082(.A(KEYINPUT72), .B(new_n506), .C1(new_n507), .C2(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT5), .B1(new_n507), .B2(KEYINPUT72), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT71), .B1(new_n514), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(G651), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(new_n518), .B1(KEYINPUT6), .B2(new_n514), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n506), .B1(new_n509), .B2(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT72), .B1(new_n507), .B2(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n522), .B1(new_n525), .B2(new_n508), .ZN(new_n526));
  AND2_X1   g101(.A1(G75), .A2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(G651), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(G50), .A3(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G166));
  NAND2_X1  g106(.A1(new_n520), .A2(G89), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n519), .A2(G543), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT74), .B(G51), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n532), .A2(new_n535), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(KEYINPUT75), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(G168));
  NAND2_X1  g117(.A1(new_n513), .A2(new_n519), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT76), .B(G90), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n519), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n514), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(G171));
  NAND2_X1  g125(.A1(new_n520), .A2(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n533), .A2(G43), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n551), .B(new_n552), .C1(new_n514), .C2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n519), .A2(G53), .A3(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n519), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n520), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n513), .A2(KEYINPUT77), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n525), .A2(new_n570), .A3(new_n508), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(G65), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n514), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  INV_X1    g154(.A(new_n528), .ZN(new_n580));
  INV_X1    g155(.A(G88), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n529), .B1(new_n543), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n579), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n521), .A2(new_n528), .A3(KEYINPUT78), .A4(new_n529), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n520), .A2(G87), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n533), .A2(G49), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  INV_X1    g166(.A(G48), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n543), .A2(new_n591), .B1(new_n545), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n513), .A2(G61), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n513), .A2(KEYINPUT79), .A3(G61), .ZN(new_n597));
  NAND2_X1  g172(.A1(G73), .A2(G543), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n593), .B1(new_n599), .B2(G651), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G305));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n543), .A2(new_n602), .B1(new_n545), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n605), .A2(KEYINPUT80), .A3(new_n514), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT80), .B1(new_n605), .B2(new_n514), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n604), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G301), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n543), .B2(new_n614), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n612), .A2(new_n615), .B1(G54), .B2(new_n533), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n569), .A2(new_n571), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n617), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G651), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n618), .A2(new_n619), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n611), .B1(new_n624), .B2(new_n610), .ZN(G284));
  AOI21_X1  g200(.A(new_n611), .B1(new_n624), .B2(new_n610), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT82), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n575), .B(KEYINPUT83), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(G868), .B2(new_n629), .ZN(G297));
  XOR2_X1   g205(.A(G297), .B(KEYINPUT84), .Z(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n624), .B1(new_n632), .B2(G860), .ZN(G148));
  OAI211_X1 g208(.A(new_n632), .B(new_n616), .C1(new_n621), .C2(new_n622), .ZN(new_n634));
  MUX2_X1   g209(.A(new_n554), .B(new_n634), .S(G868), .Z(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n486), .A2(G2104), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n640), .A2(KEYINPUT13), .B1(KEYINPUT86), .B2(G2100), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(KEYINPUT13), .B2(new_n640), .ZN(new_n642));
  OR3_X1    g217(.A1(new_n642), .A2(KEYINPUT86), .A3(G2100), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n642), .B1(KEYINPUT86), .B2(G2100), .ZN(new_n644));
  MUX2_X1   g219(.A(G99), .B(G111), .S(G2105), .Z(new_n645));
  AOI22_X1  g220(.A1(G123), .A2(new_n481), .B1(new_n645), .B2(G2104), .ZN(new_n646));
  INV_X1    g221(.A(G135), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n647), .B2(new_n469), .ZN(new_n648));
  INV_X1    g223(.A(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(G156));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2427), .ZN(new_n656));
  INV_X1    g231(.A(G2430), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(G14), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT88), .ZN(G401));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT89), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  OR2_X1    g251(.A1(new_n671), .A2(new_n674), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n673), .B1(new_n677), .B2(KEYINPUT17), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(KEYINPUT17), .ZN(new_n679));
  INV_X1    g254(.A(new_n674), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(new_n671), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n680), .B2(new_n679), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n676), .B1(new_n678), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n649), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2100), .ZN(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n688), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1981), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT90), .ZN(new_n701));
  XOR2_X1   g276(.A(G1991), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n699), .B(new_n703), .ZN(G229));
  XNOR2_X1  g279(.A(KEYINPUT91), .B(G29), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G27), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G164), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G2078), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT31), .B(G11), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT30), .B(G28), .Z(new_n711));
  OAI221_X1 g286(.A(new_n710), .B1(G29), .B2(new_n711), .C1(new_n648), .C2(new_n705), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT26), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n486), .A2(G141), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n481), .A2(G129), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n714), .B(new_n717), .C1(G105), .C2(new_n465), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G29), .ZN(new_n719));
  NOR2_X1   g294(.A1(G29), .A2(G32), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(KEYINPUT96), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT96), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n712), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n705), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n486), .A2(G140), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n481), .A2(G128), .ZN(new_n728));
  MUX2_X1   g303(.A(G104), .B(G116), .S(G2105), .Z(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G2104), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n726), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G2067), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n724), .B(new_n736), .C1(new_n722), .C2(new_n723), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  NOR2_X1   g314(.A1(G171), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G5), .B2(new_n739), .ZN(new_n741));
  AOI211_X1 g316(.A(new_n709), .B(new_n737), .C1(new_n738), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n733), .A2(G33), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n499), .A2(G127), .ZN(new_n748));
  NAND2_X1  g323(.A1(G115), .A2(G2104), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n464), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n465), .A2(G103), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT25), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n750), .B(new_n752), .C1(G139), .C2(new_n486), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT95), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n747), .B1(new_n754), .B2(new_n733), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G2072), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n739), .A2(G19), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n554), .B2(G16), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(G1341), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT24), .B(G34), .ZN(new_n762));
  AOI22_X1  g337(.A1(G160), .A2(G29), .B1(new_n705), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2084), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n741), .B2(new_n738), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n708), .A2(G2078), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G2084), .B2(new_n763), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n706), .A2(G35), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G162), .B2(new_n706), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT98), .Z(new_n770));
  XOR2_X1   g345(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n765), .B(new_n767), .C1(new_n772), .C2(G2090), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n742), .A2(new_n746), .A3(new_n761), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G4), .A2(G16), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n624), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1348), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G21), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G168), .B2(G16), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G1966), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(G1966), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n780), .B(new_n781), .C1(new_n772), .C2(G2090), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n774), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G24), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n608), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT93), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1986), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G22), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G166), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n739), .A2(G23), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n589), .B2(new_n739), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT33), .B(G1976), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G6), .A2(G16), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n600), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(KEYINPUT34), .B1(new_n796), .B2(new_n800), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT92), .B1(G95), .B2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NOR3_X1   g381(.A1(KEYINPUT92), .A2(G95), .A3(G2105), .ZN(new_n807));
  OAI221_X1 g382(.A(G2104), .B1(G107), .B2(new_n464), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n486), .A2(G131), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n481), .A2(G119), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(new_n706), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n787), .A2(new_n803), .A3(new_n804), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT36), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n783), .A2(new_n816), .ZN(G150));
  XNOR2_X1  g392(.A(G150), .B(KEYINPUT99), .ZN(G311));
  AOI22_X1  g393(.A1(G93), .A2(new_n520), .B1(new_n533), .B2(G55), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n514), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT102), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n624), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n821), .B(new_n554), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT101), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n827), .B(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n831), .B2(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n824), .B1(new_n832), .B2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(G162), .B(G160), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n648), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT103), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n493), .B1(new_n486), .B2(new_n491), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n469), .A2(new_n490), .A3(new_n492), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n504), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n494), .A2(new_n495), .A3(KEYINPUT103), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n732), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n481), .A2(G130), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT104), .Z(new_n848));
  INV_X1    g423(.A(G118), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n849), .A2(KEYINPUT105), .A3(G2105), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT105), .B1(new_n849), .B2(G2105), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n850), .A2(new_n853), .B1(new_n486), .B2(G142), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n811), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n856), .A2(new_n640), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n856), .A2(new_n640), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n846), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n754), .B(new_n718), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n857), .A2(new_n858), .A3(new_n846), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n857), .A2(new_n858), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n845), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n861), .B1(new_n866), .B2(new_n859), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n837), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n860), .B2(new_n863), .ZN(new_n870));
  INV_X1    g445(.A(new_n837), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n866), .A2(new_n859), .A3(new_n861), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n868), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g450(.A(new_n608), .B(new_n589), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n600), .B(G166), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n623), .A2(G299), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n514), .B1(new_n618), .B2(new_n619), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n619), .B2(new_n618), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n575), .B1(new_n882), .B2(new_n616), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n879), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n623), .A2(G299), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n575), .A3(new_n616), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n826), .A2(new_n632), .A3(new_n882), .A4(new_n616), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n555), .B(new_n821), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n634), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n880), .A2(new_n883), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n888), .A3(new_n890), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n878), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n892), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n900));
  INV_X1    g475(.A(new_n878), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n898), .A2(new_n903), .A3(G868), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT106), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n898), .A2(new_n903), .A3(new_n906), .A4(G868), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n821), .A2(new_n610), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(G295));
  AND2_X1   g484(.A1(new_n904), .A2(KEYINPUT106), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT107), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n905), .A2(new_n913), .A3(new_n907), .A4(new_n908), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(G331));
  XNOR2_X1  g490(.A(G168), .B(G301), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n826), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n894), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n884), .A2(new_n887), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n918), .B(new_n878), .C1(new_n919), .C2(new_n917), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n869), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n917), .A2(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n878), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n918), .B1(new_n919), .B2(new_n917), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n901), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n869), .A4(new_n920), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n844), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n475), .A2(new_n476), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n474), .B1(new_n499), .B2(G125), .ZN(new_n936));
  OAI21_X1  g511(.A(G2105), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n471), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(G40), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n933), .B1(new_n496), .B2(new_n504), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n940), .B2(KEYINPUT50), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n738), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n844), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n939), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G2078), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(KEYINPUT121), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT121), .B1(new_n948), .B2(new_n949), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G40), .ZN(new_n954));
  AOI211_X1 g529(.A(new_n954), .B(new_n471), .C1(new_n477), .C2(G2105), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n949), .A2(G2078), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n504), .B1(new_n838), .B2(new_n496), .ZN(new_n957));
  AOI21_X1  g532(.A(G1384), .B1(new_n957), .B2(new_n843), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n955), .B(new_n956), .C1(new_n958), .C2(KEYINPUT45), .ZN(new_n959));
  INV_X1    g534(.A(new_n944), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT122), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n844), .A2(new_n933), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n939), .B1(new_n962), .B2(new_n945), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT122), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n964), .A3(new_n944), .A4(new_n956), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(G171), .B1(new_n953), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n948), .A2(new_n949), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT121), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n950), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT45), .B(new_n933), .C1(new_n496), .C2(new_n504), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n963), .A2(new_n972), .A3(new_n956), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n971), .A2(G301), .A3(new_n973), .A4(new_n943), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n967), .A2(KEYINPUT54), .A3(new_n974), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n955), .B(new_n972), .C1(new_n958), .C2(KEYINPUT45), .ZN(new_n976));
  INV_X1    g551(.A(G1966), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G2084), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n934), .A2(new_n941), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT115), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n934), .A2(new_n941), .A3(new_n982), .A4(new_n979), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n978), .A2(new_n981), .A3(G168), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(KEYINPUT120), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT51), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n989), .A3(new_n986), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n978), .A2(new_n981), .A3(new_n983), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(G8), .A3(G286), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n973), .B(new_n943), .C1(new_n951), .C2(new_n952), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G171), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n961), .A2(new_n965), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n971), .A2(new_n996), .A3(G301), .A4(new_n943), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT54), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n975), .B(new_n993), .C1(new_n998), .C2(KEYINPUT123), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n589), .A2(G1976), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n844), .A2(new_n955), .A3(new_n933), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(G8), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT110), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1005), .A3(G8), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1001), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n1008));
  INV_X1    g583(.A(G1976), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G288), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1007), .A2(KEYINPUT111), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(G305), .A2(G1981), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n600), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n597), .A2(new_n598), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT79), .B1(new_n513), .B2(G61), .ZN(new_n1017));
  OAI21_X1  g592(.A(G651), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n593), .ZN(new_n1019));
  AND4_X1   g594(.A1(new_n1013), .A2(new_n1018), .A3(new_n1019), .A4(new_n1014), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1012), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1012), .B(KEYINPUT49), .C1(new_n1015), .C2(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1011), .A2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1002), .A2(new_n1005), .A3(G8), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1005), .B1(new_n1002), .B2(G8), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1000), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1009), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1031), .A2(KEYINPUT111), .B1(new_n1007), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT114), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT111), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1007), .A2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1011), .A4(new_n1026), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1971), .B1(new_n944), .B2(new_n946), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n934), .A2(new_n941), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT108), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n583), .A2(new_n584), .A3(G8), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(KEYINPUT109), .A3(new_n1047), .ZN(new_n1051));
  NAND3_X1  g626(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT108), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1041), .A2(new_n1054), .A3(new_n1043), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1045), .A2(new_n1053), .A3(G8), .A4(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1052), .A2(new_n1051), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n844), .A2(KEYINPUT50), .A3(new_n933), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n940), .A2(new_n932), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n939), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1040), .B1(new_n1042), .B2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1057), .B(new_n1050), .C1(new_n1061), .C2(new_n985), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1034), .A2(new_n1039), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1065), .B(KEYINPUT54), .C1(new_n995), .C2(new_n997), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n999), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT60), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1002), .A2(G2067), .ZN(new_n1069));
  INV_X1    g644(.A(G1348), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1069), .B1(new_n942), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n624), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n624), .B(new_n1071), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n1068), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n944), .A2(new_n946), .A3(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1060), .B2(G1956), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n572), .A2(new_n573), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G651), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n566), .A4(new_n567), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT57), .B1(new_n568), .B2(new_n574), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n1076), .C1(G1956), .C2(new_n1060), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1084), .A2(new_n1086), .A3(KEYINPUT61), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT61), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  INV_X1    g665(.A(G1996), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n944), .A2(new_n946), .A3(new_n1091), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT58), .B(G1341), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n958), .B2(new_n955), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1002), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT118), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1092), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1090), .B1(new_n1105), .B2(new_n555), .ZN(new_n1106));
  AOI211_X1 g681(.A(KEYINPUT59), .B(new_n554), .C1(new_n1100), .C2(new_n1104), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1089), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT119), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1089), .B(new_n1110), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1074), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1086), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1071), .A2(new_n623), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(KEYINPUT116), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1115), .A2(KEYINPUT116), .B1(new_n1077), .B2(new_n1083), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1113), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1067), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n990), .A2(new_n992), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n989), .B1(new_n984), .B2(new_n986), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT62), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n988), .A2(new_n1123), .A3(new_n990), .A4(new_n992), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(new_n1124), .A3(G171), .A4(new_n994), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1125), .A2(new_n1064), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n589), .A2(new_n1009), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1021), .A2(new_n1022), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1128), .B1(new_n1129), .B2(new_n1025), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1024), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1037), .A2(new_n1011), .A3(new_n1026), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1133), .B2(new_n1056), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT113), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1132), .B(KEYINPUT113), .C1(new_n1133), .C2(new_n1056), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1127), .A2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n991), .A2(G8), .A3(G168), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1064), .A2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1056), .A2(new_n1140), .A3(KEYINPUT63), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1045), .A2(G8), .A3(new_n1055), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1143), .B1(new_n1053), .B2(new_n1144), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1142), .A2(KEYINPUT63), .B1(new_n1133), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1126), .B1(new_n1125), .B2(new_n1064), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1119), .A2(new_n1139), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n958), .A2(KEYINPUT45), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n955), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n718), .B(G1996), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n731), .B(new_n735), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(G290), .A2(G1986), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n811), .B(new_n813), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G290), .A2(G1986), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1151), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1148), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1150), .B1(new_n718), .B2(new_n1153), .ZN(new_n1161));
  OR3_X1    g736(.A1(new_n1150), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT46), .B1(new_n1150), .B2(G1996), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT47), .Z(new_n1165));
  INV_X1    g740(.A(new_n811), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(new_n813), .C1(new_n1154), .C2(new_n1150), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n732), .A2(new_n735), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT125), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(KEYINPUT125), .A3(new_n1168), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1151), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1165), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1151), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1151), .A2(new_n1158), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT126), .Z(new_n1176));
  OAI21_X1  g751(.A(new_n1174), .B1(new_n1176), .B2(KEYINPUT48), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1177), .B1(KEYINPUT48), .B2(new_n1176), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1172), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1160), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n1182));
  NOR4_X1   g756(.A1(G401), .A2(G227), .A3(G229), .A4(new_n462), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n874), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g758(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1182), .B1(new_n929), .B2(new_n1185), .ZN(new_n1186));
  AOI211_X1 g760(.A(KEYINPUT127), .B(new_n1184), .C1(new_n924), .C2(new_n928), .ZN(new_n1187));
  NOR2_X1   g761(.A1(new_n1186), .A2(new_n1187), .ZN(G308));
  NAND2_X1  g762(.A1(new_n929), .A2(new_n1185), .ZN(G225));
endmodule


