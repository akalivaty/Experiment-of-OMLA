//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930;
  XNOR2_X1  g000(.A(KEYINPUT71), .B(G218gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT22), .B1(new_n202), .B2(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G197gat), .B(G204gat), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(KEYINPUT72), .A3(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(new_n203), .B2(new_n205), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n210), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n204), .A2(KEYINPUT72), .A3(new_n206), .A4(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT28), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT65), .B(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n220), .B2(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n215), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n216), .A2(new_n219), .A3(KEYINPUT28), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT26), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT26), .ZN(new_n231));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n225), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G226gat), .ZN(new_n238));
  INV_X1    g037(.A(G233gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(G176gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(new_n226), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n243), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT23), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n228), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n234), .A2(KEYINPUT24), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT24), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  INV_X1    g052(.A(G183gat), .ZN(new_n254));
  INV_X1    g053(.A(G190gat), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n251), .A2(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n241), .B1(new_n250), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G190gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n260), .A3(new_n254), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n251), .A2(new_n253), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n241), .B1(new_n229), .B2(KEYINPUT23), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(new_n249), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n257), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n237), .A2(new_n240), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n235), .B1(new_n223), .B2(new_n224), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n257), .A2(new_n270), .A3(new_n265), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n240), .A2(KEYINPUT29), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n214), .B(new_n267), .C1(new_n272), .C2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n257), .A2(new_n270), .A3(new_n265), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n270), .B1(new_n257), .B2(new_n265), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n237), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n240), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n268), .B1(new_n257), .B2(new_n265), .ZN(new_n281));
  OAI22_X1  g080(.A1(new_n279), .A2(new_n280), .B1(new_n281), .B2(new_n274), .ZN(new_n282));
  INV_X1    g081(.A(new_n214), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n273), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n285), .A2(new_n286), .A3(new_n214), .A4(new_n267), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT84), .B(KEYINPUT37), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n276), .A2(new_n284), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G8gat), .B(G36gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n283), .A3(new_n267), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT37), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n214), .B2(new_n282), .ZN(new_n299));
  OR3_X1    g098(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT38), .ZN(new_n300));
  NOR2_X1   g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT78), .B1(new_n306), .B2(new_n301), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT2), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G155gat), .ZN(new_n310));
  INV_X1    g109(.A(G162gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT77), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT77), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G155gat), .B2(G162gat), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n312), .A2(new_n314), .B1(G155gat), .B2(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT68), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n319), .B(new_n321), .C1(G113gat), .C2(new_n320), .ZN(new_n322));
  INV_X1    g121(.A(G134gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G127gat), .ZN(new_n324));
  INV_X1    g123(.A(G127gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327));
  AND3_X1   g126(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n318), .A2(G120gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n320), .A2(G113gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n324), .A2(new_n326), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n322), .A2(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(new_n310), .B2(new_n311), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n306), .A2(new_n301), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n316), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT4), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n309), .A2(new_n315), .B1(new_n336), .B2(new_n335), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n342));
  INV_X1    g141(.A(new_n333), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n316), .A2(new_n344), .A3(new_n337), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n340), .B(new_n342), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT79), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n338), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n341), .A2(new_n333), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT5), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n316), .A2(new_n337), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n344), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n343), .A3(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n360), .A2(new_n348), .A3(new_n340), .A4(new_n342), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n361), .A2(new_n354), .A3(KEYINPUT79), .ZN(new_n362));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n356), .A2(new_n362), .A3(KEYINPUT6), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n356), .A2(new_n362), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n366), .B(KEYINPUT83), .ZN(new_n370));
  OR2_X1    g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n366), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT6), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n368), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT37), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n284), .A2(new_n287), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n377), .B2(new_n276), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT38), .B1(new_n378), .B2(new_n296), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n276), .A2(new_n284), .A3(new_n287), .A4(new_n294), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT76), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n300), .A2(new_n374), .A3(new_n379), .A4(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT31), .B(G50gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  XOR2_X1   g184(.A(new_n385), .B(KEYINPUT80), .Z(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n211), .A2(new_n387), .A3(new_n213), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(new_n344), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n357), .ZN(new_n390));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(KEYINPUT81), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n359), .A2(new_n387), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n214), .A2(new_n394), .B1(KEYINPUT81), .B2(new_n391), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n214), .A2(new_n394), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n391), .A2(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n341), .B1(new_n388), .B2(new_n344), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n392), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT82), .B(G22gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n396), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n396), .B2(new_n401), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n386), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n385), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n396), .A2(new_n401), .A3(G22gat), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n396), .A2(new_n401), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(new_n403), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n295), .B1(new_n376), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n413), .B1(new_n414), .B2(new_n380), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n381), .B2(new_n414), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n347), .A2(new_n349), .ZN(new_n417));
  OR3_X1    g216(.A1(new_n351), .A2(new_n352), .A3(new_n349), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT39), .A3(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n419), .B(new_n370), .C1(KEYINPUT39), .C2(new_n417), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT40), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n371), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n382), .B(new_n411), .C1(new_n416), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n362), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n354), .B1(new_n361), .B2(KEYINPUT79), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n372), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n356), .A2(new_n362), .A3(new_n366), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n367), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n377), .A2(KEYINPUT76), .A3(new_n276), .A4(new_n294), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT76), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n380), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n414), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n294), .B1(new_n377), .B2(new_n276), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n380), .A2(new_n414), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n430), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n411), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n279), .A2(new_n333), .ZN(new_n441));
  INV_X1    g240(.A(G227gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n239), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n343), .B(new_n237), .C1(new_n277), .C2(new_n278), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT69), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT69), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  XNOR2_X1  g249(.A(G15gat), .B(G43gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n445), .B2(KEYINPUT32), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n445), .B(KEYINPUT32), .C1(new_n446), .C2(new_n453), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n443), .B1(new_n441), .B2(new_n444), .ZN(new_n457));
  XOR2_X1   g256(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n455), .B2(new_n456), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n462), .A2(KEYINPUT36), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(KEYINPUT36), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n423), .A2(new_n440), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n411), .B1(new_n460), .B2(new_n461), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT35), .B1(new_n466), .B2(new_n438), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n455), .A2(new_n456), .ZN(new_n468));
  INV_X1    g267(.A(new_n459), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n426), .B(new_n427), .C1(new_n369), .C2(new_n370), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT35), .B1(new_n473), .B2(new_n367), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(new_n416), .A3(new_n411), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n465), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G22gat), .ZN(new_n479));
  INV_X1    g278(.A(G1gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT16), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n480), .B2(new_n479), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT88), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(G8gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n482), .B2(KEYINPUT88), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g286(.A(KEYINPUT88), .B(new_n485), .C1(new_n482), .C2(new_n483), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G43gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(G50gat), .ZN(new_n491));
  INV_X1    g290(.A(G50gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n492), .A2(G43gat), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT86), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT86), .B1(new_n491), .B2(new_n493), .ZN(new_n497));
  INV_X1    g296(.A(G29gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n499));
  AND2_X1   g298(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n500));
  NOR2_X1   g299(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n502), .B2(G36gat), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n496), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n490), .A2(G50gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(new_n491), .B2(KEYINPUT87), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n507), .A2(new_n490), .A3(G50gat), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n495), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n496), .A2(new_n497), .B1(new_n509), .B2(new_n503), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT17), .B1(new_n504), .B2(new_n510), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n484), .A2(G8gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n484), .B2(new_n486), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n517), .A2(new_n518), .A3(new_n511), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n517), .B2(new_n511), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n478), .B(new_n515), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n511), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT90), .B1(new_n489), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n517), .A2(new_n518), .A3(new_n511), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n527), .A2(KEYINPUT18), .A3(new_n478), .A4(new_n515), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n489), .A2(new_n524), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n519), .B2(new_n520), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n478), .B(KEYINPUT13), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n523), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G113gat), .B(G141gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G197gat), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT11), .B(G169gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT85), .B(KEYINPUT12), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n523), .A2(new_n532), .A3(new_n528), .A4(new_n539), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n477), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546));
  XOR2_X1   g345(.A(G99gat), .B(G106gat), .Z(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  INV_X1    g351(.A(G92gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(KEYINPUT8), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n548), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n548), .A2(new_n550), .A3(new_n554), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(KEYINPUT94), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n559));
  INV_X1    g358(.A(new_n557), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n555), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n511), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT92), .Z(new_n566));
  INV_X1    g365(.A(KEYINPUT41), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n546), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n563), .B(KEYINPUT95), .C1(new_n567), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n513), .A2(new_n514), .A3(new_n558), .A4(new_n561), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT96), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n573), .B2(new_n574), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n566), .A2(new_n567), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G134gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G162gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n578), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n575), .A2(new_n579), .A3(new_n577), .A4(new_n583), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G57gat), .B(G64gat), .Z(new_n589));
  INV_X1    g388(.A(KEYINPUT9), .ZN(new_n590));
  INV_X1    g389(.A(G71gat), .ZN(new_n591));
  INV_X1    g390(.A(G78gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G71gat), .B(G78gat), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n594), .B(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n517), .B1(KEYINPUT21), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT91), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n597), .A2(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G127gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n599), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n604), .B(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n597), .B1(new_n560), .B2(new_n555), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n594), .B(new_n595), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(new_n557), .A3(new_n556), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT10), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n597), .A2(KEYINPUT10), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n558), .B2(new_n561), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n610), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n610), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n613), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n617), .A2(KEYINPUT97), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626));
  OAI211_X1 g425(.A(new_n626), .B(new_n610), .C1(new_n614), .C2(new_n616), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n624), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n623), .B1(new_n628), .B2(new_n622), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n588), .A2(new_n609), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n545), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(new_n430), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT98), .B(G1gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(G1324gat));
  INV_X1    g433(.A(new_n631), .ZN(new_n635));
  INV_X1    g434(.A(new_n416), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT16), .B(G8gat), .Z(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n485), .B1(new_n635), .B2(new_n636), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT42), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n641), .B1(KEYINPUT42), .B2(new_n639), .ZN(G1325gat));
  NAND2_X1  g441(.A1(new_n463), .A2(new_n464), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(G15gat), .B1(new_n631), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n462), .A2(G15gat), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n645), .B1(new_n631), .B2(new_n646), .ZN(G1326gat));
  NOR2_X1   g446(.A1(new_n631), .A2(new_n411), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT43), .B(G22gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(G1327gat));
  INV_X1    g449(.A(new_n629), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n609), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n587), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n545), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n430), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n498), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n541), .A2(new_n659), .A3(new_n542), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n659), .B1(new_n541), .B2(new_n542), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n652), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n467), .A2(new_n666), .A3(new_n475), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n467), .B2(new_n475), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n465), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT101), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n465), .B(new_n671), .C1(new_n667), .C2(new_n668), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n587), .A2(KEYINPUT44), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT44), .B1(new_n477), .B2(new_n587), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n665), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G29gat), .B1(new_n677), .B2(new_n430), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n658), .A2(new_n678), .ZN(G1328gat));
  AOI21_X1  g478(.A(G36gat), .B1(KEYINPUT102), .B2(KEYINPUT46), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n655), .A2(new_n636), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G36gat), .B1(new_n677), .B2(new_n416), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n676), .A2(new_n643), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n462), .A2(G43gat), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n687), .A2(G43gat), .B1(new_n655), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n686), .B(KEYINPUT47), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n689), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT104), .B1(new_n692), .B2(KEYINPUT103), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n694), .B1(new_n692), .B2(KEYINPUT104), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n691), .B1(new_n693), .B2(new_n695), .ZN(G1330gat));
  NAND3_X1  g495(.A1(new_n655), .A2(new_n492), .A3(new_n439), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n411), .B(new_n665), .C1(new_n674), .C2(new_n675), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT48), .B(new_n697), .C1(new_n698), .C2(new_n492), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT105), .B1(new_n698), .B2(new_n492), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n674), .A2(new_n675), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n439), .A3(new_n664), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n703), .A3(G50gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n704), .A3(new_n697), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(new_n705), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n699), .B1(new_n708), .B2(new_n709), .ZN(G1331gat));
  AND2_X1   g509(.A1(new_n670), .A2(new_n672), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n588), .A2(new_n609), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n629), .A3(new_n663), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n711), .A2(KEYINPUT107), .A3(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n656), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g521(.A1(new_n719), .A2(new_n416), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(G1333gat));
  NAND3_X1  g526(.A1(new_n720), .A2(new_n591), .A3(new_n472), .ZN(new_n728));
  OAI21_X1  g527(.A(G71gat), .B1(new_n719), .B2(new_n644), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT50), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1334gat));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n411), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT108), .B(G78gat), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1335gat));
  INV_X1    g536(.A(new_n609), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n738), .A2(new_n662), .A3(new_n651), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n701), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740), .B2(new_n430), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n669), .A2(new_n588), .A3(new_n609), .A4(new_n663), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT51), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n656), .A2(new_n552), .A3(new_n629), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(G1336gat));
  OAI21_X1  g544(.A(G92gat), .B1(new_n740), .B2(new_n416), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n636), .A2(new_n553), .A3(new_n629), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n746), .B(new_n747), .C1(new_n743), .C2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n743), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n748), .B(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(new_n746), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n749), .B1(new_n753), .B2(new_n747), .ZN(G1337gat));
  OAI21_X1  g553(.A(G99gat), .B1(new_n740), .B2(new_n644), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n462), .A2(G99gat), .A3(new_n651), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n743), .B2(new_n756), .ZN(G1338gat));
  OAI21_X1  g556(.A(G106gat), .B1(new_n740), .B2(new_n411), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT53), .B1(new_n758), .B2(KEYINPUT110), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n411), .A2(new_n651), .A3(G106gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n743), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n759), .B(new_n761), .Z(G1339gat));
  OR3_X1    g561(.A1(new_n614), .A2(new_n616), .A3(new_n610), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(KEYINPUT54), .A3(new_n617), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n765));
  NAND3_X1  g564(.A1(new_n625), .A2(new_n627), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n767));
  INV_X1    g566(.A(new_n622), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  OAI211_X1 g569(.A(KEYINPUT55), .B(new_n764), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n623), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(KEYINPUT113), .A3(new_n623), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n764), .B1(new_n769), .B2(new_n770), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n774), .A2(new_n662), .A3(new_n775), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n531), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n527), .A2(new_n529), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n478), .B1(new_n527), .B2(new_n515), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n537), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n629), .A3(new_n542), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n588), .B1(new_n779), .B2(new_n785), .ZN(new_n786));
  AND4_X1   g585(.A1(new_n542), .A2(new_n585), .A3(new_n586), .A4(new_n784), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(new_n774), .A3(new_n775), .A4(new_n778), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n609), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n712), .A2(new_n651), .A3(new_n663), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n430), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND4_X1   g591(.A1(new_n416), .A2(new_n792), .A3(new_n411), .A4(new_n472), .ZN(new_n793));
  AOI21_X1  g592(.A(G113gat), .B1(new_n793), .B2(new_n662), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n790), .A2(new_n791), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT114), .B1(new_n795), .B2(new_n411), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n797), .B(new_n439), .C1(new_n790), .C2(new_n791), .ZN(new_n798));
  OR2_X1    g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n416), .A2(new_n656), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n462), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n544), .A2(new_n318), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n794), .B1(new_n802), .B2(new_n803), .ZN(G1340gat));
  NAND3_X1  g603(.A1(new_n793), .A2(new_n320), .A3(new_n629), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n629), .B(new_n801), .C1(new_n796), .C2(new_n798), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n807), .B2(new_n320), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT115), .ZN(G1341gat));
  AOI21_X1  g608(.A(new_n325), .B1(new_n802), .B2(new_n738), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n793), .A2(new_n325), .A3(new_n738), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n810), .A2(new_n811), .ZN(G1342gat));
  NAND3_X1  g611(.A1(new_n793), .A2(new_n323), .A3(new_n588), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT56), .Z(new_n814));
  NAND2_X1  g613(.A1(new_n802), .A2(new_n588), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n323), .ZN(G1343gat));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n643), .A2(new_n411), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n416), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n544), .A2(G141gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n792), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT119), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n792), .A2(new_n826), .A3(new_n822), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n643), .A2(new_n800), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n795), .B2(new_n439), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n439), .A2(KEYINPUT57), .ZN(new_n832));
  XOR2_X1   g631(.A(new_n785), .B(KEYINPUT116), .Z(new_n833));
  NAND4_X1  g632(.A1(new_n778), .A2(new_n543), .A3(new_n623), .A4(new_n771), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n588), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n788), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n609), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n832), .B1(new_n839), .B2(new_n791), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n662), .B(new_n830), .C1(new_n831), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(G141gat), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n818), .B1(new_n829), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n818), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n543), .B(new_n830), .C1(new_n831), .C2(new_n840), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(G141gat), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT120), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n846), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n828), .B1(G141gat), .B2(new_n841), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n848), .B(new_n849), .C1(new_n850), .C2(new_n818), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(G1344gat));
  AND2_X1   g651(.A1(new_n792), .A2(new_n822), .ZN(new_n853));
  INV_X1    g652(.A(G148gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n629), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT121), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT59), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n795), .A2(KEYINPUT57), .A3(new_n439), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n789), .A2(new_n835), .A3(KEYINPUT122), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT122), .B1(new_n789), .B2(new_n835), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n609), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n630), .A2(new_n544), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n411), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n858), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n629), .A3(new_n830), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n857), .B1(new_n865), .B2(G148gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n830), .B1(new_n831), .B2(new_n840), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n867), .A2(new_n651), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(KEYINPUT59), .A3(new_n854), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n856), .B1(new_n866), .B2(new_n869), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n738), .A2(G155gat), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT123), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(G155gat), .B1(new_n853), .B2(new_n738), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n867), .B2(new_n587), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n853), .A2(new_n311), .A3(new_n588), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NOR3_X1   g677(.A1(new_n462), .A2(new_n416), .A3(new_n656), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n795), .A2(new_n411), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n880), .A2(new_n245), .A3(new_n246), .A4(new_n662), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n799), .A2(new_n543), .A3(new_n879), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n883), .B2(new_n226), .ZN(G1348gat));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n227), .A3(new_n629), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n799), .A2(new_n629), .A3(new_n879), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n227), .ZN(G1349gat));
  OAI211_X1 g687(.A(new_n738), .B(new_n879), .C1(new_n796), .C2(new_n798), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n738), .A2(new_n216), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n889), .A2(G183gat), .B1(new_n880), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT60), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(KEYINPUT60), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n892), .A2(KEYINPUT60), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n893), .A2(new_n896), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n219), .A3(new_n588), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n588), .B(new_n879), .C1(new_n796), .C2(new_n798), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n899), .A2(new_n900), .A3(G190gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n899), .B2(G190gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT125), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g704(.A(KEYINPUT125), .B(new_n898), .C1(new_n901), .C2(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1351gat));
  XOR2_X1   g706(.A(KEYINPUT126), .B(G197gat), .Z(new_n908));
  NOR3_X1   g707(.A1(new_n643), .A2(new_n656), .A3(new_n416), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n864), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n910), .B2(new_n544), .ZN(new_n911));
  NOR4_X1   g710(.A1(new_n643), .A2(new_n656), .A3(new_n416), .A4(new_n411), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n795), .A2(new_n912), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n663), .A2(new_n908), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1352gat));
  OAI21_X1  g714(.A(G204gat), .B1(new_n910), .B2(new_n651), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n913), .A2(G204gat), .A3(new_n651), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1353gat));
  OR3_X1    g718(.A1(new_n913), .A2(G211gat), .A3(new_n609), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n864), .A2(new_n738), .A3(new_n909), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n921), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT63), .B1(new_n921), .B2(G211gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1354gat));
  INV_X1    g723(.A(new_n913), .ZN(new_n925));
  AOI21_X1  g724(.A(G218gat), .B1(new_n925), .B2(new_n588), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n910), .A2(KEYINPUT127), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n588), .A2(new_n202), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n910), .A2(KEYINPUT127), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(G1355gat));
endmodule


