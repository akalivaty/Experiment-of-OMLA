//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n548, new_n549, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(KEYINPUT65), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(KEYINPUT65), .B2(new_n459), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n472), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n468), .B1(new_n475), .B2(G2105), .ZN(G160));
  NOR2_X1   g051(.A1(new_n469), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT67), .Z(new_n479));
  OAI21_X1  g054(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n483));
  INV_X1    g058(.A(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n479), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  XNOR2_X1  g070(.A(KEYINPUT69), .B(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n462), .A2(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n469), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT69), .A2(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n487), .A2(G138), .A3(new_n462), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n502));
  OR2_X1    g077(.A1(G102), .A2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G2105), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n503), .A2(new_n505), .A3(G2104), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n517), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n515), .B2(new_n525), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT5), .B(G543), .Z(new_n527));
  NAND2_X1  g102(.A1(new_n512), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(new_n513), .ZN(new_n532));
  INV_X1    g107(.A(new_n515), .ZN(new_n533));
  AOI22_X1  g108(.A1(G90), .A2(new_n532), .B1(new_n533), .B2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n519), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT70), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n519), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n532), .A2(G81), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT71), .B(G43), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n513), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT73), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(G91), .A3(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n519), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT72), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n512), .A2(G543), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G168), .ZN(G286));
  NOR2_X1   g139(.A1(new_n511), .A2(G74), .ZN(new_n565));
  INV_X1    g140(.A(G49), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n519), .B1(new_n515), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n552), .A2(new_n553), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G87), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n568), .A2(KEYINPUT74), .A3(G87), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI211_X1 g150(.A(KEYINPUT75), .B(new_n567), .C1(new_n571), .C2(new_n572), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n568), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n527), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n533), .B2(G48), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(G305));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n513), .A2(new_n586), .B1(new_n515), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n519), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(new_n568), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n519), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n598), .A2(new_n599), .B1(G54), .B2(new_n533), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  MUX2_X1   g177(.A(G301), .B(new_n601), .S(new_n602), .Z(G284));
  MUX2_X1   g178(.A(G301), .B(new_n601), .S(new_n602), .Z(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(new_n601), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NOR2_X1   g186(.A1(new_n544), .A2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n610), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT78), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n612), .B1(new_n614), .B2(G868), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g191(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XOR2_X1   g193(.A(KEYINPUT79), .B(KEYINPUT13), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n477), .A2(G135), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n622), .A2(KEYINPUT80), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(KEYINPUT80), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G111), .B2(new_n462), .ZN(new_n625));
  INV_X1    g200(.A(G123), .ZN(new_n626));
  OAI221_X1 g201(.A(new_n621), .B1(new_n623), .B2(new_n625), .C1(new_n489), .C2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n620), .A2(G2100), .B1(new_n627), .B2(G2096), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n628), .B(new_n629), .C1(G2100), .C2(new_n620), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT81), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  INV_X1    g230(.A(new_n648), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n655), .B1(new_n651), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n662), .A2(new_n667), .A3(new_n665), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n667), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n670));
  AOI211_X1 g245(.A(new_n666), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n669), .B2(new_n670), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1981), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G5), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G171), .B2(new_n679), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(G1961), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G34), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(G29), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G160), .B2(G29), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G32), .ZN(new_n688));
  INV_X1    g263(.A(G129), .ZN(new_n689));
  OAI21_X1  g264(.A(KEYINPUT91), .B1(new_n489), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT91), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n482), .A2(new_n488), .A3(new_n691), .A4(G129), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n477), .A2(G141), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  NAND3_X1  g271(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n698), .B1(new_n690), .B2(new_n692), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(KEYINPUT92), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n688), .B1(new_n706), .B2(new_n687), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT93), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  OAI221_X1 g284(.A(new_n682), .B1(G2084), .B2(new_n686), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n609), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G4), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n687), .A2(G26), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n482), .A2(new_n488), .A3(G128), .ZN(new_n720));
  OAI211_X1 g295(.A(G140), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(KEYINPUT88), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT88), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n487), .A2(new_n723), .A3(G140), .A4(new_n462), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(G104), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n720), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n719), .B1(new_n728), .B2(new_n687), .ZN(new_n729));
  INV_X1    g304(.A(G2067), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n717), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G19), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n545), .B2(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n679), .A2(G21), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G168), .B2(new_n679), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT94), .B(G1966), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n734), .A2(G1341), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n736), .B2(new_n738), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n681), .B2(G1961), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n687), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n687), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT29), .B(G2090), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n686), .A2(G2084), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n687), .A2(G33), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n748));
  NAND3_X1  g323(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n477), .A2(G139), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n487), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(new_n462), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n747), .B1(new_n755), .B2(new_n687), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G2072), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n687), .A2(G27), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n687), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2078), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(G2078), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n756), .A2(G2072), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n757), .A2(new_n760), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT30), .B(G28), .ZN(new_n764));
  OR2_X1    g339(.A1(KEYINPUT31), .A2(G11), .ZN(new_n765));
  NAND2_X1  g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n764), .A2(new_n687), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI221_X1 g342(.A(new_n767), .B1(new_n687), .B2(new_n627), .C1(new_n734), .C2(G1341), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n763), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n741), .A2(new_n745), .A3(new_n746), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n679), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n606), .B2(new_n679), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n715), .A2(new_n716), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n732), .A2(new_n770), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n711), .A2(new_n712), .A3(new_n713), .A4(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G6), .B(G305), .S(G16), .Z(new_n778));
  XOR2_X1   g353(.A(KEYINPUT32), .B(G1981), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n679), .A2(G23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n573), .B2(new_n679), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT33), .B(G1976), .Z(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n679), .A2(G22), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G166), .B2(new_n679), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G1971), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n782), .B2(new_n783), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n780), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT34), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n780), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n591), .A2(KEYINPUT87), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n591), .A2(KEYINPUT87), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n794), .A2(G16), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n679), .A2(G24), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT86), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1986), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n687), .A2(G25), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n490), .A2(G119), .ZN(new_n802));
  OAI21_X1  g377(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(G107), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n477), .B2(G131), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n801), .B1(new_n808), .B2(new_n687), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT35), .B(G1991), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT85), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n809), .B(new_n811), .Z(new_n812));
  NOR2_X1   g387(.A1(new_n800), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n791), .A2(new_n793), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT36), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n791), .A2(new_n816), .A3(new_n793), .A4(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n777), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n777), .B2(new_n818), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n820), .A2(new_n821), .ZN(G311));
  NAND2_X1  g397(.A1(new_n777), .A2(new_n818), .ZN(G150));
  NOR2_X1   g398(.A1(new_n601), .A2(new_n610), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n527), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n519), .B1(new_n829), .B2(KEYINPUT98), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(KEYINPUT98), .B2(new_n829), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT99), .B(G55), .ZN(new_n832));
  AOI22_X1  g407(.A1(G93), .A2(new_n532), .B1(new_n533), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n545), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n826), .B(new_n835), .Z(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n837), .A2(new_n838), .A3(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n834), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT37), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n839), .A2(new_n841), .ZN(G145));
  XOR2_X1   g417(.A(new_n627), .B(G160), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n494), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n502), .A2(new_n845), .A3(new_n506), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n502), .B2(new_n506), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n501), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n728), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n507), .A2(KEYINPUT100), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n502), .A2(new_n845), .A3(new_n506), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n850), .A2(new_n851), .B1(new_n498), .B2(new_n500), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n720), .A2(new_n725), .A3(new_n727), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n849), .A2(new_n854), .A3(KEYINPUT101), .ZN(new_n855));
  AOI21_X1  g430(.A(KEYINPUT101), .B1(new_n849), .B2(new_n854), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n700), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n858));
  INV_X1    g433(.A(new_n854), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n852), .A2(new_n853), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n849), .A2(new_n854), .A3(KEYINPUT101), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(new_n703), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n755), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n857), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n700), .A2(new_n701), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n703), .A2(KEYINPUT92), .ZN(new_n867));
  OAI22_X1  g442(.A1(new_n866), .A2(new_n867), .B1(new_n860), .B2(new_n859), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n702), .A2(new_n704), .A3(new_n849), .A4(new_n854), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n755), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n477), .A2(G142), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT102), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n490), .A2(G130), .ZN(new_n873));
  OR2_X1    g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n874), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n865), .A2(new_n870), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n865), .B2(new_n870), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n618), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n865), .A2(new_n870), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n876), .ZN(new_n882));
  INV_X1    g457(.A(new_n618), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n865), .A2(new_n870), .A3(new_n877), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n880), .A2(new_n885), .A3(new_n808), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n808), .B1(new_n880), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n844), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n878), .A2(new_n879), .A3(new_n618), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n883), .B1(new_n882), .B2(new_n884), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n807), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n844), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n880), .A2(new_n885), .A3(new_n808), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n888), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n888), .A2(new_n894), .A3(KEYINPUT103), .A4(new_n895), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n898), .A2(KEYINPUT40), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT40), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(G395));
  XNOR2_X1  g477(.A(new_n835), .B(KEYINPUT104), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n614), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT78), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n613), .B(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n601), .B(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n601), .B(new_n606), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n910), .A2(KEYINPUT41), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n912), .A2(KEYINPUT105), .A3(new_n913), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n904), .A3(new_n908), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  XNOR2_X1  g497(.A(G305), .B(G303), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n573), .B(new_n591), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n911), .A2(new_n920), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n922), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n930), .B1(new_n922), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n834), .A2(new_n602), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(G331));
  XNOR2_X1  g513(.A(G171), .B(new_n835), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G286), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n835), .B(G301), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(G168), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n917), .A2(new_n943), .A3(new_n918), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n942), .A3(new_n912), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n946), .B2(new_n930), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(new_n929), .A3(new_n928), .A4(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n940), .A2(new_n942), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n914), .A2(new_n915), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n930), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n949), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n951), .B1(new_n956), .B2(KEYINPUT43), .ZN(new_n957));
  AOI211_X1 g532(.A(KEYINPUT108), .B(new_n948), .C1(new_n955), .C2(new_n949), .ZN(new_n958));
  OAI211_X1 g533(.A(KEYINPUT44), .B(new_n950), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n948), .B1(new_n947), .B2(new_n949), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n955), .A2(new_n948), .A3(new_n949), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(G397));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n848), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G40), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n967), .B(new_n468), .C1(new_n475), .C2(G2105), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n970), .A2(G1986), .A3(G290), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT109), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n728), .A2(new_n730), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n853), .A2(G2067), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(G1996), .B2(new_n700), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n705), .B2(G1996), .ZN(new_n979));
  XOR2_X1   g554(.A(new_n807), .B(new_n811), .Z(new_n980));
  OAI21_X1  g555(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n470), .B1(new_n485), .B2(new_n486), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n474), .B1(new_n983), .B2(new_n472), .ZN(new_n984));
  INV_X1    g559(.A(new_n473), .ZN(new_n985));
  OAI21_X1  g560(.A(G2105), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n468), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(G40), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT114), .B1(new_n966), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n850), .A2(new_n851), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n501), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n968), .B(new_n990), .C1(new_n992), .C2(KEYINPUT45), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n737), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n501), .B2(new_n508), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n848), .A2(new_n965), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1002));
  OAI221_X1 g577(.A(new_n968), .B1(new_n999), .B2(new_n1000), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(G2084), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n995), .A2(KEYINPUT115), .A3(new_n737), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n998), .A2(G168), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(new_n994), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n988), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(new_n1011), .B2(new_n990), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n738), .B1(new_n1012), .B2(new_n989), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1004), .B1(new_n1013), .B2(KEYINPUT115), .ZN(new_n1014));
  AOI21_X1  g589(.A(G168), .B1(new_n1014), .B2(new_n998), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT51), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT62), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1007), .A2(new_n1018), .A3(G8), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1022));
  OAI211_X1 g597(.A(G160), .B(G40), .C1(new_n1000), .C2(KEYINPUT45), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT110), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n992), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G1971), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1003), .A2(G2090), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G303), .A2(G8), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT55), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1001), .A2(new_n988), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n571), .A2(new_n572), .ZN(new_n1037));
  INV_X1    g612(.A(new_n567), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1976), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT52), .ZN(new_n1042));
  INV_X1    g617(.A(G86), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n582), .B1(new_n1043), .B2(new_n513), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G1981), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(G1981), .B2(new_n583), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1045), .B(KEYINPUT49), .C1(G1981), .C2(new_n583), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1036), .A3(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT112), .B(G1976), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n575), .A2(new_n576), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(new_n1036), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1042), .B(new_n1050), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1032), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n988), .B1(new_n999), .B2(new_n1000), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1027), .A2(G1971), .B1(new_n1059), .B2(G2090), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1056), .B1(new_n1060), .B2(G8), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1033), .A2(new_n1055), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2078), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1027), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1065));
  INV_X1    g640(.A(G1961), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1064), .A2(new_n1065), .B1(new_n1066), .B2(new_n1003), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1012), .A2(KEYINPUT53), .A3(new_n1063), .A4(new_n989), .ZN(new_n1068));
  AOI21_X1  g643(.A(G301), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1062), .A2(new_n1069), .ZN(new_n1070));
  NOR4_X1   g645(.A1(new_n1021), .A2(new_n1022), .A3(KEYINPUT126), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT126), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(KEYINPUT62), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(new_n1074), .B2(new_n1020), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n583), .A2(G1981), .ZN(new_n1077));
  NOR2_X1   g652(.A1(G288), .A2(G1976), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1077), .B1(new_n1078), .B2(new_n1050), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1079), .A2(KEYINPUT113), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1036), .B1(new_n1079), .B2(KEYINPUT113), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1033), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1080), .A2(new_n1081), .B1(new_n1082), .B2(new_n1055), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1014), .A2(new_n998), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G286), .A2(new_n1035), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1062), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1033), .A2(new_n1055), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1093), .B(new_n1094), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1083), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1027), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n557), .A2(KEYINPUT117), .ZN(new_n1099));
  INV_X1    g674(.A(new_n562), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n554), .B2(new_n556), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n562), .A2(new_n554), .A3(new_n556), .A4(KEYINPUT57), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT118), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1104), .A2(KEYINPUT118), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1103), .A2(KEYINPUT57), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1956), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1098), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1003), .A2(new_n716), .B1(new_n730), .B2(new_n1034), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1113), .A2(new_n601), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1102), .A2(new_n1100), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(KEYINPUT117), .B2(new_n557), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1104), .A2(KEYINPUT118), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1116), .A2(new_n1117), .B1(new_n1118), .B2(new_n1105), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1097), .ZN(new_n1120));
  AOI211_X1 g695(.A(new_n1120), .B(new_n1023), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1119), .B1(new_n1121), .B2(new_n1109), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1112), .B1(new_n1114), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1113), .A2(KEYINPUT60), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1124), .B(new_n601), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1113), .A2(KEYINPUT60), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT61), .B1(new_n1122), .B2(new_n1111), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT119), .B(G1996), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1027), .A2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(KEYINPUT58), .B(G1341), .Z(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n1001), .B2(new_n988), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT120), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n545), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1136), .B(new_n545), .C1(new_n1130), .C2(new_n1133), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1128), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1122), .A2(new_n1111), .A3(KEYINPUT61), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT121), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1122), .A2(new_n1111), .A3(new_n1141), .A4(KEYINPUT61), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1138), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1127), .B1(new_n1144), .B2(KEYINPUT122), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1138), .A2(new_n1143), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1123), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n968), .B(KEYINPUT124), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT53), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT125), .B(G2078), .Z(new_n1153));
  NOR3_X1   g728(.A1(new_n966), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1150), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1067), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(G171), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1149), .B1(new_n1157), .B2(new_n1069), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(G171), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1067), .A2(new_n1068), .A3(G301), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(KEYINPUT54), .A3(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1073), .A2(new_n1062), .A3(new_n1158), .A4(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1096), .B1(new_n1148), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n982), .B1(new_n1076), .B2(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n969), .A2(G1996), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT46), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT127), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n970), .B1(new_n700), .B2(new_n977), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT47), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n972), .B(KEYINPUT48), .Z(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n981), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n808), .A2(new_n811), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n975), .B1(new_n979), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n970), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1164), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g755(.A(G227), .ZN(new_n1182));
  NAND2_X1  g756(.A1(new_n1182), .A2(G319), .ZN(new_n1183));
  NOR3_X1   g757(.A1(G229), .A2(G401), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g758(.A(new_n1184), .B1(new_n961), .B2(new_n962), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1185), .B1(new_n898), .B2(new_n899), .ZN(G308));
  NAND2_X1  g760(.A1(new_n898), .A2(new_n899), .ZN(new_n1187));
  OAI211_X1 g761(.A(new_n1187), .B(new_n1184), .C1(new_n961), .C2(new_n962), .ZN(G225));
endmodule


