//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G169gat), .ZN(new_n205));
  INV_X1    g004(.A(G176gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT23), .ZN(new_n207));
  NAND3_X1  g006(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT25), .B1(new_n211), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n207), .A2(KEYINPUT66), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT23), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT25), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  AND2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(KEYINPUT24), .ZN(new_n227));
  NAND2_X1  g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n210), .A2(KEYINPUT65), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n224), .A2(new_n234), .A3(new_n212), .A4(new_n216), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  INV_X1    g035(.A(G190gat), .ZN(new_n237));
  AND2_X1   g036(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n236), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n238), .B2(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT27), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(KEYINPUT68), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(G190gat), .B1(new_n242), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n228), .B(new_n240), .C1(new_n248), .C2(new_n236), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n221), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n212), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n219), .B(new_n235), .C1(new_n249), .C2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT29), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n204), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT75), .ZN(new_n258));
  INV_X1    g057(.A(G197gat), .ZN(new_n259));
  INV_X1    g058(.A(G204gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT74), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n265), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G211gat), .B(G218gat), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT22), .ZN(new_n270));
  INV_X1    g069(.A(G211gat), .ZN(new_n271));
  INV_X1    g070(.A(G218gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n267), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n270), .B1(new_n264), .B2(new_n266), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(new_n269), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n258), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n264), .A2(new_n266), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n268), .B1(new_n279), .B2(new_n270), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(KEYINPUT75), .A3(new_n274), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n235), .A2(new_n219), .ZN(new_n283));
  NOR3_X1   g082(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT68), .B1(new_n245), .B2(new_n246), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n237), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT28), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n287), .A2(new_n228), .A3(new_n240), .A4(new_n253), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n203), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n257), .A2(new_n282), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n255), .A2(new_n256), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n203), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n255), .A2(KEYINPUT76), .A3(new_n204), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT76), .B1(new_n255), .B2(new_n204), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n290), .B1(new_n295), .B2(new_n282), .ZN(new_n296));
  XOR2_X1   g095(.A(G8gat), .B(G36gat), .Z(new_n297));
  XNOR2_X1  g096(.A(new_n297), .B(G64gat), .ZN(new_n298));
  INV_X1    g097(.A(G92gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n202), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n282), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n255), .A2(new_n204), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n292), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT76), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n255), .A2(KEYINPUT76), .A3(new_n204), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n257), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n304), .B1(new_n308), .B2(new_n302), .ZN(new_n309));
  INV_X1    g108(.A(new_n300), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(KEYINPUT77), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n301), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n300), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n309), .A2(KEYINPUT30), .A3(new_n310), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G127gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n321));
  AND2_X1   g120(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n320), .B(new_n321), .C1(new_n324), .C2(new_n317), .ZN(new_n325));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n326), .A2(KEYINPUT1), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n317), .A2(G127gat), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n326), .A2(KEYINPUT1), .A3(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n325), .A2(new_n327), .B1(new_n329), .B2(new_n318), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G141gat), .B(G148gat), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n336), .B(KEYINPUT78), .C1(KEYINPUT2), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n339));
  INV_X1    g138(.A(G141gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G148gat), .ZN(new_n341));
  INV_X1    g140(.A(G148gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G141gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT2), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n339), .B1(new_n344), .B2(new_n335), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT79), .B(G148gat), .Z(new_n347));
  OAI21_X1  g146(.A(new_n341), .B1(new_n347), .B2(new_n340), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n334), .B1(new_n333), .B2(KEYINPUT2), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n330), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n338), .A2(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT3), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n354), .B1(new_n353), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n330), .ZN(new_n359));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n353), .A2(new_n364), .A3(new_n330), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n330), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n359), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n361), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(KEYINPUT5), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n361), .A2(KEYINPUT5), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n366), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(G85gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G1gat), .B(G29gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n360), .B1(new_n358), .B2(new_n366), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT39), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n370), .A2(new_n361), .ZN(new_n384));
  OR3_X1    g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n385), .A2(KEYINPUT40), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT40), .B1(new_n385), .B2(new_n386), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n316), .A2(new_n381), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT31), .B(G50gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G228gat), .ZN(new_n393));
  INV_X1    g192(.A(G233gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n280), .B2(new_n274), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n351), .B(new_n395), .C1(new_n396), .C2(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n393), .B2(new_n394), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT80), .B1(new_n351), .B2(KEYINPUT3), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT29), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n397), .B(new_n398), .C1(new_n401), .C2(new_n282), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n282), .ZN(new_n403));
  OR3_X1    g202(.A1(new_n276), .A2(KEYINPUT82), .A3(new_n269), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT82), .B1(new_n276), .B2(new_n269), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n274), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n256), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n355), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n403), .A2(KEYINPUT83), .B1(new_n351), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n392), .B(new_n402), .C1(new_n409), .C2(new_n395), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n351), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n256), .B1(new_n356), .B2(new_n357), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(new_n302), .A3(KEYINPUT83), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n395), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n402), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n391), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G78gat), .B(G106gat), .Z(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G22gat), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n410), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n410), .B2(new_n416), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n390), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n372), .A2(new_n379), .A3(new_n374), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n372), .A2(KEYINPUT81), .A3(new_n379), .A4(new_n374), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n425), .A2(new_n381), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT38), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n300), .C1(new_n296), .C2(KEYINPUT37), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT37), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n302), .B1(new_n292), .B2(new_n303), .ZN(new_n434));
  AOI211_X1 g233(.A(new_n433), .B(new_n434), .C1(new_n302), .C2(new_n308), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n301), .B(new_n311), .C1(new_n432), .C2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n310), .B1(new_n309), .B2(new_n433), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n296), .A2(KEYINPUT37), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n431), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n430), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT84), .B1(new_n422), .B2(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n428), .A2(new_n429), .ZN(new_n442));
  INV_X1    g241(.A(new_n436), .ZN(new_n443));
  INV_X1    g242(.A(new_n439), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n421), .A4(new_n390), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n316), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n421), .B1(new_n430), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT36), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n249), .A2(new_n254), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n235), .A2(new_n219), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n283), .A2(new_n288), .A3(KEYINPUT71), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n368), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT64), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n255), .A2(new_n453), .A3(new_n330), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT72), .B(G71gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(G99gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G43gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT33), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n462), .A2(KEYINPUT32), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT73), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT73), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n462), .A2(new_n470), .A3(KEYINPUT32), .A4(new_n467), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT33), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n462), .B1(KEYINPUT32), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n466), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n473), .B1(new_n472), .B2(new_n476), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n461), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n460), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n477), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n472), .A2(new_n476), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT34), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n452), .B1(new_n483), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n482), .B1(new_n477), .B2(new_n478), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n481), .A3(new_n486), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT36), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n448), .A2(new_n451), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT86), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n483), .A2(new_n487), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n449), .A2(new_n421), .A3(new_n430), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT35), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n489), .A2(new_n490), .A3(new_n497), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n449), .A2(new_n421), .A3(new_n430), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT35), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n493), .A2(new_n494), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n494), .B1(new_n493), .B2(new_n503), .ZN(new_n505));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n508), .B(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT12), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT89), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(G50gat), .ZN(new_n519));
  INV_X1    g318(.A(G50gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(G43gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n517), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n522), .A3(KEYINPUT15), .ZN(new_n523));
  NAND2_X1  g322(.A1(G29gat), .A2(G36gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT90), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g326(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n523), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n515), .A2(KEYINPUT15), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n514), .B(new_n530), .C1(new_n532), .C2(new_n529), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n523), .B2(new_n531), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n523), .A2(new_n529), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT17), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT16), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(G1gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G1gat), .B2(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G8gat), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n539), .B(new_n542), .C1(G1gat), .C2(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n533), .A2(new_n536), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n534), .A2(new_n535), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n544), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT18), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n546), .A2(KEYINPUT18), .A3(new_n547), .A4(new_n549), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n547), .B(KEYINPUT13), .Z(new_n554));
  AND2_X1   g353(.A1(new_n548), .A2(new_n544), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n548), .A2(new_n544), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n512), .B(new_n513), .C1(new_n552), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT91), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n550), .A2(new_n551), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n557), .A3(new_n553), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT91), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n562), .A2(new_n563), .A3(new_n512), .A4(new_n513), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(KEYINPUT92), .ZN(new_n565));
  INV_X1    g364(.A(new_n558), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n565), .A2(new_n566), .A3(new_n511), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n561), .A2(KEYINPUT92), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n560), .A2(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n504), .A2(new_n505), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n571));
  XOR2_X1   g370(.A(G57gat), .B(G64gat), .Z(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  INV_X1    g372(.A(G71gat), .ZN(new_n574));
  INV_X1    g373(.A(G78gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n579), .A2(KEYINPUT21), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(KEYINPUT21), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n545), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G183gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n545), .A2(new_n584), .A3(new_n244), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n591));
  INV_X1    g390(.A(G231gat), .ZN(new_n592));
  OAI22_X1  g391(.A1(new_n590), .A2(new_n591), .B1(new_n592), .B2(new_n394), .ZN(new_n593));
  INV_X1    g392(.A(new_n591), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n592), .A2(new_n394), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n595), .A3(new_n589), .ZN(new_n596));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n271), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n593), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n599), .B1(new_n593), .B2(new_n596), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n583), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n596), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(new_n598), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n593), .A2(new_n596), .A3(new_n599), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(new_n582), .A3(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  OAI21_X1  g408(.A(KEYINPUT94), .B1(new_n609), .B2(new_n299), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT94), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n612), .A3(KEYINPUT7), .ZN(new_n613));
  NAND2_X1  g412(.A1(G99gat), .A2(G106gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(KEYINPUT8), .A2(new_n614), .B1(new_n609), .B2(new_n299), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT7), .ZN(new_n616));
  OAI211_X1 g415(.A(KEYINPUT94), .B(new_n616), .C1(new_n609), .C2(new_n299), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G99gat), .B(G106gat), .Z(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(KEYINPUT95), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT95), .ZN(new_n622));
  INV_X1    g421(.A(new_n619), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(new_n615), .A3(new_n613), .A4(new_n617), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n533), .A2(new_n536), .A3(new_n620), .A4(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n620), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(new_n548), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n237), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n237), .B1(new_n626), .B2(new_n629), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n631), .A2(new_n272), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n629), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(G190gat), .ZN(new_n635));
  AOI21_X1  g434(.A(G218gat), .B1(new_n635), .B2(new_n630), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT96), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n272), .B1(new_n631), .B2(new_n632), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n635), .A2(G218gat), .A3(new_n630), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT96), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n638), .A2(new_n646), .A3(new_n641), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n571), .B1(new_n608), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n638), .ZN(new_n650));
  INV_X1    g449(.A(new_n641), .ZN(new_n651));
  INV_X1    g450(.A(new_n646), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n642), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n607), .A3(KEYINPUT97), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT98), .Z(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n579), .A2(new_n621), .A3(new_n624), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n659), .B(new_n660), .C1(new_n628), .C2(new_n579), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n579), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n660), .B1(new_n628), .B2(new_n579), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n658), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(new_n206), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n260), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(new_n666), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n656), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n570), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n430), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT99), .B(G1gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  NAND3_X1  g479(.A1(new_n570), .A2(new_n316), .A3(new_n676), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n683), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n681), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT100), .B1(new_n683), .B2(KEYINPUT42), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n686), .B(new_n687), .C1(new_n681), .C2(new_n682), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT36), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT36), .B1(new_n489), .B2(new_n490), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT101), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n488), .A2(new_n694), .A3(new_n491), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n677), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n570), .A2(new_n495), .A3(new_n676), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n698), .B2(new_n690), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n677), .A2(new_n421), .ZN(new_n700));
  XNOR2_X1  g499(.A(KEYINPUT43), .B(G22gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT102), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n700), .B(new_n702), .ZN(G1327gat));
  AOI221_X4 g502(.A(new_n450), .B1(new_n488), .B2(new_n491), .C1(new_n441), .C2(new_n447), .ZN(new_n704));
  INV_X1    g503(.A(new_n503), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT86), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n493), .A2(new_n494), .A3(new_n503), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n560), .A2(new_n564), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n568), .A2(new_n565), .A3(new_n511), .A4(new_n566), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n607), .A2(new_n654), .A3(new_n675), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n706), .A2(new_n707), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n430), .A2(G29gat), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n712), .A2(KEYINPUT103), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT103), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n654), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n706), .A2(new_n707), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n450), .B1(new_n441), .B2(new_n447), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n696), .A2(new_n722), .B1(new_n502), .B2(new_n499), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n723), .B2(new_n654), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n607), .B(KEYINPUT104), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n674), .B(KEYINPUT105), .Z(new_n728));
  NOR3_X1   g527(.A1(new_n727), .A2(new_n569), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n725), .A2(new_n442), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G29gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n715), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n718), .A2(new_n731), .A3(new_n732), .ZN(G1328gat));
  NAND4_X1  g532(.A1(new_n721), .A2(new_n316), .A3(new_n724), .A4(new_n729), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n735), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(G36gat), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n449), .A2(G36gat), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT46), .B1(new_n712), .B2(new_n739), .ZN(new_n740));
  OR3_X1    g539(.A1(new_n712), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(G1329gat));
  INV_X1    g541(.A(new_n495), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n570), .A2(KEYINPUT107), .A3(new_n711), .A4(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746));
  INV_X1    g545(.A(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n712), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n696), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n721), .A2(new_n750), .A3(new_n724), .A4(new_n729), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1330gat));
  INV_X1    g556(.A(new_n421), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n721), .A2(new_n758), .A3(new_n724), .A4(new_n729), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G50gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n570), .A2(new_n520), .A3(new_n758), .A4(new_n711), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n760), .B2(new_n761), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n696), .A2(new_n722), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n503), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n649), .A2(new_n569), .A3(new_n655), .A4(new_n728), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n430), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(G57gat), .Z(G1332gat));
  NAND3_X1  g571(.A1(new_n767), .A2(KEYINPUT108), .A3(new_n769), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n723), .B2(new_n768), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n449), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  AND2_X1   g576(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n776), .B2(new_n777), .ZN(G1333gat));
  OAI21_X1  g579(.A(new_n574), .B1(new_n770), .B2(new_n743), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n773), .A2(new_n775), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n696), .A2(new_n574), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT109), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n785));
  INV_X1    g584(.A(new_n783), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n785), .B(new_n786), .C1(new_n773), .C2(new_n775), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n781), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT50), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n790), .B(new_n781), .C1(new_n784), .C2(new_n787), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(G1334gat));
  NAND2_X1  g591(.A1(new_n782), .A2(new_n758), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT110), .B(G78gat), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1335gat));
  NOR2_X1   g594(.A1(new_n607), .A2(new_n710), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n674), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n721), .A2(new_n442), .A3(new_n724), .A4(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(G85gat), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n654), .B1(new_n766), .B2(new_n503), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT51), .B1(new_n804), .B2(new_n796), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  NOR4_X1   g605(.A1(new_n723), .A2(new_n806), .A3(new_n654), .A4(new_n797), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n675), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n442), .A2(new_n609), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  INV_X1    g609(.A(new_n728), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n811), .A2(new_n449), .A3(G92gat), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n805), .B2(new_n807), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n723), .A2(new_n654), .A3(new_n797), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT112), .B1(new_n816), .B2(KEYINPUT51), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n813), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n721), .A2(new_n316), .A3(new_n724), .A4(new_n798), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(G92gat), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT52), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(G92gat), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n805), .A2(new_n807), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n822), .B(new_n823), .C1(new_n824), .C2(new_n813), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n821), .A2(new_n825), .ZN(G1337gat));
  NAND3_X1  g625(.A1(new_n725), .A2(new_n750), .A3(new_n798), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G99gat), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n743), .A2(G99gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n828), .B1(new_n808), .B2(new_n829), .ZN(G1338gat));
  OR3_X1    g629(.A1(new_n811), .A2(G106gat), .A3(new_n421), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT113), .Z(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n815), .B2(new_n817), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n721), .A2(new_n758), .A3(new_n724), .A4(new_n798), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(G106gat), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT53), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(G106gat), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n837), .B(new_n838), .C1(new_n824), .C2(new_n832), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(G1339gat));
  NOR3_X1   g639(.A1(new_n555), .A2(new_n556), .A3(new_n554), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n547), .B1(new_n546), .B2(new_n549), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n510), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n709), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n675), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n661), .A2(new_n658), .A3(new_n662), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT114), .B(new_n672), .C1(new_n663), .C2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n661), .A2(new_n662), .ZN(new_n851));
  INV_X1    g650(.A(new_n658), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n850), .B1(new_n853), .B2(new_n670), .ZN(new_n854));
  OAI211_X1 g653(.A(KEYINPUT55), .B(new_n847), .C1(new_n849), .C2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n673), .ZN(new_n856));
  AOI211_X1 g655(.A(KEYINPUT54), .B(new_n658), .C1(new_n661), .C2(new_n662), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT114), .B1(new_n857), .B2(new_n672), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n853), .A2(new_n850), .A3(new_n670), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n847), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT55), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n710), .A2(new_n856), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n648), .B1(new_n845), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n855), .A2(new_n673), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n863), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n654), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT115), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT55), .B1(new_n860), .B2(new_n847), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n569), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n844), .A2(new_n675), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n654), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n648), .A2(new_n844), .A3(new_n856), .A4(new_n863), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n869), .A2(new_n726), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n649), .A2(new_n569), .A3(new_n655), .A4(new_n674), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n743), .A2(new_n758), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n442), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT116), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n881), .A2(KEYINPUT116), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n449), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(new_n449), .C1(new_n883), .C2(new_n884), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n569), .A2(G113gat), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT118), .Z(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n879), .A2(new_n880), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n442), .A3(new_n449), .ZN(new_n893));
  OAI21_X1  g692(.A(G113gat), .B1(new_n893), .B2(new_n569), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(G1340gat));
  NOR2_X1   g694(.A1(new_n674), .A2(G120gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n886), .A2(new_n888), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G120gat), .B1(new_n893), .B2(new_n811), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g699(.A(KEYINPUT119), .B(G120gat), .C1(new_n893), .C2(new_n811), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(new_n902), .ZN(G1341gat));
  INV_X1    g702(.A(new_n324), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n893), .A2(new_n904), .A3(new_n726), .ZN(new_n905));
  INV_X1    g704(.A(new_n884), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n316), .B1(new_n906), .B2(new_n882), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n607), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n905), .B1(new_n908), .B2(new_n904), .ZN(G1342gat));
  OAI211_X1 g708(.A(new_n449), .B(new_n648), .C1(new_n883), .C2(new_n884), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT56), .B1(new_n910), .B2(G134gat), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n907), .A2(new_n912), .A3(new_n317), .A4(new_n648), .ZN(new_n913));
  OAI21_X1  g712(.A(G134gat), .B1(new_n893), .B2(new_n654), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(G1343gat));
  NAND2_X1  g714(.A1(new_n879), .A2(new_n758), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n430), .B(new_n316), .C1(new_n693), .C2(new_n695), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n340), .A3(new_n710), .ZN(new_n920));
  INV_X1    g719(.A(new_n878), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n871), .B2(new_n872), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n864), .A2(KEYINPUT120), .A3(new_n845), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n654), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n607), .B1(new_n925), .B2(new_n874), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n758), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT57), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n879), .A2(new_n929), .A3(new_n758), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n928), .A2(new_n930), .A3(new_n710), .A4(new_n918), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n931), .A2(G141gat), .B1(KEYINPUT121), .B2(KEYINPUT58), .ZN(new_n932));
  NOR2_X1   g731(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT122), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n920), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n920), .B2(new_n932), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1344gat));
  INV_X1    g736(.A(new_n347), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n919), .A2(new_n938), .A3(new_n675), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n918), .A2(KEYINPUT123), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n674), .B1(new_n918), .B2(KEYINPUT123), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n874), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n608), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n878), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n945), .B2(new_n758), .ZN(new_n946));
  AOI211_X1 g745(.A(new_n929), .B(new_n421), .C1(new_n877), .C2(new_n878), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n941), .B(new_n942), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n342), .B1(new_n948), .B2(KEYINPUT124), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n927), .A2(new_n929), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n950), .B1(new_n929), .B2(new_n916), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n951), .A2(new_n952), .A3(new_n941), .A4(new_n942), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n940), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n928), .A2(new_n918), .A3(new_n930), .ZN(new_n955));
  AOI211_X1 g754(.A(KEYINPUT59), .B(new_n938), .C1(new_n955), .C2(new_n675), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n939), .B1(new_n954), .B2(new_n956), .ZN(G1345gat));
  AOI21_X1  g756(.A(G155gat), .B1(new_n919), .B2(new_n607), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n955), .A2(G155gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n727), .ZN(G1346gat));
  AOI21_X1  g759(.A(G162gat), .B1(new_n919), .B2(new_n648), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n955), .A2(G162gat), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n648), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n442), .A2(new_n449), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n892), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n965), .A2(new_n569), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(new_n205), .ZN(G1348gat));
  NOR3_X1   g766(.A1(new_n965), .A2(new_n206), .A3(new_n811), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n892), .A2(new_n675), .A3(new_n964), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n968), .B1(new_n206), .B2(new_n969), .ZN(G1349gat));
  OAI21_X1  g769(.A(G183gat), .B1(new_n965), .B2(new_n726), .ZN(new_n971));
  NAND2_X1  g770(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n242), .A2(new_n247), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n892), .A2(new_n973), .A3(new_n607), .A4(new_n964), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n971), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OR2_X1    g774(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(G1350gat));
  XNOR2_X1  g776(.A(KEYINPUT61), .B(G190gat), .ZN(new_n978));
  NAND2_X1  g777(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n965), .A2(new_n654), .ZN(new_n980));
  MUX2_X1   g779(.A(new_n978), .B(new_n979), .S(new_n980), .Z(G1351gat));
  AND2_X1   g780(.A1(new_n696), .A2(new_n964), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n951), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(G197gat), .B1(new_n983), .B2(new_n569), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n917), .A2(new_n982), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(new_n259), .A3(new_n710), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n984), .A2(new_n987), .ZN(G1352gat));
  NOR3_X1   g787(.A1(new_n985), .A2(G204gat), .A3(new_n674), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(G204gat), .B1(new_n983), .B2(new_n811), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n989), .A2(new_n990), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(G1353gat));
  NAND3_X1  g793(.A1(new_n951), .A2(new_n607), .A3(new_n982), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(G211gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n996), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n986), .A2(new_n271), .A3(new_n607), .ZN(new_n998));
  NAND2_X1  g797(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n999));
  OR2_X1    g798(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1000));
  NAND4_X1  g799(.A1(new_n995), .A2(G211gat), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n997), .A2(new_n998), .A3(new_n1001), .ZN(G1354gat));
  OAI21_X1  g801(.A(G218gat), .B1(new_n983), .B2(new_n654), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n986), .A2(new_n272), .A3(new_n648), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1355gat));
endmodule


