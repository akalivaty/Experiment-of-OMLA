

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U553 ( .A(n563), .B(n562), .ZN(n894) );
  XNOR2_X1 U554 ( .A(n567), .B(n566), .ZN(G164) );
  AND2_X1 U555 ( .A1(n539), .A2(n538), .ZN(n537) );
  NAND2_X1 U556 ( .A1(n807), .A2(n522), .ZN(n538) );
  NAND2_X1 U557 ( .A1(n797), .A2(n526), .ZN(n539) );
  NAND2_X1 U558 ( .A1(n548), .A2(n546), .ZN(n752) );
  NAND2_X1 U559 ( .A1(n773), .A2(n520), .ZN(n778) );
  NAND2_X1 U560 ( .A1(n533), .A2(n523), .ZN(n532) );
  NAND2_X1 U561 ( .A1(n534), .A2(n537), .ZN(n533) );
  OR2_X1 U562 ( .A1(n540), .A2(n544), .ZN(n534) );
  XNOR2_X1 U563 ( .A(n528), .B(n527), .ZN(n786) );
  XNOR2_X1 U564 ( .A(n733), .B(KEYINPUT64), .ZN(n808) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n733) );
  XNOR2_X1 U566 ( .A(n558), .B(n556), .ZN(n555) );
  INV_X1 U567 ( .A(KEYINPUT91), .ZN(n556) );
  XNOR2_X1 U568 ( .A(n553), .B(KEYINPUT102), .ZN(n547) );
  NAND2_X1 U569 ( .A1(n746), .A2(n552), .ZN(n545) );
  OR2_X1 U570 ( .A1(n745), .A2(KEYINPUT101), .ZN(n551) );
  NAND2_X1 U571 ( .A1(n550), .A2(n554), .ZN(n549) );
  INV_X1 U572 ( .A(n746), .ZN(n550) );
  AND2_X1 U573 ( .A1(n808), .A2(n734), .ZN(n760) );
  INV_X1 U574 ( .A(KEYINPUT29), .ZN(n757) );
  NAND2_X1 U575 ( .A1(n542), .A2(n541), .ZN(n540) );
  INV_X1 U576 ( .A(n807), .ZN(n541) );
  INV_X1 U577 ( .A(n797), .ZN(n542) );
  NAND2_X1 U578 ( .A1(n529), .A2(n785), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n778), .A2(G286), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n842) );
  NAND2_X1 U581 ( .A1(n804), .A2(n518), .ZN(n530) );
  AND2_X1 U582 ( .A1(n535), .A2(n532), .ZN(n531) );
  XNOR2_X1 U583 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n563) );
  NAND2_X1 U584 ( .A1(n557), .A2(n555), .ZN(n566) );
  AND2_X1 U585 ( .A1(n565), .A2(n524), .ZN(n557) );
  AND2_X1 U586 ( .A1(n537), .A2(KEYINPUT105), .ZN(n518) );
  OR2_X1 U587 ( .A1(G299), .A2(n753), .ZN(n519) );
  XOR2_X1 U588 ( .A(n772), .B(KEYINPUT31), .Z(n520) );
  AND2_X1 U589 ( .A1(n519), .A2(n551), .ZN(n521) );
  NAND2_X1 U590 ( .A1(n803), .A2(n802), .ZN(n522) );
  OR2_X1 U591 ( .A1(n537), .A2(n544), .ZN(n523) );
  INV_X1 U592 ( .A(n804), .ZN(n543) );
  AND2_X1 U593 ( .A1(n561), .A2(n560), .ZN(n524) );
  AND2_X1 U594 ( .A1(n545), .A2(n521), .ZN(n525) );
  NAND2_X1 U595 ( .A1(n790), .A2(n789), .ZN(n526) );
  XOR2_X1 U596 ( .A(KEYINPUT32), .B(KEYINPUT104), .Z(n527) );
  INV_X1 U597 ( .A(KEYINPUT105), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n543), .A2(n536), .ZN(n535) );
  AND2_X1 U599 ( .A1(n540), .A2(n544), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n547), .A2(n519), .ZN(n546) );
  NAND2_X1 U601 ( .A1(n525), .A2(n549), .ZN(n548) );
  AND2_X1 U602 ( .A1(n745), .A2(KEYINPUT101), .ZN(n552) );
  NOR2_X1 U603 ( .A1(n747), .A2(n941), .ZN(n553) );
  INV_X1 U604 ( .A(KEYINPUT101), .ZN(n554) );
  NAND2_X1 U605 ( .A1(n894), .A2(G138), .ZN(n558) );
  XNOR2_X1 U606 ( .A(n758), .B(n757), .ZN(n763) );
  INV_X1 U607 ( .A(n760), .ZN(n779) );
  OR2_X1 U608 ( .A1(G301), .A2(n769), .ZN(n559) );
  INV_X1 U609 ( .A(n809), .ZN(n734) );
  NOR2_X1 U610 ( .A1(G2104), .A2(G2105), .ZN(n562) );
  NOR2_X1 U611 ( .A1(G651), .A2(n672), .ZN(n685) );
  NOR2_X1 U612 ( .A1(G651), .A2(G543), .ZN(n692) );
  INV_X1 U613 ( .A(KEYINPUT92), .ZN(n567) );
  INV_X1 U614 ( .A(G2105), .ZN(n564) );
  AND2_X1 U615 ( .A1(n564), .A2(G2104), .ZN(n893) );
  NAND2_X1 U616 ( .A1(G102), .A2(n893), .ZN(n561) );
  AND2_X1 U617 ( .A1(G2104), .A2(G2105), .ZN(n889) );
  NAND2_X1 U618 ( .A1(G114), .A2(n889), .ZN(n560) );
  NOR2_X1 U619 ( .A1(G2104), .A2(n564), .ZN(n890) );
  NAND2_X1 U620 ( .A1(n890), .A2(G126), .ZN(n565) );
  XNOR2_X1 U621 ( .A(G2446), .B(KEYINPUT106), .ZN(n577) );
  XOR2_X1 U622 ( .A(G2430), .B(G2427), .Z(n569) );
  XNOR2_X1 U623 ( .A(G2435), .B(G2438), .ZN(n568) );
  XNOR2_X1 U624 ( .A(n569), .B(n568), .ZN(n573) );
  XOR2_X1 U625 ( .A(G2454), .B(KEYINPUT107), .Z(n571) );
  XNOR2_X1 U626 ( .A(G1348), .B(G1341), .ZN(n570) );
  XNOR2_X1 U627 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U628 ( .A(n573), .B(n572), .Z(n575) );
  XNOR2_X1 U629 ( .A(G2443), .B(G2451), .ZN(n574) );
  XNOR2_X1 U630 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U631 ( .A(n577), .B(n576), .ZN(n578) );
  AND2_X1 U632 ( .A1(n578), .A2(G14), .ZN(G401) );
  AND2_X1 U633 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U634 ( .A(G132), .ZN(G219) );
  INV_X1 U635 ( .A(G69), .ZN(G235) );
  INV_X1 U636 ( .A(G651), .ZN(n582) );
  NOR2_X1 U637 ( .A1(G543), .A2(n582), .ZN(n579) );
  XOR2_X1 U638 ( .A(KEYINPUT1), .B(n579), .Z(n684) );
  NAND2_X1 U639 ( .A1(G64), .A2(n684), .ZN(n581) );
  XOR2_X1 U640 ( .A(KEYINPUT0), .B(G543), .Z(n672) );
  NAND2_X1 U641 ( .A1(G52), .A2(n685), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n587) );
  NOR2_X1 U643 ( .A1(n672), .A2(n582), .ZN(n688) );
  NAND2_X1 U644 ( .A1(G77), .A2(n688), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G90), .A2(n692), .ZN(n583) );
  NAND2_X1 U646 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT9), .B(n585), .Z(n586) );
  NOR2_X1 U648 ( .A1(n587), .A2(n586), .ZN(G171) );
  NAND2_X1 U649 ( .A1(n684), .A2(G63), .ZN(n588) );
  XNOR2_X1 U650 ( .A(n588), .B(KEYINPUT76), .ZN(n590) );
  NAND2_X1 U651 ( .A1(G51), .A2(n685), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U653 ( .A(KEYINPUT6), .B(n591), .ZN(n599) );
  NAND2_X1 U654 ( .A1(G89), .A2(n692), .ZN(n592) );
  XNOR2_X1 U655 ( .A(n592), .B(KEYINPUT74), .ZN(n593) );
  XNOR2_X1 U656 ( .A(n593), .B(KEYINPUT4), .ZN(n595) );
  NAND2_X1 U657 ( .A1(G76), .A2(n688), .ZN(n594) );
  NAND2_X1 U658 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U659 ( .A(KEYINPUT75), .B(n596), .ZN(n597) );
  XNOR2_X1 U660 ( .A(KEYINPUT5), .B(n597), .ZN(n598) );
  NOR2_X1 U661 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U662 ( .A(KEYINPUT7), .B(n600), .Z(G168) );
  XOR2_X1 U663 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U664 ( .A1(G7), .A2(G661), .ZN(n601) );
  XNOR2_X1 U665 ( .A(n601), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U666 ( .A(G223), .ZN(n857) );
  NAND2_X1 U667 ( .A1(n857), .A2(G567), .ZN(n602) );
  XOR2_X1 U668 ( .A(KEYINPUT11), .B(n602), .Z(G234) );
  NAND2_X1 U669 ( .A1(n684), .A2(G56), .ZN(n603) );
  XOR2_X1 U670 ( .A(KEYINPUT14), .B(n603), .Z(n611) );
  NAND2_X1 U671 ( .A1(G68), .A2(n688), .ZN(n607) );
  XOR2_X1 U672 ( .A(KEYINPUT71), .B(KEYINPUT12), .Z(n605) );
  NAND2_X1 U673 ( .A1(G81), .A2(n692), .ZN(n604) );
  XNOR2_X1 U674 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U675 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U676 ( .A(n608), .B(KEYINPUT13), .ZN(n609) );
  XOR2_X1 U677 ( .A(KEYINPUT72), .B(n609), .Z(n610) );
  NOR2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n685), .A2(G43), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n944) );
  INV_X1 U681 ( .A(G860), .ZN(n634) );
  OR2_X1 U682 ( .A1(n944), .A2(n634), .ZN(G153) );
  INV_X1 U683 ( .A(G868), .ZN(n705) );
  NOR2_X1 U684 ( .A1(n705), .A2(G171), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n614), .B(KEYINPUT73), .ZN(n623) );
  NAND2_X1 U686 ( .A1(G79), .A2(n688), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G66), .A2(n684), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U689 ( .A1(G92), .A2(n692), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G54), .A2(n685), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT15), .B(n621), .Z(n941) );
  OR2_X1 U694 ( .A1(G868), .A2(n941), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(G284) );
  NAND2_X1 U696 ( .A1(G78), .A2(n688), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G65), .A2(n684), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G53), .A2(n685), .ZN(n626) );
  XNOR2_X1 U700 ( .A(KEYINPUT69), .B(n626), .ZN(n627) );
  NOR2_X1 U701 ( .A1(n628), .A2(n627), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n692), .A2(G91), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(G299) );
  XNOR2_X1 U704 ( .A(KEYINPUT77), .B(G868), .ZN(n631) );
  NOR2_X1 U705 ( .A1(G286), .A2(n631), .ZN(n633) );
  NOR2_X1 U706 ( .A1(G868), .A2(G299), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(G297) );
  NAND2_X1 U708 ( .A1(n634), .A2(G559), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n635), .A2(n941), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n636), .B(KEYINPUT16), .ZN(n638) );
  XOR2_X1 U711 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n637) );
  XNOR2_X1 U712 ( .A(n638), .B(n637), .ZN(G148) );
  NOR2_X1 U713 ( .A1(G868), .A2(n944), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G868), .A2(n941), .ZN(n639) );
  NOR2_X1 U715 ( .A1(G559), .A2(n639), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n641), .A2(n640), .ZN(G282) );
  NAND2_X1 U717 ( .A1(G99), .A2(n893), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G111), .A2(n889), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U720 ( .A(KEYINPUT80), .B(n644), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n890), .A2(G123), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT18), .B(n645), .Z(n646) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n894), .A2(G135), .ZN(n648) );
  NAND2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n992) );
  XNOR2_X1 U726 ( .A(n992), .B(G2096), .ZN(n650) );
  XNOR2_X1 U727 ( .A(n650), .B(KEYINPUT81), .ZN(n652) );
  INV_X1 U728 ( .A(G2100), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(G156) );
  NAND2_X1 U730 ( .A1(n941), .A2(G559), .ZN(n702) );
  XNOR2_X1 U731 ( .A(n944), .B(n702), .ZN(n653) );
  NOR2_X1 U732 ( .A1(n653), .A2(G860), .ZN(n660) );
  NAND2_X1 U733 ( .A1(G80), .A2(n688), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G67), .A2(n684), .ZN(n654) );
  NAND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U736 ( .A1(G93), .A2(n692), .ZN(n657) );
  NAND2_X1 U737 ( .A1(G55), .A2(n685), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n657), .A2(n656), .ZN(n658) );
  OR2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n704) );
  XOR2_X1 U740 ( .A(n660), .B(n704), .Z(G145) );
  NAND2_X1 U741 ( .A1(G62), .A2(n684), .ZN(n662) );
  NAND2_X1 U742 ( .A1(G50), .A2(n685), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U744 ( .A(KEYINPUT85), .B(n663), .ZN(n667) );
  NAND2_X1 U745 ( .A1(G75), .A2(n688), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G88), .A2(n692), .ZN(n664) );
  AND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U748 ( .A1(n667), .A2(n666), .ZN(G303) );
  INV_X1 U749 ( .A(G303), .ZN(G166) );
  NAND2_X1 U750 ( .A1(G49), .A2(n685), .ZN(n669) );
  NAND2_X1 U751 ( .A1(G74), .A2(G651), .ZN(n668) );
  NAND2_X1 U752 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U753 ( .A(KEYINPUT82), .B(n670), .ZN(n671) );
  NOR2_X1 U754 ( .A1(n684), .A2(n671), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n672), .A2(G87), .ZN(n673) );
  NAND2_X1 U756 ( .A1(n674), .A2(n673), .ZN(G288) );
  NAND2_X1 U757 ( .A1(n692), .A2(G86), .ZN(n675) );
  XOR2_X1 U758 ( .A(KEYINPUT83), .B(n675), .Z(n677) );
  NAND2_X1 U759 ( .A1(n684), .A2(G61), .ZN(n676) );
  NAND2_X1 U760 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U761 ( .A(KEYINPUT84), .B(n678), .ZN(n681) );
  NAND2_X1 U762 ( .A1(n688), .A2(G73), .ZN(n679) );
  XOR2_X1 U763 ( .A(KEYINPUT2), .B(n679), .Z(n680) );
  NOR2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U765 ( .A1(n685), .A2(G48), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n683), .A2(n682), .ZN(G305) );
  NAND2_X1 U767 ( .A1(G60), .A2(n684), .ZN(n687) );
  NAND2_X1 U768 ( .A1(G47), .A2(n685), .ZN(n686) );
  NAND2_X1 U769 ( .A1(n687), .A2(n686), .ZN(n691) );
  NAND2_X1 U770 ( .A1(G72), .A2(n688), .ZN(n689) );
  XOR2_X1 U771 ( .A(KEYINPUT68), .B(n689), .Z(n690) );
  NOR2_X1 U772 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U773 ( .A1(n692), .A2(G85), .ZN(n693) );
  NAND2_X1 U774 ( .A1(n694), .A2(n693), .ZN(G290) );
  XNOR2_X1 U775 ( .A(KEYINPUT19), .B(KEYINPUT86), .ZN(n695) );
  XOR2_X1 U776 ( .A(n695), .B(n704), .Z(n696) );
  XNOR2_X1 U777 ( .A(G166), .B(n696), .ZN(n699) );
  XOR2_X1 U778 ( .A(n944), .B(G305), .Z(n697) );
  XNOR2_X1 U779 ( .A(G288), .B(n697), .ZN(n698) );
  XNOR2_X1 U780 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U781 ( .A(n700), .B(G290), .ZN(n701) );
  XNOR2_X1 U782 ( .A(n701), .B(G299), .ZN(n906) );
  XNOR2_X1 U783 ( .A(n702), .B(n906), .ZN(n703) );
  NAND2_X1 U784 ( .A1(n703), .A2(G868), .ZN(n707) );
  NAND2_X1 U785 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U786 ( .A1(n707), .A2(n706), .ZN(G295) );
  NAND2_X1 U787 ( .A1(G2078), .A2(G2084), .ZN(n708) );
  XOR2_X1 U788 ( .A(KEYINPUT20), .B(n708), .Z(n709) );
  NAND2_X1 U789 ( .A1(G2090), .A2(n709), .ZN(n711) );
  XOR2_X1 U790 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n710) );
  XNOR2_X1 U791 ( .A(n711), .B(n710), .ZN(n712) );
  NAND2_X1 U792 ( .A1(G2072), .A2(n712), .ZN(G158) );
  XNOR2_X1 U793 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U794 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NAND2_X1 U795 ( .A1(G120), .A2(G57), .ZN(n713) );
  NOR2_X1 U796 ( .A1(G235), .A2(n713), .ZN(n714) );
  XNOR2_X1 U797 ( .A(KEYINPUT88), .B(n714), .ZN(n715) );
  NAND2_X1 U798 ( .A1(n715), .A2(G108), .ZN(n864) );
  NAND2_X1 U799 ( .A1(G567), .A2(n864), .ZN(n720) );
  NOR2_X1 U800 ( .A1(G220), .A2(G219), .ZN(n716) );
  XOR2_X1 U801 ( .A(KEYINPUT22), .B(n716), .Z(n717) );
  NOR2_X1 U802 ( .A1(G218), .A2(n717), .ZN(n718) );
  NAND2_X1 U803 ( .A1(G96), .A2(n718), .ZN(n865) );
  NAND2_X1 U804 ( .A1(G2106), .A2(n865), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U806 ( .A(KEYINPUT89), .B(n721), .ZN(G319) );
  INV_X1 U807 ( .A(G319), .ZN(n724) );
  NAND2_X1 U808 ( .A1(G661), .A2(G483), .ZN(n722) );
  XNOR2_X1 U809 ( .A(KEYINPUT90), .B(n722), .ZN(n723) );
  NOR2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n863) );
  NAND2_X1 U811 ( .A1(n863), .A2(G36), .ZN(G176) );
  XOR2_X1 U812 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n726) );
  NAND2_X1 U813 ( .A1(G101), .A2(n893), .ZN(n725) );
  XNOR2_X1 U814 ( .A(n726), .B(n725), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n889), .A2(G113), .ZN(n727) );
  NAND2_X1 U816 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U817 ( .A1(G137), .A2(n894), .ZN(n730) );
  NAND2_X1 U818 ( .A1(G125), .A2(n890), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U820 ( .A1(n732), .A2(n731), .ZN(G160) );
  INV_X1 U821 ( .A(G171), .ZN(G301) );
  NAND2_X1 U822 ( .A1(G160), .A2(G40), .ZN(n809) );
  NOR2_X1 U823 ( .A1(n779), .A2(G2084), .ZN(n735) );
  XNOR2_X1 U824 ( .A(n735), .B(KEYINPUT98), .ZN(n764) );
  NAND2_X1 U825 ( .A1(n764), .A2(G8), .ZN(n777) );
  NAND2_X1 U826 ( .A1(G8), .A2(n779), .ZN(n805) );
  NOR2_X1 U827 ( .A1(G1966), .A2(n805), .ZN(n775) );
  NAND2_X1 U828 ( .A1(n779), .A2(G1341), .ZN(n737) );
  INV_X1 U829 ( .A(n944), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n740) );
  AND2_X1 U831 ( .A1(n760), .A2(G1996), .ZN(n738) );
  XNOR2_X1 U832 ( .A(n738), .B(KEYINPUT26), .ZN(n739) );
  NOR2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n742) );
  INV_X1 U834 ( .A(KEYINPUT65), .ZN(n741) );
  XNOR2_X1 U835 ( .A(n742), .B(n741), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n747), .A2(n941), .ZN(n746) );
  NOR2_X1 U837 ( .A1(n760), .A2(G1348), .ZN(n744) );
  NOR2_X1 U838 ( .A1(G2067), .A2(n779), .ZN(n743) );
  NOR2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U840 ( .A1(n760), .A2(G2072), .ZN(n749) );
  XNOR2_X1 U841 ( .A(KEYINPUT27), .B(KEYINPUT100), .ZN(n748) );
  XNOR2_X1 U842 ( .A(n749), .B(n748), .ZN(n751) );
  NAND2_X1 U843 ( .A1(n779), .A2(G1956), .ZN(n750) );
  NAND2_X1 U844 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U845 ( .A(n752), .B(KEYINPUT103), .ZN(n756) );
  NAND2_X1 U846 ( .A1(G299), .A2(n753), .ZN(n754) );
  XNOR2_X1 U847 ( .A(KEYINPUT28), .B(n754), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U849 ( .A(G2078), .B(KEYINPUT25), .ZN(n759) );
  XNOR2_X1 U850 ( .A(n759), .B(KEYINPUT99), .ZN(n1022) );
  NOR2_X1 U851 ( .A1(n1022), .A2(n779), .ZN(n762) );
  NOR2_X1 U852 ( .A1(n760), .A2(G1961), .ZN(n761) );
  NOR2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n763), .A2(n559), .ZN(n773) );
  INV_X1 U855 ( .A(n764), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G8), .A2(n765), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n775), .A2(n766), .ZN(n767) );
  XOR2_X1 U858 ( .A(KEYINPUT30), .B(n767), .Z(n768) );
  NOR2_X1 U859 ( .A1(G168), .A2(n768), .ZN(n771) );
  AND2_X1 U860 ( .A1(G301), .A2(n769), .ZN(n770) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  INV_X1 U862 ( .A(n778), .ZN(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n787) );
  INV_X1 U865 ( .A(G8), .ZN(n784) );
  NOR2_X1 U866 ( .A1(G1971), .A2(n805), .ZN(n781) );
  NOR2_X1 U867 ( .A1(G2090), .A2(n779), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n782), .A2(G303), .ZN(n783) );
  OR2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n787), .A2(n786), .ZN(n804) );
  NOR2_X1 U872 ( .A1(G1976), .A2(G288), .ZN(n949) );
  NOR2_X1 U873 ( .A1(G1971), .A2(G303), .ZN(n788) );
  NOR2_X1 U874 ( .A1(n949), .A2(n788), .ZN(n790) );
  INV_X1 U875 ( .A(KEYINPUT33), .ZN(n789) );
  INV_X1 U876 ( .A(n805), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n951) );
  AND2_X1 U878 ( .A1(n791), .A2(n951), .ZN(n792) );
  NOR2_X1 U879 ( .A1(KEYINPUT33), .A2(n792), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n949), .A2(KEYINPUT33), .ZN(n793) );
  NOR2_X1 U881 ( .A1(n793), .A2(n805), .ZN(n794) );
  NOR2_X1 U882 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U883 ( .A(G1981), .B(G305), .Z(n937) );
  AND2_X1 U884 ( .A1(n796), .A2(n937), .ZN(n797) );
  NOR2_X1 U885 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U886 ( .A1(G8), .A2(n798), .ZN(n803) );
  NOR2_X1 U887 ( .A1(G1981), .A2(G305), .ZN(n799) );
  XNOR2_X1 U888 ( .A(n799), .B(KEYINPUT24), .ZN(n800) );
  XNOR2_X1 U889 ( .A(KEYINPUT97), .B(n800), .ZN(n801) );
  NOR2_X1 U890 ( .A1(n805), .A2(n801), .ZN(n806) );
  INV_X1 U891 ( .A(n806), .ZN(n802) );
  OR2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n943) );
  NOR2_X1 U894 ( .A1(n809), .A2(n808), .ZN(n852) );
  NAND2_X1 U895 ( .A1(n943), .A2(n852), .ZN(n840) );
  XOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .Z(n810) );
  XNOR2_X1 U897 ( .A(KEYINPUT93), .B(n810), .ZN(n843) );
  NAND2_X1 U898 ( .A1(G104), .A2(n893), .ZN(n812) );
  NAND2_X1 U899 ( .A1(G140), .A2(n894), .ZN(n811) );
  NAND2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U901 ( .A(KEYINPUT34), .B(n813), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G116), .A2(n889), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G128), .A2(n890), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U905 ( .A(KEYINPUT35), .B(n816), .Z(n817) );
  NOR2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U907 ( .A(KEYINPUT36), .B(n819), .ZN(n902) );
  NOR2_X1 U908 ( .A1(n843), .A2(n902), .ZN(n1000) );
  NAND2_X1 U909 ( .A1(n852), .A2(n1000), .ZN(n849) );
  INV_X1 U910 ( .A(n849), .ZN(n838) );
  NAND2_X1 U911 ( .A1(G95), .A2(n893), .ZN(n821) );
  NAND2_X1 U912 ( .A1(G107), .A2(n889), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n890), .A2(G119), .ZN(n822) );
  XOR2_X1 U915 ( .A(KEYINPUT94), .B(n822), .Z(n823) );
  NOR2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n894), .A2(G131), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n873) );
  NAND2_X1 U919 ( .A1(G1991), .A2(n873), .ZN(n835) );
  NAND2_X1 U920 ( .A1(G117), .A2(n889), .ZN(n828) );
  NAND2_X1 U921 ( .A1(G129), .A2(n890), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n893), .A2(G105), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT38), .B(n829), .Z(n830) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n894), .A2(G141), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n833), .A2(n832), .ZN(n874) );
  NAND2_X1 U928 ( .A1(G1996), .A2(n874), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT95), .B(n836), .Z(n999) );
  NAND2_X1 U931 ( .A1(n999), .A2(n852), .ZN(n837) );
  XOR2_X1 U932 ( .A(KEYINPUT96), .B(n837), .Z(n846) );
  NOR2_X1 U933 ( .A1(n838), .A2(n846), .ZN(n839) );
  AND2_X1 U934 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U935 ( .A1(n842), .A2(n841), .ZN(n855) );
  NAND2_X1 U936 ( .A1(n843), .A2(n902), .ZN(n1004) );
  NOR2_X1 U937 ( .A1(G1996), .A2(n874), .ZN(n995) );
  NOR2_X1 U938 ( .A1(G1991), .A2(n873), .ZN(n991) );
  NOR2_X1 U939 ( .A1(G1986), .A2(G290), .ZN(n844) );
  NOR2_X1 U940 ( .A1(n991), .A2(n844), .ZN(n845) );
  NOR2_X1 U941 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U942 ( .A1(n995), .A2(n847), .ZN(n848) );
  XNOR2_X1 U943 ( .A(n848), .B(KEYINPUT39), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n850), .A2(n849), .ZN(n851) );
  NAND2_X1 U945 ( .A1(n1004), .A2(n851), .ZN(n853) );
  NAND2_X1 U946 ( .A1(n853), .A2(n852), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U948 ( .A(KEYINPUT40), .B(n856), .ZN(G329) );
  NAND2_X1 U949 ( .A1(n857), .A2(G2106), .ZN(n858) );
  XNOR2_X1 U950 ( .A(n858), .B(KEYINPUT108), .ZN(G217) );
  NAND2_X1 U951 ( .A1(G15), .A2(G2), .ZN(n860) );
  INV_X1 U952 ( .A(G661), .ZN(n859) );
  NOR2_X1 U953 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U954 ( .A(n861), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U955 ( .A1(G3), .A2(G1), .ZN(n862) );
  NAND2_X1 U956 ( .A1(n863), .A2(n862), .ZN(G188) );
  XOR2_X1 U957 ( .A(G120), .B(KEYINPUT110), .Z(G236) );
  INV_X1 U959 ( .A(G108), .ZN(G238) );
  INV_X1 U960 ( .A(G96), .ZN(G221) );
  INV_X1 U961 ( .A(G57), .ZN(G237) );
  NOR2_X1 U962 ( .A1(n865), .A2(n864), .ZN(G325) );
  INV_X1 U963 ( .A(G325), .ZN(G261) );
  NAND2_X1 U964 ( .A1(G124), .A2(n890), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n889), .A2(G112), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G100), .A2(n893), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G136), .A2(n894), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n875) );
  XNOR2_X1 U973 ( .A(n992), .B(n875), .ZN(n886) );
  XOR2_X1 U974 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n884) );
  NAND2_X1 U975 ( .A1(G103), .A2(n893), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G139), .A2(n894), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G115), .A2(n889), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G127), .A2(n890), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n1006) );
  XNOR2_X1 U983 ( .A(n1006), .B(KEYINPUT115), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U985 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U986 ( .A(G160), .B(G162), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n904) );
  NAND2_X1 U988 ( .A1(G118), .A2(n889), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G130), .A2(n890), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U991 ( .A1(G106), .A2(n893), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G142), .A2(n894), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U994 ( .A(n897), .B(KEYINPUT45), .Z(n898) );
  NOR2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n900), .B(G164), .ZN(n901) );
  XOR2_X1 U997 ( .A(n902), .B(n901), .Z(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U999 ( .A1(G37), .A2(n905), .ZN(G395) );
  XOR2_X1 U1000 ( .A(n906), .B(n941), .Z(n908) );
  XNOR2_X1 U1001 ( .A(G286), .B(G171), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2474), .B(KEYINPUT112), .Z(n911) );
  XNOR2_X1 U1005 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1007 ( .A(n912), .B(KEYINPUT113), .Z(n914) );
  XNOR2_X1 U1008 ( .A(G1996), .B(G1991), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n922) );
  XOR2_X1 U1010 ( .A(G1976), .B(G1956), .Z(n916) );
  XNOR2_X1 U1011 ( .A(G1986), .B(G1971), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n920) );
  XOR2_X1 U1013 ( .A(KEYINPUT114), .B(G1981), .Z(n918) );
  XNOR2_X1 U1014 ( .A(G1961), .B(G1966), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n918), .B(n917), .ZN(n919) );
  XOR2_X1 U1016 ( .A(n920), .B(n919), .Z(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(G229) );
  XOR2_X1 U1018 ( .A(G2100), .B(G2096), .Z(n924) );
  XNOR2_X1 U1019 ( .A(KEYINPUT42), .B(G2678), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n924), .B(n923), .ZN(n928) );
  XOR2_X1 U1021 ( .A(KEYINPUT43), .B(G2072), .Z(n926) );
  XNOR2_X1 U1022 ( .A(G2067), .B(G2090), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n926), .B(n925), .ZN(n927) );
  XOR2_X1 U1024 ( .A(n928), .B(n927), .Z(n930) );
  XNOR2_X1 U1025 ( .A(G2078), .B(G2084), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n930), .B(n929), .ZN(G227) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(KEYINPUT116), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(G319), .A2(n932), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(G401), .A2(n933), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(G229), .A2(G227), .ZN(n934) );
  XOR2_X1 U1032 ( .A(KEYINPUT49), .B(n934), .Z(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(G225) );
  INV_X1 U1034 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1035 ( .A(KEYINPUT56), .B(G16), .ZN(n964) );
  XNOR2_X1 U1036 ( .A(G168), .B(G1966), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(n939), .B(KEYINPUT57), .ZN(n940) );
  XOR2_X1 U1039 ( .A(KEYINPUT121), .B(n940), .Z(n962) );
  XOR2_X1 U1040 ( .A(G1348), .B(n941), .Z(n942) );
  NOR2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G301), .B(G1961), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n944), .B(G1341), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n959) );
  INV_X1 U1046 ( .A(n949), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1048 ( .A(KEYINPUT122), .B(n952), .Z(n956) );
  XNOR2_X1 U1049 ( .A(G303), .B(G1971), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G299), .B(G1956), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1053 ( .A(KEYINPUT123), .B(n957), .Z(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(KEYINPUT124), .B(n960), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n1020) );
  XNOR2_X1 U1058 ( .A(KEYINPUT127), .B(G1966), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n965), .B(G21), .ZN(n978) );
  XOR2_X1 U1060 ( .A(G1956), .B(G20), .Z(n970) );
  XNOR2_X1 U1061 ( .A(G1341), .B(G19), .ZN(n967) );
  XNOR2_X1 U1062 ( .A(G1981), .B(G6), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(KEYINPUT126), .B(n968), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT59), .B(G1348), .Z(n971) );
  XNOR2_X1 U1067 ( .A(G4), .B(n971), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1069 ( .A(KEYINPUT60), .B(n974), .Z(n976) );
  XNOR2_X1 U1070 ( .A(G1961), .B(G5), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n985) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G22), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(G23), .B(G1976), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n982) );
  XOR2_X1 U1076 ( .A(G1986), .B(G24), .Z(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(KEYINPUT58), .B(n983), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(n986), .B(KEYINPUT61), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(G16), .B(KEYINPUT125), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(G11), .A2(n989), .ZN(n1018) );
  XOR2_X1 U1084 ( .A(G160), .B(G2084), .Z(n990) );
  NOR2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n998) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(n996), .B(KEYINPUT51), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n1002) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(KEYINPUT117), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1011) );
  XOR2_X1 U1095 ( .A(G2072), .B(n1006), .Z(n1008) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1009), .Z(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT52), .B(n1012), .ZN(n1014) );
  INV_X1 U1101 ( .A(KEYINPUT55), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(G29), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT118), .B(n1016), .Z(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1042) );
  XOR2_X1 U1107 ( .A(G2090), .B(G35), .Z(n1035) );
  XOR2_X1 U1108 ( .A(G1991), .B(G25), .Z(n1021) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(G28), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(G1996), .B(G32), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(n1022), .B(G27), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(n1025), .B(KEYINPUT119), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1031) );
  XNOR2_X1 U1115 ( .A(G2067), .B(G26), .ZN(n1029) );
  XNOR2_X1 U1116 ( .A(G2072), .B(G33), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(n1032), .B(KEYINPUT120), .ZN(n1033) );
  XNOR2_X1 U1120 ( .A(n1033), .B(KEYINPUT53), .ZN(n1034) );
  NAND2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(G34), .B(G2084), .ZN(n1036) );
  XNOR2_X1 U1123 ( .A(KEYINPUT54), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1125 ( .A(KEYINPUT55), .B(n1039), .Z(n1040) );
  NOR2_X1 U1126 ( .A1(G29), .A2(n1040), .ZN(n1041) );
  NOR2_X1 U1127 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XNOR2_X1 U1128 ( .A(n1043), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1129 ( .A(G311), .ZN(G150) );
endmodule

