

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U555 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X2 U556 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  INV_X1 U557 ( .A(KEYINPUT66), .ZN(n541) );
  NOR2_X1 U558 ( .A1(n636), .A2(n605), .ZN(n607) );
  INV_X1 U559 ( .A(KEYINPUT96), .ZN(n652) );
  BUF_X1 U560 ( .A(n734), .Z(n896) );
  NOR2_X2 U561 ( .A1(n547), .A2(n546), .ZN(G160) );
  AND2_X1 U562 ( .A1(n759), .A2(n1002), .ZN(n523) );
  NOR2_X1 U563 ( .A1(n536), .A2(n535), .ZN(G164) );
  XNOR2_X2 U564 ( .A(n529), .B(KEYINPUT65), .ZN(n734) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n524) );
  INV_X1 U566 ( .A(KEYINPUT26), .ZN(n606) );
  XNOR2_X1 U567 ( .A(n607), .B(n606), .ZN(n622) );
  INV_X1 U568 ( .A(KEYINPUT94), .ZN(n633) );
  INV_X1 U569 ( .A(KEYINPUT27), .ZN(n645) );
  XNOR2_X1 U570 ( .A(n646), .B(n645), .ZN(n649) );
  XNOR2_X1 U571 ( .A(n653), .B(n652), .ZN(n657) );
  NOR2_X1 U572 ( .A1(n673), .A2(n672), .ZN(n674) );
  BUF_X1 U573 ( .A(n636), .Z(n667) );
  NOR2_X1 U574 ( .A1(G164), .A2(G1384), .ZN(n746) );
  NAND2_X1 U575 ( .A1(n528), .A2(G2104), .ZN(n529) );
  INV_X1 U576 ( .A(KEYINPUT101), .ZN(n763) );
  NOR2_X2 U577 ( .A1(G2104), .A2(n525), .ZN(n900) );
  NOR2_X1 U578 ( .A1(G651), .A2(n588), .ZN(n807) );
  NAND2_X1 U579 ( .A1(n618), .A2(n617), .ZN(n996) );
  INV_X1 U580 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U581 ( .A1(G126), .A2(n900), .ZN(n527) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U583 ( .A1(G114), .A2(n901), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n527), .A2(n526), .ZN(n536) );
  INV_X1 U585 ( .A(G2105), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n734), .A2(G102), .ZN(n530) );
  XNOR2_X1 U587 ( .A(n530), .B(KEYINPUT86), .ZN(n533) );
  XOR2_X2 U588 ( .A(KEYINPUT17), .B(n531), .Z(n897) );
  NAND2_X1 U589 ( .A1(G138), .A2(n897), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U591 ( .A(KEYINPUT87), .B(n534), .Z(n535) );
  NAND2_X1 U592 ( .A1(n734), .A2(G101), .ZN(n537) );
  XNOR2_X1 U593 ( .A(n537), .B(KEYINPUT23), .ZN(n538) );
  INV_X1 U594 ( .A(n538), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n900), .A2(G125), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(n541), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n897), .A2(G137), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U600 ( .A1(G113), .A2(n901), .ZN(n545) );
  XNOR2_X1 U601 ( .A(KEYINPUT67), .B(n545), .ZN(n546) );
  XNOR2_X1 U602 ( .A(KEYINPUT68), .B(n524), .ZN(n588) );
  NAND2_X1 U603 ( .A1(G53), .A2(n807), .ZN(n550) );
  INV_X1 U604 ( .A(G651), .ZN(n551) );
  NOR2_X1 U605 ( .A1(G543), .A2(n551), .ZN(n548) );
  XOR2_X1 U606 ( .A(KEYINPUT1), .B(n548), .Z(n808) );
  NAND2_X1 U607 ( .A1(G65), .A2(n808), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n555) );
  NOR2_X1 U609 ( .A1(G543), .A2(G651), .ZN(n811) );
  NAND2_X1 U610 ( .A1(G91), .A2(n811), .ZN(n553) );
  NOR2_X2 U611 ( .A1(n551), .A2(n588), .ZN(n812) );
  NAND2_X1 U612 ( .A1(G78), .A2(n812), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n999) );
  INV_X1 U615 ( .A(n999), .ZN(G299) );
  NAND2_X1 U616 ( .A1(G52), .A2(n807), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G64), .A2(n808), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G90), .A2(n811), .ZN(n559) );
  NAND2_X1 U620 ( .A1(G77), .A2(n812), .ZN(n558) );
  NAND2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U623 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U624 ( .A1(n811), .A2(G89), .ZN(n563) );
  XNOR2_X1 U625 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G76), .A2(n812), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U628 ( .A(n566), .B(KEYINPUT5), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G51), .A2(n807), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G63), .A2(n808), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U632 ( .A(KEYINPUT6), .B(n569), .Z(n570) );
  NAND2_X1 U633 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n572), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U635 ( .A(G168), .B(KEYINPUT8), .Z(n573) );
  XNOR2_X1 U636 ( .A(KEYINPUT76), .B(n573), .ZN(G286) );
  NAND2_X1 U637 ( .A1(G88), .A2(n811), .ZN(n575) );
  NAND2_X1 U638 ( .A1(G75), .A2(n812), .ZN(n574) );
  NAND2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n808), .A2(G62), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G50), .A2(n807), .ZN(n576) );
  XOR2_X1 U642 ( .A(KEYINPUT81), .B(n576), .Z(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(G166) );
  INV_X1 U645 ( .A(G166), .ZN(G303) );
  NAND2_X1 U646 ( .A1(G86), .A2(n811), .ZN(n582) );
  NAND2_X1 U647 ( .A1(G61), .A2(n808), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n812), .A2(G73), .ZN(n583) );
  XOR2_X1 U650 ( .A(KEYINPUT2), .B(n583), .Z(n584) );
  NOR2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n807), .A2(G48), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U654 ( .A1(G74), .A2(G651), .ZN(n593) );
  NAND2_X1 U655 ( .A1(G49), .A2(n807), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G87), .A2(n588), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U658 ( .A1(n808), .A2(n591), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n594), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U661 ( .A1(G60), .A2(n808), .ZN(n601) );
  NAND2_X1 U662 ( .A1(G47), .A2(n807), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G85), .A2(n811), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U665 ( .A1(G72), .A2(n812), .ZN(n597) );
  XNOR2_X1 U666 ( .A(KEYINPUT69), .B(n597), .ZN(n598) );
  NOR2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U669 ( .A(n602), .B(KEYINPUT70), .ZN(G290) );
  INV_X1 U670 ( .A(KEYINPUT64), .ZN(n624) );
  NAND2_X1 U671 ( .A1(G160), .A2(G40), .ZN(n747) );
  INV_X1 U672 ( .A(KEYINPUT90), .ZN(n603) );
  XNOR2_X1 U673 ( .A(n747), .B(n603), .ZN(n604) );
  NAND2_X2 U674 ( .A1(n604), .A2(n746), .ZN(n636) );
  INV_X1 U675 ( .A(G1996), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n636), .A2(G1341), .ZN(n620) );
  NAND2_X1 U677 ( .A1(G68), .A2(n812), .ZN(n611) );
  NAND2_X1 U678 ( .A1(G81), .A2(n811), .ZN(n608) );
  XNOR2_X1 U679 ( .A(n608), .B(KEYINPUT72), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n609), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n613) );
  XNOR2_X1 U682 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n612) );
  XNOR2_X1 U683 ( .A(n613), .B(n612), .ZN(n616) );
  NAND2_X1 U684 ( .A1(n808), .A2(G56), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT14), .B(n614), .Z(n615) );
  NOR2_X1 U686 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U687 ( .A1(n807), .A2(G43), .ZN(n617) );
  INV_X1 U688 ( .A(n996), .ZN(n619) );
  AND2_X1 U689 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U690 ( .A(n624), .B(n623), .ZN(n641) );
  NAND2_X1 U691 ( .A1(n807), .A2(G54), .ZN(n631) );
  NAND2_X1 U692 ( .A1(G79), .A2(n812), .ZN(n626) );
  NAND2_X1 U693 ( .A1(G66), .A2(n808), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U695 ( .A1(n811), .A2(G92), .ZN(n627) );
  XOR2_X1 U696 ( .A(KEYINPUT74), .B(n627), .Z(n628) );
  NOR2_X1 U697 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U699 ( .A(KEYINPUT15), .B(n632), .ZN(n991) );
  INV_X1 U700 ( .A(n991), .ZN(n642) );
  NOR2_X1 U701 ( .A1(n641), .A2(n642), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(n633), .ZN(n640) );
  INV_X1 U703 ( .A(n636), .ZN(n659) );
  XOR2_X2 U704 ( .A(KEYINPUT93), .B(n659), .Z(n661) );
  NAND2_X1 U705 ( .A1(n661), .A2(G2067), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT95), .B(n635), .Z(n638) );
  NAND2_X1 U707 ( .A1(G1348), .A2(n667), .ZN(n637) );
  NAND2_X1 U708 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U710 ( .A1(n641), .A2(n642), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n651) );
  NAND2_X1 U712 ( .A1(n661), .A2(G2072), .ZN(n646) );
  INV_X1 U713 ( .A(n661), .ZN(n647) );
  NAND2_X1 U714 ( .A1(G1956), .A2(n647), .ZN(n648) );
  NAND2_X1 U715 ( .A1(n649), .A2(n648), .ZN(n654) );
  OR2_X1 U716 ( .A1(G299), .A2(n654), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U718 ( .A1(G299), .A2(n654), .ZN(n655) );
  XOR2_X1 U719 ( .A(KEYINPUT28), .B(n655), .Z(n656) );
  NOR2_X1 U720 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U721 ( .A(n658), .B(KEYINPUT29), .ZN(n665) );
  NOR2_X1 U722 ( .A1(n659), .A2(G1961), .ZN(n660) );
  XOR2_X1 U723 ( .A(KEYINPUT92), .B(n660), .Z(n663) );
  XNOR2_X1 U724 ( .A(G2078), .B(KEYINPUT25), .ZN(n968) );
  NAND2_X1 U725 ( .A1(n661), .A2(n968), .ZN(n662) );
  NAND2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U727 ( .A1(G171), .A2(n666), .ZN(n664) );
  NAND2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n676) );
  NOR2_X1 U729 ( .A1(G171), .A2(n666), .ZN(n673) );
  NAND2_X1 U730 ( .A1(G8), .A2(n667), .ZN(n668) );
  XNOR2_X2 U731 ( .A(KEYINPUT91), .B(n668), .ZN(n714) );
  INV_X1 U732 ( .A(n714), .ZN(n705) );
  NOR2_X2 U733 ( .A1(G1966), .A2(n705), .ZN(n689) );
  NOR2_X1 U734 ( .A1(G2084), .A2(n667), .ZN(n687) );
  NOR2_X1 U735 ( .A1(n689), .A2(n687), .ZN(n669) );
  NAND2_X1 U736 ( .A1(G8), .A2(n669), .ZN(n670) );
  XNOR2_X1 U737 ( .A(KEYINPUT30), .B(n670), .ZN(n671) );
  NOR2_X1 U738 ( .A1(G168), .A2(n671), .ZN(n672) );
  XOR2_X1 U739 ( .A(KEYINPUT31), .B(n674), .Z(n675) );
  NAND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n688) );
  AND2_X1 U741 ( .A1(G286), .A2(G8), .ZN(n677) );
  NAND2_X1 U742 ( .A1(n688), .A2(n677), .ZN(n684) );
  INV_X1 U743 ( .A(G8), .ZN(n682) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n705), .ZN(n679) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n667), .ZN(n678) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U747 ( .A1(n680), .A2(G303), .ZN(n681) );
  OR2_X1 U748 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n686) );
  INV_X1 U750 ( .A(KEYINPUT32), .ZN(n685) );
  XNOR2_X1 U751 ( .A(n686), .B(n685), .ZN(n694) );
  NAND2_X1 U752 ( .A1(G8), .A2(n687), .ZN(n692) );
  XNOR2_X1 U753 ( .A(KEYINPUT97), .B(n688), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U756 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U757 ( .A(n695), .B(KEYINPUT98), .ZN(n709) );
  NOR2_X1 U758 ( .A1(G2090), .A2(G303), .ZN(n696) );
  NAND2_X1 U759 ( .A1(G8), .A2(n696), .ZN(n697) );
  NAND2_X1 U760 ( .A1(n709), .A2(n697), .ZN(n698) );
  NAND2_X1 U761 ( .A1(n698), .A2(n705), .ZN(n728) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n1006) );
  XOR2_X1 U763 ( .A(n1006), .B(KEYINPUT99), .Z(n699) );
  NOR2_X1 U764 ( .A1(KEYINPUT33), .A2(n699), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n714), .A2(KEYINPUT100), .ZN(n700) );
  XNOR2_X1 U766 ( .A(G1981), .B(G305), .ZN(n989) );
  NOR2_X1 U767 ( .A1(n700), .A2(n989), .ZN(n711) );
  INV_X1 U768 ( .A(n711), .ZN(n701) );
  OR2_X1 U769 ( .A1(G1976), .A2(G288), .ZN(n1003) );
  OR2_X1 U770 ( .A1(n701), .A2(n1003), .ZN(n710) );
  AND2_X1 U771 ( .A1(n702), .A2(n710), .ZN(n707) );
  NOR2_X1 U772 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U773 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  NOR2_X1 U774 ( .A1(n705), .A2(n704), .ZN(n724) );
  INV_X1 U775 ( .A(n724), .ZN(n706) );
  AND2_X1 U776 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n726) );
  INV_X1 U778 ( .A(n710), .ZN(n713) );
  AND2_X1 U779 ( .A1(KEYINPUT100), .A2(n711), .ZN(n712) );
  NOR2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n722) );
  NAND2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n995) );
  AND2_X1 U782 ( .A1(n714), .A2(KEYINPUT100), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n995), .A2(n717), .ZN(n715) );
  INV_X1 U784 ( .A(KEYINPUT33), .ZN(n716) );
  NAND2_X1 U785 ( .A1(n715), .A2(n716), .ZN(n720) );
  NOR2_X1 U786 ( .A1(n716), .A2(n1003), .ZN(n718) );
  NAND2_X1 U787 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n723) );
  OR2_X1 U790 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U792 ( .A1(n728), .A2(n727), .ZN(n762) );
  NAND2_X1 U793 ( .A1(G131), .A2(n897), .ZN(n730) );
  NAND2_X1 U794 ( .A1(G119), .A2(n900), .ZN(n729) );
  NAND2_X1 U795 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U796 ( .A1(G107), .A2(n901), .ZN(n731) );
  XNOR2_X1 U797 ( .A(KEYINPUT89), .B(n731), .ZN(n732) );
  NOR2_X1 U798 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U799 ( .A1(n896), .A2(G95), .ZN(n735) );
  NAND2_X1 U800 ( .A1(n736), .A2(n735), .ZN(n891) );
  AND2_X1 U801 ( .A1(n891), .A2(G1991), .ZN(n745) );
  NAND2_X1 U802 ( .A1(G129), .A2(n900), .ZN(n738) );
  NAND2_X1 U803 ( .A1(G117), .A2(n901), .ZN(n737) );
  NAND2_X1 U804 ( .A1(n738), .A2(n737), .ZN(n741) );
  NAND2_X1 U805 ( .A1(n896), .A2(G105), .ZN(n739) );
  XOR2_X1 U806 ( .A(KEYINPUT38), .B(n739), .Z(n740) );
  NOR2_X1 U807 ( .A1(n741), .A2(n740), .ZN(n743) );
  NAND2_X1 U808 ( .A1(n897), .A2(G141), .ZN(n742) );
  NAND2_X1 U809 ( .A1(n743), .A2(n742), .ZN(n907) );
  AND2_X1 U810 ( .A1(n907), .A2(G1996), .ZN(n744) );
  NOR2_X1 U811 ( .A1(n745), .A2(n744), .ZN(n1027) );
  NOR2_X1 U812 ( .A1(n747), .A2(n746), .ZN(n759) );
  INV_X1 U813 ( .A(n759), .ZN(n777) );
  NOR2_X1 U814 ( .A1(n1027), .A2(n777), .ZN(n767) );
  INV_X1 U815 ( .A(n767), .ZN(n758) );
  NAND2_X1 U816 ( .A1(n897), .A2(G140), .ZN(n748) );
  XNOR2_X1 U817 ( .A(n748), .B(KEYINPUT88), .ZN(n750) );
  NAND2_X1 U818 ( .A1(G104), .A2(n896), .ZN(n749) );
  NAND2_X1 U819 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U820 ( .A(KEYINPUT34), .B(n751), .ZN(n756) );
  NAND2_X1 U821 ( .A1(G128), .A2(n900), .ZN(n753) );
  NAND2_X1 U822 ( .A1(G116), .A2(n901), .ZN(n752) );
  NAND2_X1 U823 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U824 ( .A(KEYINPUT35), .B(n754), .Z(n755) );
  NOR2_X1 U825 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U826 ( .A(KEYINPUT36), .B(n757), .Z(n912) );
  XOR2_X1 U827 ( .A(G2067), .B(KEYINPUT37), .Z(n774) );
  AND2_X1 U828 ( .A1(n912), .A2(n774), .ZN(n1041) );
  NAND2_X1 U829 ( .A1(n759), .A2(n1041), .ZN(n771) );
  NAND2_X1 U830 ( .A1(n758), .A2(n771), .ZN(n760) );
  XNOR2_X1 U831 ( .A(G1986), .B(G290), .ZN(n1002) );
  NOR2_X1 U832 ( .A1(n760), .A2(n523), .ZN(n761) );
  NAND2_X1 U833 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U834 ( .A(n764), .B(n763), .ZN(n780) );
  NOR2_X1 U835 ( .A1(G1996), .A2(n907), .ZN(n1024) );
  NOR2_X1 U836 ( .A1(G1986), .A2(G290), .ZN(n765) );
  NOR2_X1 U837 ( .A1(G1991), .A2(n891), .ZN(n1020) );
  NOR2_X1 U838 ( .A1(n765), .A2(n1020), .ZN(n766) );
  NOR2_X1 U839 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U840 ( .A1(n1024), .A2(n768), .ZN(n769) );
  XNOR2_X1 U841 ( .A(KEYINPUT39), .B(n769), .ZN(n770) );
  XNOR2_X1 U842 ( .A(n770), .B(KEYINPUT102), .ZN(n772) );
  NAND2_X1 U843 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U844 ( .A(KEYINPUT103), .B(n773), .ZN(n775) );
  NOR2_X1 U845 ( .A1(n912), .A2(n774), .ZN(n1037) );
  NOR2_X1 U846 ( .A1(n775), .A2(n1037), .ZN(n776) );
  NOR2_X1 U847 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U848 ( .A(KEYINPUT104), .B(n778), .Z(n779) );
  NAND2_X1 U849 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U850 ( .A(n781), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U851 ( .A(G171), .ZN(G301) );
  AND2_X1 U852 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U853 ( .A(G132), .ZN(G219) );
  INV_X1 U854 ( .A(G82), .ZN(G220) );
  INV_X1 U855 ( .A(G57), .ZN(G237) );
  INV_X1 U856 ( .A(G69), .ZN(G235) );
  INV_X1 U857 ( .A(G108), .ZN(G238) );
  INV_X1 U858 ( .A(G120), .ZN(G236) );
  XOR2_X1 U859 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n783) );
  NAND2_X1 U860 ( .A1(G7), .A2(G661), .ZN(n782) );
  XOR2_X1 U861 ( .A(n783), .B(n782), .Z(n847) );
  NAND2_X1 U862 ( .A1(n847), .A2(G567), .ZN(n784) );
  XOR2_X1 U863 ( .A(KEYINPUT11), .B(n784), .Z(G234) );
  INV_X1 U864 ( .A(G860), .ZN(n791) );
  OR2_X1 U865 ( .A1(n996), .A2(n791), .ZN(G153) );
  NOR2_X1 U866 ( .A1(n991), .A2(G868), .ZN(n785) );
  XNOR2_X1 U867 ( .A(n785), .B(KEYINPUT75), .ZN(n787) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n787), .A2(n786), .ZN(G284) );
  INV_X1 U870 ( .A(G868), .ZN(n829) );
  NAND2_X1 U871 ( .A1(n999), .A2(n829), .ZN(n788) );
  XNOR2_X1 U872 ( .A(n788), .B(KEYINPUT77), .ZN(n790) );
  NOR2_X1 U873 ( .A1(G286), .A2(n829), .ZN(n789) );
  NOR2_X1 U874 ( .A1(n790), .A2(n789), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n791), .A2(G559), .ZN(n792) );
  NAND2_X1 U876 ( .A1(n792), .A2(n991), .ZN(n793) );
  XNOR2_X1 U877 ( .A(n793), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U878 ( .A1(n991), .A2(G868), .ZN(n794) );
  NOR2_X1 U879 ( .A1(G559), .A2(n794), .ZN(n795) );
  XNOR2_X1 U880 ( .A(n795), .B(KEYINPUT78), .ZN(n797) );
  NOR2_X1 U881 ( .A1(n996), .A2(G868), .ZN(n796) );
  NOR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(G282) );
  NAND2_X1 U883 ( .A1(G123), .A2(n900), .ZN(n798) );
  XNOR2_X1 U884 ( .A(n798), .B(KEYINPUT18), .ZN(n800) );
  NAND2_X1 U885 ( .A1(n896), .A2(G99), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G135), .A2(n897), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G111), .A2(n901), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n1019) );
  XNOR2_X1 U891 ( .A(G2096), .B(n1019), .ZN(n805) );
  INV_X1 U892 ( .A(G2100), .ZN(n870) );
  NAND2_X1 U893 ( .A1(n805), .A2(n870), .ZN(G156) );
  NAND2_X1 U894 ( .A1(n991), .A2(G559), .ZN(n826) );
  XNOR2_X1 U895 ( .A(n996), .B(n826), .ZN(n806) );
  NOR2_X1 U896 ( .A1(n806), .A2(G860), .ZN(n818) );
  NAND2_X1 U897 ( .A1(G55), .A2(n807), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G67), .A2(n808), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n817) );
  NAND2_X1 U900 ( .A1(G93), .A2(n811), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G80), .A2(n812), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U903 ( .A(KEYINPUT79), .B(n815), .Z(n816) );
  OR2_X1 U904 ( .A1(n817), .A2(n816), .ZN(n828) );
  XOR2_X1 U905 ( .A(n818), .B(n828), .Z(G145) );
  XNOR2_X1 U906 ( .A(n828), .B(KEYINPUT82), .ZN(n820) );
  XOR2_X1 U907 ( .A(G299), .B(KEYINPUT19), .Z(n819) );
  XNOR2_X1 U908 ( .A(n820), .B(n819), .ZN(n823) );
  XOR2_X1 U909 ( .A(G290), .B(G166), .Z(n821) );
  XNOR2_X1 U910 ( .A(n821), .B(G305), .ZN(n822) );
  XNOR2_X1 U911 ( .A(n823), .B(n822), .ZN(n825) );
  XNOR2_X1 U912 ( .A(n996), .B(G288), .ZN(n824) );
  XNOR2_X1 U913 ( .A(n825), .B(n824), .ZN(n917) );
  XNOR2_X1 U914 ( .A(n826), .B(n917), .ZN(n827) );
  NAND2_X1 U915 ( .A1(n827), .A2(G868), .ZN(n831) );
  NAND2_X1 U916 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U917 ( .A1(n831), .A2(n830), .ZN(G295) );
  NAND2_X1 U918 ( .A1(G2084), .A2(G2078), .ZN(n832) );
  XOR2_X1 U919 ( .A(KEYINPUT20), .B(n832), .Z(n833) );
  NAND2_X1 U920 ( .A1(G2090), .A2(n833), .ZN(n834) );
  XNOR2_X1 U921 ( .A(KEYINPUT21), .B(n834), .ZN(n835) );
  NAND2_X1 U922 ( .A1(n835), .A2(G2072), .ZN(n836) );
  XOR2_X1 U923 ( .A(KEYINPUT83), .B(n836), .Z(G158) );
  XNOR2_X1 U924 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U925 ( .A1(G236), .A2(G238), .ZN(n838) );
  NOR2_X1 U926 ( .A1(G235), .A2(G237), .ZN(n837) );
  NAND2_X1 U927 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U928 ( .A(KEYINPUT84), .B(n839), .ZN(n853) );
  NAND2_X1 U929 ( .A1(G567), .A2(n853), .ZN(n844) );
  NOR2_X1 U930 ( .A1(G220), .A2(G219), .ZN(n840) );
  XOR2_X1 U931 ( .A(KEYINPUT22), .B(n840), .Z(n841) );
  NOR2_X1 U932 ( .A1(G218), .A2(n841), .ZN(n842) );
  NAND2_X1 U933 ( .A1(G96), .A2(n842), .ZN(n852) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n852), .ZN(n843) );
  NAND2_X1 U935 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U936 ( .A(KEYINPUT85), .B(n845), .Z(n851) );
  NAND2_X1 U937 ( .A1(G661), .A2(G483), .ZN(n846) );
  NOR2_X1 U938 ( .A1(n851), .A2(n846), .ZN(n850) );
  NAND2_X1 U939 ( .A1(n850), .A2(G36), .ZN(G176) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n847), .ZN(G217) );
  INV_X1 U941 ( .A(n847), .ZN(G223) );
  AND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n848) );
  NAND2_X1 U943 ( .A1(G661), .A2(n848), .ZN(G259) );
  NAND2_X1 U944 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(G188) );
  INV_X1 U946 ( .A(n851), .ZN(G319) );
  INV_X1 U948 ( .A(G96), .ZN(G221) );
  NOR2_X1 U949 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U950 ( .A(G325), .ZN(G261) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1986), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1971), .B(G1976), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U954 ( .A(n856), .B(KEYINPUT109), .Z(n858) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U957 ( .A(G1981), .B(G1956), .Z(n860) );
  XNOR2_X1 U958 ( .A(G1966), .B(G1961), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U960 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U961 ( .A(KEYINPUT110), .B(G2474), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(G229) );
  XOR2_X1 U963 ( .A(G2096), .B(G2678), .Z(n866) );
  XNOR2_X1 U964 ( .A(G2072), .B(KEYINPUT43), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U966 ( .A(n867), .B(KEYINPUT42), .Z(n869) );
  XNOR2_X1 U967 ( .A(G2090), .B(G2067), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n874) );
  XNOR2_X1 U969 ( .A(KEYINPUT108), .B(n870), .ZN(n872) );
  XNOR2_X1 U970 ( .A(G2084), .B(G2078), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(G227) );
  NAND2_X1 U973 ( .A1(G124), .A2(n900), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U975 ( .A1(n896), .A2(G100), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G136), .A2(n897), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G112), .A2(n901), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U980 ( .A1(n881), .A2(n880), .ZN(G162) );
  NAND2_X1 U981 ( .A1(G118), .A2(n901), .ZN(n890) );
  NAND2_X1 U982 ( .A1(n900), .A2(G130), .ZN(n882) );
  XNOR2_X1 U983 ( .A(KEYINPUT111), .B(n882), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G106), .A2(n896), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G142), .A2(n897), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U987 ( .A(KEYINPUT112), .B(n885), .Z(n886) );
  XNOR2_X1 U988 ( .A(KEYINPUT45), .B(n886), .ZN(n887) );
  NOR2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n895) );
  XOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n893) );
  XOR2_X1 U992 ( .A(n891), .B(KEYINPUT113), .Z(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n911) );
  XOR2_X1 U995 ( .A(n1019), .B(G162), .Z(n909) );
  NAND2_X1 U996 ( .A1(G103), .A2(n896), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G139), .A2(n897), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n906) );
  NAND2_X1 U999 ( .A1(G127), .A2(n900), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n901), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n1030) );
  XOR2_X1 U1004 ( .A(n907), .B(n1030), .Z(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n911), .B(n910), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G164), .B(n912), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(G160), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n916), .ZN(G395) );
  XOR2_X1 U1011 ( .A(n917), .B(n991), .Z(n918) );
  XNOR2_X1 U1012 ( .A(n918), .B(G286), .ZN(n919) );
  XOR2_X1 U1013 ( .A(n919), .B(G301), .Z(n920) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n920), .ZN(G397) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n922) );
  XNOR2_X1 U1016 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n936) );
  XOR2_X1 U1018 ( .A(KEYINPUT106), .B(G2443), .Z(n924) );
  XNOR2_X1 U1019 ( .A(G2451), .B(G2427), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1021 ( .A(n925), .B(G2430), .Z(n927) );
  XNOR2_X1 U1022 ( .A(G1348), .B(G1341), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n931) );
  XOR2_X1 U1024 ( .A(KEYINPUT107), .B(G2435), .Z(n929) );
  XNOR2_X1 U1025 ( .A(G2438), .B(G2454), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(n929), .B(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(n931), .B(n930), .Z(n933) );
  XNOR2_X1 U1028 ( .A(G2446), .B(KEYINPUT105), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n933), .B(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(G14), .ZN(n939) );
  NAND2_X1 U1031 ( .A1(G319), .A2(n939), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(G395), .A2(G397), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(G225) );
  INV_X1 U1035 ( .A(G225), .ZN(G308) );
  INV_X1 U1036 ( .A(n939), .ZN(G401) );
  XNOR2_X1 U1037 ( .A(G1986), .B(G24), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G1971), .B(G22), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G23), .B(G1976), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(KEYINPUT125), .B(n942), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(KEYINPUT58), .B(n945), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(n946), .B(KEYINPUT126), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G21), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G5), .B(G1961), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n961) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(G6), .B(G1981), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n958) );
  XOR2_X1 U1052 ( .A(KEYINPUT124), .B(G4), .Z(n954) );
  XNOR2_X1 U1053 ( .A(G1348), .B(KEYINPUT59), .ZN(n953) );
  XNOR2_X1 U1054 ( .A(n954), .B(n953), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(G1956), .B(G20), .ZN(n955) );
  NOR2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(KEYINPUT60), .B(n959), .ZN(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(n962), .B(KEYINPUT127), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(KEYINPUT61), .B(n963), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(G16), .A2(n964), .ZN(n1049) );
  XNOR2_X1 U1063 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n1043) );
  XNOR2_X1 U1064 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1065 ( .A(G1991), .B(G25), .ZN(n965) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n975) );
  XOR2_X1 U1067 ( .A(G2072), .B(G33), .Z(n967) );
  NAND2_X1 U1068 ( .A1(n967), .A2(G28), .ZN(n973) );
  XOR2_X1 U1069 ( .A(n968), .B(G27), .Z(n970) );
  XNOR2_X1 U1070 ( .A(G32), .B(G1996), .ZN(n969) );
  NOR2_X1 U1071 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1072 ( .A(n971), .B(KEYINPUT119), .ZN(n972) );
  NOR2_X1 U1073 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1074 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1075 ( .A(n976), .B(KEYINPUT53), .ZN(n979) );
  XOR2_X1 U1076 ( .A(G2084), .B(G34), .Z(n977) );
  XNOR2_X1 U1077 ( .A(KEYINPUT54), .B(n977), .ZN(n978) );
  NAND2_X1 U1078 ( .A1(n979), .A2(n978), .ZN(n982) );
  XNOR2_X1 U1079 ( .A(KEYINPUT118), .B(G2090), .ZN(n980) );
  XNOR2_X1 U1080 ( .A(G35), .B(n980), .ZN(n981) );
  NOR2_X1 U1081 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1082 ( .A(n1043), .B(n983), .Z(n985) );
  INV_X1 U1083 ( .A(G29), .ZN(n984) );
  NAND2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1085 ( .A1(n986), .A2(G11), .ZN(n987) );
  XNOR2_X1 U1086 ( .A(n987), .B(KEYINPUT120), .ZN(n1018) );
  XOR2_X1 U1087 ( .A(G168), .B(G1966), .Z(n988) );
  NOR2_X1 U1088 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1089 ( .A(KEYINPUT57), .B(n990), .Z(n1012) );
  XOR2_X1 U1090 ( .A(G301), .B(G1961), .Z(n993) );
  XNOR2_X1 U1091 ( .A(G1348), .B(n991), .ZN(n992) );
  NAND2_X1 U1092 ( .A1(n993), .A2(n992), .ZN(n1010) );
  NAND2_X1 U1093 ( .A1(G1971), .A2(G303), .ZN(n994) );
  NAND2_X1 U1094 ( .A1(n995), .A2(n994), .ZN(n998) );
  XNOR2_X1 U1095 ( .A(G1341), .B(n996), .ZN(n997) );
  NOR2_X1 U1096 ( .A1(n998), .A2(n997), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G1956), .B(KEYINPUT122), .ZN(n1000) );
  XOR2_X1 U1098 ( .A(n1000), .B(n999), .Z(n1001) );
  NOR2_X1 U1099 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1100 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1101 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1102 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(KEYINPUT123), .B(n1013), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(G16), .B(KEYINPUT121), .ZN(n1014) );
  XNOR2_X1 U1107 ( .A(n1014), .B(KEYINPUT56), .ZN(n1015) );
  NOR2_X1 U1108 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1047) );
  XNOR2_X1 U1110 ( .A(G160), .B(G2084), .ZN(n1022) );
  NOR2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(G2090), .B(G162), .Z(n1023) );
  NOR2_X1 U1114 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1115 ( .A(KEYINPUT51), .B(n1025), .Z(n1026) );
  NAND2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1039) );
  XNOR2_X1 U1118 ( .A(G2072), .B(n1030), .ZN(n1033) );
  XOR2_X1 U1119 ( .A(G164), .B(G2078), .Z(n1031) );
  XNOR2_X1 U1120 ( .A(KEYINPUT115), .B(n1031), .ZN(n1032) );
  NAND2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1122 ( .A(n1034), .B(KEYINPUT116), .ZN(n1035) );
  XNOR2_X1 U1123 ( .A(n1035), .B(KEYINPUT50), .ZN(n1036) );
  NOR2_X1 U1124 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1125 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NOR2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1127 ( .A(KEYINPUT52), .B(n1042), .ZN(n1044) );
  NAND2_X1 U1128 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NAND2_X1 U1129 ( .A1(n1045), .A2(G29), .ZN(n1046) );
  NAND2_X1 U1130 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NOR2_X1 U1131 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  XOR2_X1 U1132 ( .A(KEYINPUT62), .B(n1050), .Z(G150) );
  INV_X1 U1133 ( .A(G150), .ZN(G311) );
endmodule

