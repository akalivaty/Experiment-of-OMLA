//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT5), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT81), .B(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n219), .B2(KEYINPUT2), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G141gat), .B(G148gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n216), .B(new_n219), .C1(new_n222), .C2(KEYINPUT2), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n211), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n221), .A2(KEYINPUT83), .A3(new_n226), .A4(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n221), .A2(KEYINPUT82), .A3(new_n223), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(KEYINPUT3), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT85), .ZN(new_n238));
  INV_X1    g037(.A(new_n235), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n234), .B(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n221), .A3(new_n223), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n238), .B1(new_n241), .B2(KEYINPUT4), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n236), .A2(new_n224), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(KEYINPUT85), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(new_n243), .B2(new_n244), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(new_n248), .A3(new_n245), .ZN(new_n251));
  AOI221_X4 g050(.A(new_n210), .B1(new_n228), .B2(new_n237), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n228), .A2(new_n236), .A3(new_n232), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n243), .A2(new_n244), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n253), .B(new_n207), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT5), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n230), .A2(new_n236), .A3(new_n231), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n241), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n257), .B1(new_n259), .B2(new_n208), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n206), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n250), .A2(new_n251), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n253), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n205), .B(new_n261), .C1(new_n265), .C2(new_n210), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(KEYINPUT6), .B(new_n206), .C1(new_n252), .C2(new_n262), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT69), .B1(new_n273), .B2(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT27), .B(G183gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n272), .B(new_n274), .C1(new_n275), .C2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(KEYINPUT28), .A3(new_n272), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(KEYINPUT70), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n282), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n293), .A2(KEYINPUT71), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT71), .B1(new_n293), .B2(new_n294), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n280), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n290), .B1(KEYINPUT23), .B2(new_n281), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT23), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT25), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT67), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n273), .A2(new_n272), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n301), .B(new_n302), .C1(new_n309), .C2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n310), .B(new_n311), .C1(new_n306), .C2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n304), .A2(KEYINPUT65), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT66), .B(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n321));
  OAI22_X1  g120(.A1(new_n319), .A2(new_n320), .B1(new_n321), .B2(new_n290), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n314), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n312), .B1(new_n305), .B2(new_n308), .ZN(new_n324));
  OAI211_X1 g123(.A(KEYINPUT25), .B(new_n299), .C1(new_n321), .C2(new_n290), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT68), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n313), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n271), .B1(new_n297), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n297), .A2(new_n327), .ZN(new_n329));
  XOR2_X1   g128(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n331), .B2(new_n271), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  AND2_X1   g133(.A1(G211gat), .A2(G218gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n334), .B1(KEYINPUT22), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT76), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n328), .ZN(new_n341));
  INV_X1    g140(.A(new_n338), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT29), .B1(new_n297), .B2(new_n327), .ZN(new_n343));
  INV_X1    g142(.A(new_n271), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT78), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n340), .A2(new_n352), .A3(new_n345), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n347), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n340), .A2(KEYINPUT30), .A3(new_n345), .A4(new_n350), .ZN(new_n355));
  INV_X1    g154(.A(new_n339), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n345), .B(new_n350), .C1(new_n332), .C2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n354), .B(new_n355), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n270), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT89), .ZN(new_n364));
  INV_X1    g163(.A(G22gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n230), .A2(new_n231), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n226), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n330), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n370), .B1(new_n225), .B2(new_n227), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT87), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n339), .B1(new_n371), .B2(KEYINPUT87), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n226), .B1(new_n338), .B2(new_n370), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n224), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n371), .B2(new_n342), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n366), .B(KEYINPUT86), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n365), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n375), .A2(new_n365), .A3(new_n380), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n364), .B1(new_n384), .B2(KEYINPUT88), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387));
  AOI211_X1 g186(.A(new_n387), .B(KEYINPUT89), .C1(new_n382), .C2(new_n383), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G78gat), .B(G106gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT31), .ZN(new_n391));
  INV_X1    g190(.A(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n382), .A2(new_n383), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n387), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n386), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n393), .B1(new_n384), .B2(KEYINPUT88), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n398), .B1(new_n385), .B2(new_n388), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n363), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT39), .B1(new_n259), .B2(new_n208), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT90), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n250), .A2(new_n251), .B1(new_n228), .B2(new_n237), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n402), .B1(new_n403), .B2(new_n207), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT39), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n265), .A2(new_n405), .A3(new_n208), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n406), .A3(new_n205), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT40), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT40), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n408), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n410), .A2(new_n362), .A3(new_n263), .A4(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n413), .A2(new_n397), .A3(new_n399), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n347), .A2(KEYINPUT37), .A3(new_n353), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n340), .A2(new_n416), .A3(new_n345), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n351), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT38), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n343), .A2(new_n344), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n338), .B1(new_n420), .B2(new_n328), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n333), .B2(new_n339), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT38), .B1(new_n422), .B2(KEYINPUT37), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n423), .A2(new_n351), .A3(new_n417), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n268), .A2(new_n424), .A3(new_n269), .A4(new_n357), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT92), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n425), .A2(new_n426), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n419), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n400), .B1(new_n414), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n297), .A2(new_n240), .A3(new_n327), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT72), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n297), .A2(new_n327), .A3(new_n434), .A4(new_n240), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n329), .A2(new_n236), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT34), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n437), .A2(KEYINPUT73), .A3(new_n438), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT73), .B1(new_n437), .B2(new_n438), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT32), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n443), .B2(new_n444), .ZN(new_n447));
  XOR2_X1   g246(.A(G15gat), .B(G43gat), .Z(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT74), .ZN(new_n452));
  INV_X1    g251(.A(new_n450), .ZN(new_n453));
  OAI221_X1 g252(.A(KEYINPUT32), .B1(new_n446), .B2(new_n453), .C1(new_n443), .C2(new_n444), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n451), .B2(new_n454), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n442), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n451), .A2(new_n441), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT36), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n431), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n431), .A3(new_n460), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  INV_X1    g262(.A(new_n458), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n441), .B1(new_n451), .B2(new_n454), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n430), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n397), .A2(new_n399), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(new_n457), .A3(new_n363), .A4(new_n458), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT35), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n397), .A2(new_n399), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n464), .A2(new_n465), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n475), .A3(new_n363), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT15), .ZN(new_n479));
  OR2_X1    g278(.A1(G43gat), .A2(G50gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(G43gat), .A2(G50gat), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(KEYINPUT93), .B(G43gat), .Z(new_n483));
  OAI211_X1 g282(.A(new_n479), .B(new_n481), .C1(new_n483), .C2(G50gat), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n486));
  XOR2_X1   g285(.A(KEYINPUT14), .B(G29gat), .Z(new_n487));
  OAI21_X1  g286(.A(new_n486), .B1(new_n487), .B2(G36gat), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n488), .A2(new_n482), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT17), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n491), .B(KEYINPUT94), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n493), .B1(new_n494), .B2(new_n492), .ZN(new_n495));
  INV_X1    g294(.A(G8gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT95), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT16), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(G1gat), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(G1gat), .B2(new_n498), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI221_X1 g303(.A(new_n500), .B1(new_n501), .B2(new_n496), .C1(G1gat), .C2(new_n498), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n495), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n506), .A3(KEYINPUT97), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT97), .B1(new_n494), .B2(new_n506), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n508), .B(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT18), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n512), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n516), .A2(new_n510), .B1(new_n495), .B2(new_n507), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT18), .A3(new_n509), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n494), .A2(new_n506), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n511), .B2(new_n512), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n509), .B(KEYINPUT13), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(G197gat), .ZN(new_n525));
  XOR2_X1   g324(.A(KEYINPUT11), .B(G169gat), .Z(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n527), .B(KEYINPUT12), .Z(new_n528));
  NAND2_X1  g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n528), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n515), .A2(new_n518), .A3(new_n530), .A4(new_n522), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n478), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT21), .ZN(new_n534));
  INV_X1    g333(.A(G64gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(G57gat), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(KEYINPUT98), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(KEYINPUT98), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(G64gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  OR2_X1    g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT9), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n539), .A2(G64gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT9), .B1(new_n536), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(new_n541), .A3(new_n542), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n507), .B1(new_n534), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT99), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n534), .ZN(new_n552));
  NAND2_X1  g351(.A1(G231gat), .A2(G233gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G127gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n551), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(new_n217), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT7), .ZN(new_n567));
  NAND2_X1  g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  INV_X1    g367(.A(G85gat), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G99gat), .B(G106gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n494), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577));
  AND2_X1   g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n576), .A2(new_n577), .B1(KEYINPUT41), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n574), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n495), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n576), .A2(new_n577), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n578), .A2(KEYINPUT41), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n580), .B(new_n582), .C1(new_n577), .C2(new_n576), .ZN(new_n589));
  AND3_X1   g388(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n588), .B1(new_n585), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n565), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n549), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT10), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n574), .A2(new_n545), .A3(new_n548), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n574), .A2(KEYINPUT10), .A3(new_n545), .A4(new_n548), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n604), .B(KEYINPUT101), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT102), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608));
  AOI211_X1 g407(.A(new_n608), .B(new_n605), .C1(new_n601), .C2(new_n602), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n598), .A2(new_n600), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(G230gat), .A3(G233gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n597), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n603), .A2(new_n604), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n612), .A3(new_n597), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT103), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT103), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n606), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n608), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n603), .A2(KEYINPUT102), .A3(new_n606), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n620), .A2(new_n612), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n618), .B(new_n615), .C1(new_n622), .C2(new_n597), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n594), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n533), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n270), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G1gat), .ZN(G1324gat));
  INV_X1    g428(.A(new_n627), .ZN(new_n630));
  INV_X1    g429(.A(new_n362), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n632), .A2(KEYINPUT104), .A3(new_n496), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT104), .B1(new_n632), .B2(new_n496), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT42), .ZN(new_n635));
  XOR2_X1   g434(.A(KEYINPUT16), .B(G8gat), .Z(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n633), .B(new_n634), .C1(new_n637), .C2(new_n638), .ZN(G1325gat));
  OR3_X1    g438(.A1(new_n630), .A2(G15gat), .A3(new_n473), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT105), .B1(new_n467), .B2(new_n461), .ZN(new_n641));
  INV_X1    g440(.A(new_n456), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n441), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT75), .B1(new_n644), .B2(new_n459), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n466), .A4(new_n462), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT106), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(G15gat), .B1(new_n630), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n640), .A2(new_n651), .ZN(G1326gat));
  NAND2_X1  g451(.A1(new_n627), .A2(new_n472), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT43), .B(G22gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  INV_X1    g454(.A(new_n624), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n564), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n533), .A2(new_n593), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n485), .A3(new_n270), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT45), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n641), .A2(new_n430), .A3(new_n647), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(new_n477), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(new_n592), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n478), .A2(KEYINPUT44), .A3(new_n592), .ZN(new_n666));
  INV_X1    g465(.A(new_n532), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n657), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n270), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n660), .A2(new_n671), .ZN(G1328gat));
  INV_X1    g471(.A(new_n658), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(G36gat), .A3(new_n631), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT46), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n669), .A2(new_n676), .A3(new_n631), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n676), .B1(new_n669), .B2(new_n631), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G36gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n675), .B1(new_n677), .B2(new_n679), .ZN(G1329gat));
  NOR2_X1   g479(.A1(new_n473), .A2(new_n483), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n658), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(KEYINPUT47), .ZN(new_n683));
  INV_X1    g482(.A(new_n648), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n483), .B1(new_n669), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(KEYINPUT109), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n483), .B1(new_n669), .B2(new_n650), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(new_n682), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n690));
  OAI22_X1  g489(.A1(new_n686), .A2(new_n687), .B1(new_n689), .B2(new_n690), .ZN(G1330gat));
  OAI21_X1  g490(.A(G50gat), .B1(new_n669), .B2(new_n469), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n658), .A2(new_n392), .A3(new_n472), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT48), .Z(G1331gat));
  NOR3_X1   g494(.A1(new_n594), .A2(new_n656), .A3(new_n532), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n662), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n670), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(new_n539), .ZN(G1332gat));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n631), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT49), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n535), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT49), .B(G64gat), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT110), .Z(G1333gat));
  INV_X1    g504(.A(G71gat), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n650), .A2(new_n697), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n706), .B1(new_n697), .B2(new_n473), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT50), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n709), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(G1334gat));
  NOR2_X1   g514(.A1(new_n697), .A2(new_n469), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g516(.A1(new_n565), .A2(new_n532), .A3(new_n656), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n665), .A2(new_n666), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G85gat), .B1(new_n719), .B2(new_n670), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n565), .A2(new_n532), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n662), .A2(new_n592), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n662), .A2(KEYINPUT51), .A3(new_n592), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n270), .A2(new_n624), .A3(new_n569), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n720), .B1(new_n727), .B2(new_n728), .ZN(G1336gat));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730));
  OAI21_X1  g529(.A(G92gat), .B1(new_n719), .B2(new_n631), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n631), .A2(new_n656), .A3(G92gat), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n726), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n726), .B2(new_n733), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n730), .B(new_n731), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n722), .A2(KEYINPUT113), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n725), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT113), .B1(new_n722), .B2(new_n739), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n733), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n731), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n737), .B1(new_n744), .B2(KEYINPUT52), .ZN(new_n745));
  AOI211_X1 g544(.A(KEYINPUT114), .B(new_n730), .C1(new_n743), .C2(new_n731), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n736), .B1(new_n745), .B2(new_n746), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n719), .B2(new_n650), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n473), .A2(G99gat), .A3(new_n656), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n727), .B2(new_n749), .ZN(G1338gat));
  OR2_X1    g549(.A1(new_n719), .A2(new_n469), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G106gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n469), .A2(G106gat), .A3(new_n656), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT53), .B1(new_n726), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n741), .A2(new_n742), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n756), .A2(new_n753), .B1(new_n751), .B2(G106gat), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n757), .B2(new_n758), .ZN(G1339gat));
  NAND4_X1  g558(.A1(new_n565), .A2(new_n667), .A3(new_n593), .A4(new_n656), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n517), .A2(new_n509), .B1(new_n520), .B2(new_n521), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762));
  AND3_X1   g561(.A1(new_n761), .A2(new_n762), .A3(new_n527), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n762), .B1(new_n761), .B2(new_n527), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n531), .A3(new_n592), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n767), .B1(new_n607), .B2(new_n609), .ZN(new_n768));
  INV_X1    g567(.A(new_n597), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n614), .B(KEYINPUT54), .C1(new_n603), .C2(new_n606), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n768), .A2(KEYINPUT55), .A3(new_n769), .A4(new_n770), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n773), .A2(new_n615), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT116), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n773), .A2(new_n777), .A3(new_n615), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n766), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n527), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT117), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n761), .A2(new_n762), .A3(new_n527), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n624), .A2(new_n782), .A3(new_n531), .A4(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT118), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n765), .A2(KEYINPUT118), .A3(new_n531), .A4(new_n624), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n532), .A2(new_n776), .A3(new_n778), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n780), .B1(new_n789), .B2(new_n593), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n760), .B1(new_n790), .B2(new_n565), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n791), .A2(new_n270), .A3(new_n631), .A4(new_n474), .ZN(new_n792));
  INV_X1    g591(.A(G113gat), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n792), .A2(new_n793), .A3(new_n667), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n791), .A2(new_n270), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n472), .A2(new_n644), .A3(new_n464), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(new_n631), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n532), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n794), .B1(new_n800), .B2(new_n793), .ZN(G1340gat));
  INV_X1    g600(.A(G120gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n792), .A2(new_n802), .A3(new_n656), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n799), .A2(new_n624), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n802), .ZN(G1341gat));
  OAI21_X1  g604(.A(G127gat), .B1(new_n792), .B2(new_n564), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n565), .A2(new_n555), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n798), .B2(new_n807), .ZN(G1342gat));
  OR3_X1    g607(.A1(new_n798), .A2(G134gat), .A3(new_n593), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n810));
  OAI21_X1  g609(.A(G134gat), .B1(new_n792), .B2(new_n593), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(KEYINPUT56), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(G1343gat));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n791), .A2(new_n814), .A3(new_n270), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n791), .B2(new_n270), .ZN(new_n816));
  NOR4_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n362), .A4(new_n469), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n667), .A2(G141gat), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n650), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n648), .A2(new_n670), .A3(new_n362), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n775), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n775), .A2(new_n822), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n532), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n592), .B1(new_n825), .B2(new_n784), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n780), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n565), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n760), .ZN(new_n830));
  OAI211_X1 g629(.A(KEYINPUT57), .B(new_n472), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n791), .B2(new_n472), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g633(.A(KEYINPUT119), .B(KEYINPUT57), .C1(new_n791), .C2(new_n472), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n532), .B(new_n821), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT124), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(G141gat), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n836), .A2(KEYINPUT124), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n819), .B(new_n820), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n836), .A2(G141gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n819), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n841), .B1(new_n843), .B2(KEYINPUT58), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  AOI211_X1 g644(.A(KEYINPUT122), .B(new_n845), .C1(new_n842), .C2(new_n819), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n844), .B2(new_n846), .ZN(G1344gat));
  NAND2_X1  g646(.A1(new_n817), .A2(new_n650), .ZN(new_n848));
  OR3_X1    g647(.A1(new_n848), .A2(new_n214), .A3(new_n656), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n821), .B1(new_n834), .B2(new_n835), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(new_n656), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n214), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n791), .A2(new_n472), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT125), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n766), .A2(new_n775), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n564), .B1(new_n826), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n469), .B1(new_n858), .B2(new_n760), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n859), .B2(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT57), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n624), .A3(new_n821), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n852), .B1(new_n864), .B2(G148gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n849), .B1(new_n853), .B2(new_n865), .ZN(G1345gat));
  OR3_X1    g665(.A1(new_n850), .A2(new_n217), .A3(new_n564), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n848), .A2(new_n564), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(KEYINPUT126), .ZN(new_n870));
  AOI21_X1  g669(.A(G155gat), .B1(new_n869), .B2(KEYINPUT126), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(G1346gat));
  OAI21_X1  g671(.A(G162gat), .B1(new_n850), .B2(new_n593), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n592), .A2(new_n218), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n848), .B2(new_n874), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n631), .A2(new_n270), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n791), .A2(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n796), .ZN(new_n878));
  AOI21_X1  g677(.A(G169gat), .B1(new_n878), .B2(new_n532), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n474), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(new_n284), .A3(new_n667), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(G1348gat));
  AOI21_X1  g681(.A(G176gat), .B1(new_n878), .B2(new_n624), .ZN(new_n883));
  INV_X1    g682(.A(new_n880), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n624), .A2(new_n319), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(G1349gat));
  NAND3_X1  g685(.A1(new_n878), .A2(new_n275), .A3(new_n565), .ZN(new_n887));
  OAI21_X1  g686(.A(G183gat), .B1(new_n880), .B2(new_n564), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n878), .A2(new_n272), .A3(new_n592), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT127), .Z(new_n892));
  OAI21_X1  g691(.A(G190gat), .B1(new_n880), .B2(new_n593), .ZN(new_n893));
  XNOR2_X1  g692(.A(new_n893), .B(KEYINPUT61), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1351gat));
  INV_X1    g694(.A(G197gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n650), .A2(new_n876), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n532), .A3(new_n854), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n861), .B2(new_n862), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n667), .A2(new_n896), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n896), .A2(new_n899), .B1(new_n900), .B2(new_n901), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n854), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n656), .A2(G204gat), .ZN(new_n904));
  OR3_X1    g703(.A1(new_n903), .A2(KEYINPUT62), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n863), .A2(new_n624), .A3(new_n898), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G204gat), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT62), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(G1353gat));
  OR3_X1    g708(.A1(new_n903), .A2(G211gat), .A3(new_n564), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n900), .A2(new_n565), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n911), .B2(G211gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1354gat));
  NAND2_X1  g713(.A1(new_n900), .A2(new_n592), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G218gat), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n593), .A2(G218gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n903), .B2(new_n917), .ZN(G1355gat));
endmodule


