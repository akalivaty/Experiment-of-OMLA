//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978, new_n979, new_n980;
  XOR2_X1   g000(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT91), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G141gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G169gat), .B(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT12), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(G1gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(G1gat), .B2(new_n210), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n217));
  AOI21_X1  g016(.A(G36gat), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n219), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT93), .ZN(new_n227));
  INV_X1    g026(.A(G50gat), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n227), .A2(new_n228), .A3(G43gat), .ZN(new_n229));
  AOI211_X1 g028(.A(KEYINPUT15), .B(new_n229), .C1(new_n227), .C2(new_n224), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n223), .A2(new_n225), .B1(new_n230), .B2(new_n221), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(KEYINPUT17), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n226), .A2(new_n231), .A3(KEYINPUT17), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n215), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n215), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n231), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT94), .B1(new_n242), .B2(new_n215), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n238), .A2(new_n243), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n236), .B(KEYINPUT13), .Z(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n241), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n239), .A2(new_n240), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n209), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n239), .A2(new_n240), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n252), .A2(new_n208), .A3(new_n248), .A4(new_n241), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT95), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n255), .B(new_n209), .C1(new_n249), .C2(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G228gat), .A2(G233gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT85), .Z(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT79), .B(G155gat), .ZN(new_n260));
  INV_X1    g059(.A(G162gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT2), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G141gat), .B(G148gat), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(G155gat), .ZN(new_n264));
  INV_X1    g063(.A(G155gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G162gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT78), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n266), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT78), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n262), .A2(new_n263), .A3(new_n267), .A4(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n268), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n277));
  NAND2_X1  g076(.A1(G211gat), .A2(G218gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT22), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n282), .A3(new_n279), .ZN(new_n283));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G211gat), .ZN(new_n286));
  INV_X1    g085(.A(G218gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n278), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT29), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(new_n289), .B2(new_n285), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n276), .B1(new_n277), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n289), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n295), .A2(new_n281), .A3(new_n283), .A4(new_n284), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n294), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n270), .A2(new_n267), .A3(new_n263), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT79), .B(G155gat), .Z(new_n300));
  AOI21_X1  g099(.A(new_n272), .B1(new_n300), .B2(G162gat), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n274), .B(new_n277), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n259), .B1(new_n292), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n303), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n296), .A2(new_n297), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n258), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT29), .B1(new_n296), .B2(new_n297), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n275), .B1(new_n309), .B2(KEYINPUT3), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n308), .A2(KEYINPUT86), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT86), .B1(new_n308), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n305), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G22gat), .ZN(new_n314));
  INV_X1    g113(.A(G22gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n315), .B(new_n305), .C1(new_n311), .C2(new_n312), .ZN(new_n316));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT31), .B(G50gat), .ZN(new_n318));
  XOR2_X1   g117(.A(new_n317), .B(new_n318), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT88), .A4(new_n320), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT87), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n314), .A2(new_n316), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n319), .ZN(new_n328));
  AOI211_X1 g127(.A(KEYINPUT87), .B(new_n320), .C1(new_n314), .C2(new_n316), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n323), .A2(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT35), .ZN(new_n331));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(G169gat), .A2(G176gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT23), .ZN(new_n337));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(G169gat), .B2(G176gat), .ZN(new_n340));
  AND4_X1   g139(.A1(KEYINPUT25), .A2(new_n337), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(KEYINPUT64), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n342), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  NAND3_X1  g146(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT65), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  INV_X1    g150(.A(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT65), .B1(new_n353), .B2(new_n348), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n341), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n344), .A2(new_n348), .A3(new_n353), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(KEYINPUT27), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT27), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G183gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(new_n364), .A3(new_n352), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT27), .B(G183gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT28), .A3(new_n352), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n336), .A2(KEYINPUT26), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n342), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n338), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(new_n336), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n360), .A2(new_n361), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n361), .B1(new_n360), .B2(new_n377), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT66), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n377), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT66), .A3(new_n376), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n360), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n383), .B1(new_n387), .B2(new_n303), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n381), .A2(new_n383), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n387), .A2(new_n303), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT76), .B1(new_n391), .B2(new_n383), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n298), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n380), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n394), .A2(new_n303), .A3(new_n382), .A4(new_n378), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n387), .A2(new_n382), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n307), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n335), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n388), .A2(new_n389), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n394), .A2(new_n383), .A3(new_n378), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n388), .A2(new_n389), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n307), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n397), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n334), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n398), .A2(KEYINPUT30), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n392), .A2(new_n400), .A3(new_n399), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n397), .B1(new_n407), .B2(new_n307), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n409), .A3(new_n334), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n330), .A2(new_n331), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n413));
  AND2_X1   g212(.A1(G113gat), .A2(G120gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(G113gat), .A2(G120gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G113gat), .ZN(new_n417));
  INV_X1    g216(.A(G120gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G113gat), .A2(G120gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(KEYINPUT67), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G127gat), .ZN(new_n424));
  INV_X1    g223(.A(G134gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(G127gat), .A2(G134gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT68), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n414), .B2(new_n415), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n419), .A2(KEYINPUT68), .A3(new_n420), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(G127gat), .A2(G134gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(G127gat), .A2(G134gat), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT69), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n426), .A2(new_n437), .A3(new_n427), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  AND4_X1   g238(.A1(new_n429), .A2(new_n433), .A3(new_n439), .A4(new_n422), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT1), .B1(new_n436), .B2(new_n438), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n429), .B1(new_n441), .B2(new_n433), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n428), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n443), .A2(new_n360), .A3(new_n385), .A4(new_n386), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT69), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n437), .B1(new_n426), .B2(new_n427), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n422), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n431), .A2(new_n432), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT70), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n441), .A2(new_n429), .A3(new_n433), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n387), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(G227gat), .A2(G233gat), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n444), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(G15gat), .B(G43gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  OR2_X1    g257(.A1(new_n458), .A2(KEYINPUT72), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(KEYINPUT72), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(KEYINPUT33), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(KEYINPUT32), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n458), .B1(new_n455), .B2(KEYINPUT32), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n455), .A2(KEYINPUT71), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT71), .B1(new_n455), .B2(new_n464), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n454), .B1(new_n444), .B2(new_n453), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT34), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI211_X1 g270(.A(KEYINPUT34), .B(new_n454), .C1(new_n444), .C2(new_n453), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT73), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n473), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n468), .A2(KEYINPUT73), .A3(new_n474), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n440), .A2(new_n442), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n428), .A2(new_n271), .A3(new_n274), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n482), .A2(KEYINPUT4), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n428), .A2(new_n271), .A3(new_n274), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n450), .A2(new_n451), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT3), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n302), .B1(new_n276), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n492), .B2(new_n452), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT5), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT81), .B1(new_n452), .B2(new_n276), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n443), .A2(new_n496), .A3(new_n275), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n486), .A2(new_n487), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT4), .B1(new_n482), .B2(new_n483), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n485), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT83), .ZN(new_n504));
  INV_X1    g303(.A(new_n490), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n491), .B1(new_n271), .B2(new_n274), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n506), .B1(new_n276), .B2(new_n277), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n507), .B2(new_n443), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT83), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n488), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n504), .A2(new_n508), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(G1gat), .B(G29gat), .Z(new_n513));
  XNOR2_X1  g312(.A(G57gat), .B(G85gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n515), .B(new_n516), .Z(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n481), .B1(new_n501), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n443), .B(new_n302), .C1(new_n491), .C2(new_n276), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n520), .B(new_n490), .C1(new_n484), .C2(new_n488), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n495), .A2(new_n497), .B1(new_n487), .B2(new_n486), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n521), .B(KEYINPUT5), .C1(new_n522), .C2(new_n490), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n517), .B1(new_n523), .B2(new_n512), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT89), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n512), .B1(new_n494), .B2(new_n500), .ZN(new_n526));
  INV_X1    g325(.A(new_n517), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n523), .A2(new_n512), .A3(new_n517), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n528), .A2(new_n529), .A3(new_n481), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(KEYINPUT6), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n480), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n412), .A2(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n475), .A2(new_n477), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(new_n519), .B2(new_n524), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n528), .A2(KEYINPUT84), .A3(new_n481), .A4(new_n530), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n539), .A3(new_n532), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n330), .A2(new_n536), .A3(new_n540), .A4(new_n411), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n452), .A2(KEYINPUT81), .A3(new_n276), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n496), .B1(new_n443), .B2(new_n275), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n499), .B(new_n490), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT39), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n504), .A2(new_n511), .A3(new_n520), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n505), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT39), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n550), .A3(new_n505), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n517), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT40), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n548), .A2(new_n505), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT39), .A3(new_n546), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT40), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n517), .A4(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(new_n528), .A3(new_n410), .A4(new_n406), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n298), .B1(new_n401), .B2(new_n402), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n395), .A2(new_n396), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n307), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT38), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n334), .B1(new_n403), .B2(new_n404), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n334), .A2(new_n561), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n524), .A2(KEYINPUT6), .B1(new_n408), .B2(new_n334), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n525), .A2(new_n567), .A3(new_n531), .A4(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT38), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n334), .B1(new_n408), .B2(new_n561), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT37), .B1(new_n393), .B2(new_n397), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n559), .B(new_n330), .C1(new_n569), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n540), .A2(new_n411), .ZN(new_n575));
  INV_X1    g374(.A(new_n328), .ZN(new_n576));
  INV_X1    g375(.A(new_n329), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n321), .A2(new_n322), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n576), .A2(new_n577), .B1(new_n578), .B2(new_n324), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n478), .A2(new_n581), .A3(new_n479), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n475), .A2(KEYINPUT36), .A3(new_n477), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n574), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n257), .B1(new_n543), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT96), .B(G57gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  INV_X1    g388(.A(G64gat), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n589), .B1(G57gat), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  OR2_X1    g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n592), .B(new_n596), .C1(KEYINPUT97), .C2(new_n588), .ZN(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n593), .B(new_n594), .C1(new_n598), .C2(new_n595), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT21), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(G127gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n215), .B1(new_n601), .B2(new_n600), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT98), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(G155gat), .ZN(new_n610));
  XOR2_X1   g409(.A(G183gat), .B(G211gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n597), .A2(new_n599), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT10), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT8), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n624), .B2(new_n623), .ZN(new_n626));
  INV_X1    g425(.A(G92gat), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n627), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n628));
  OAI21_X1  g427(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n626), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G99gat), .B(G106gat), .Z(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(KEYINPUT100), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n621), .A2(KEYINPUT101), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n619), .A2(new_n633), .A3(new_n634), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT10), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n636), .A2(new_n600), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n638), .A2(new_n635), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT101), .B1(new_n645), .B2(new_n621), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n618), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n642), .ZN(new_n648));
  INV_X1    g447(.A(new_n618), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(KEYINPUT102), .A3(new_n649), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  AND2_X1   g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n647), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(KEYINPUT103), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(KEYINPUT103), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n656), .B1(new_n647), .B2(new_n650), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n233), .A2(new_n234), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n645), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n645), .A2(new_n232), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n667));
  NAND2_X1  g466(.A1(G232gat), .A2(G233gat), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(G190gat), .B(G218gat), .Z(new_n670));
  OR3_X1    g469(.A1(new_n665), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n665), .B2(new_n669), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n668), .A2(new_n667), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n671), .A2(new_n676), .A3(new_n672), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n617), .A2(new_n663), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n586), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n538), .A2(new_n539), .A3(new_n532), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT105), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT104), .B(G1gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1324gat));
  INV_X1    g488(.A(new_n411), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT16), .B(G8gat), .Z(new_n691));
  NAND3_X1  g490(.A1(new_n684), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n694), .A2(KEYINPUT106), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(KEYINPUT106), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n214), .B1(new_n684), .B2(new_n690), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n692), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(new_n696), .B2(new_n698), .ZN(G1325gat));
  OAI21_X1  g498(.A(G15gat), .B1(new_n683), .B2(new_n584), .ZN(new_n700));
  INV_X1    g499(.A(new_n480), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(G15gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n683), .B2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n683), .A2(new_n330), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  INV_X1    g505(.A(new_n663), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n586), .A2(new_n617), .A3(new_n681), .A4(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(G29gat), .A3(new_n540), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n412), .A2(new_n534), .B1(new_n541), .B2(KEYINPUT35), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n585), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g514(.A1(new_n575), .A2(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(KEYINPUT108), .A3(new_n574), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n712), .B1(new_n718), .B2(new_n680), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n543), .A2(new_n585), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(KEYINPUT44), .A3(new_n681), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n663), .A2(new_n257), .A3(new_n616), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G29gat), .B1(new_n724), .B2(new_n540), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n711), .A2(new_n725), .ZN(G1328gat));
  NOR3_X1   g525(.A1(new_n708), .A2(G36gat), .A3(new_n411), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT46), .ZN(new_n728));
  OAI21_X1  g527(.A(G36gat), .B1(new_n724), .B2(new_n411), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(G1329gat));
  INV_X1    g529(.A(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n708), .B2(new_n701), .ZN(new_n732));
  INV_X1    g531(.A(new_n584), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G43gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n732), .B1(new_n724), .B2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1330gat));
  OAI21_X1  g536(.A(new_n228), .B1(new_n708), .B2(new_n330), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n579), .A2(G50gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n724), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g540(.A1(new_n663), .A2(new_n257), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n718), .A2(new_n617), .A3(new_n681), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n685), .B(KEYINPUT110), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g545(.A(new_n746), .B(new_n587), .Z(G1332gat));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n690), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT49), .B(G64gat), .Z(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(G1333gat));
  NAND2_X1  g550(.A1(new_n743), .A2(new_n733), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n701), .A2(G71gat), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n752), .A2(G71gat), .B1(new_n743), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n743), .A2(new_n579), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n616), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n722), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n540), .ZN(new_n761));
  AND4_X1   g560(.A1(KEYINPUT108), .A2(new_n574), .A3(new_n580), .A4(new_n584), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT108), .B1(new_n716), .B2(new_n574), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n543), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n617), .A2(new_n257), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n764), .A2(new_n681), .A3(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT112), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n764), .A2(KEYINPUT112), .A3(new_n681), .A4(new_n767), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n770), .A2(KEYINPUT113), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n764), .A2(new_n257), .A3(new_n617), .A4(new_n681), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n766), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT113), .B1(new_n770), .B2(new_n771), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n707), .A2(G85gat), .A3(new_n540), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n761), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  NAND3_X1  g578(.A1(new_n663), .A2(new_n627), .A3(new_n690), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n772), .A2(new_n774), .ZN(new_n781));
  INV_X1    g580(.A(new_n776), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n719), .A2(new_n690), .A3(new_n721), .A4(new_n759), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n771), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n718), .A2(new_n680), .A3(new_n765), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n790));
  OAI21_X1  g589(.A(KEYINPUT115), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT115), .ZN(new_n792));
  INV_X1    g591(.A(new_n790), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n773), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n788), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n780), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n795), .A2(new_n796), .B1(G92gat), .B2(new_n784), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n783), .A2(new_n787), .B1(new_n797), .B2(new_n786), .ZN(G1337gat));
  NOR3_X1   g597(.A1(new_n707), .A2(new_n701), .A3(G99gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n775), .B2(new_n776), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n760), .B2(new_n584), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G99gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n760), .A2(new_n801), .A3(new_n584), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n800), .B1(new_n803), .B2(new_n804), .ZN(G1338gat));
  NOR3_X1   g604(.A1(new_n707), .A2(G106gat), .A3(new_n330), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(new_n781), .B2(new_n782), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n719), .A2(new_n579), .A3(new_n721), .A4(new_n759), .ZN(new_n809));
  XNOR2_X1  g608(.A(KEYINPUT117), .B(G106gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n795), .A2(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n808), .A2(new_n813), .B1(new_n814), .B2(new_n812), .ZN(G1339gat));
  AND2_X1   g614(.A1(new_n254), .A2(new_n256), .ZN(new_n816));
  INV_X1    g615(.A(new_n656), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n647), .B2(KEYINPUT54), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n645), .A2(new_n621), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT101), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n821), .A2(new_n649), .A3(new_n643), .A4(new_n639), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(KEYINPUT54), .A3(new_n647), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT118), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n822), .A2(new_n647), .A3(new_n825), .A4(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n818), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n661), .B1(new_n827), .B2(KEYINPUT55), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n827), .A2(KEYINPUT55), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n816), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n246), .A2(new_n247), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n236), .B1(new_n235), .B2(new_n238), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n207), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n253), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n663), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n681), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n828), .A2(new_n829), .A3(new_n681), .A4(new_n834), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n617), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n682), .A2(new_n257), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n330), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n685), .A2(new_n411), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n842), .A2(new_n701), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n257), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n744), .B1(new_n839), .B2(new_n840), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n330), .A2(new_n536), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n847), .A2(new_n411), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n816), .A2(new_n417), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n846), .A2(new_n853), .ZN(G1340gat));
  AOI21_X1  g653(.A(G120gat), .B1(new_n850), .B2(new_n663), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n707), .A2(new_n418), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n844), .B2(new_n856), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n845), .B2(new_n617), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n850), .A2(new_n424), .A3(new_n616), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  OAI21_X1  g659(.A(G134gat), .B1(new_n845), .B2(new_n680), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n680), .A2(new_n690), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n425), .A3(new_n849), .A4(new_n862), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT120), .B1(new_n863), .B2(KEYINPUT56), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n863), .A2(KEYINPUT120), .A3(KEYINPUT56), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n861), .B(new_n864), .C1(new_n865), .C2(new_n866), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n733), .A2(new_n843), .ZN(new_n868));
  INV_X1    g667(.A(G141gat), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n257), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n841), .B2(new_n579), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n872), .B(new_n330), .C1(new_n839), .C2(new_n840), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n868), .B(new_n870), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n733), .A2(new_n330), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n847), .A2(new_n411), .A3(new_n816), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n869), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n874), .A2(KEYINPUT58), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1344gat));
  AND2_X1   g681(.A1(new_n847), .A2(new_n875), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(new_n411), .ZN(new_n884));
  INV_X1    g683(.A(G148gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n663), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n663), .B(new_n868), .C1(new_n871), .C2(new_n873), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n887), .A2(new_n888), .A3(G148gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n887), .B2(G148gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1345gat));
  NAND3_X1  g690(.A1(new_n884), .A2(new_n260), .A3(new_n616), .ZN(new_n892));
  INV_X1    g691(.A(new_n840), .ZN(new_n893));
  INV_X1    g692(.A(new_n661), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n824), .A2(new_n826), .ZN(new_n895));
  INV_X1    g694(.A(new_n818), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(KEYINPUT55), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n827), .A2(KEYINPUT55), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n898), .A2(new_n257), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n663), .A2(new_n834), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n680), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n837), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n893), .B1(new_n903), .B2(new_n617), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n872), .B1(new_n904), .B2(new_n330), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n841), .A2(KEYINPUT57), .A3(new_n579), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(new_n616), .A3(new_n868), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n892), .B1(new_n908), .B2(new_n260), .ZN(G1346gat));
  INV_X1    g708(.A(KEYINPUT121), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n907), .A2(new_n910), .A3(new_n681), .A4(new_n868), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n681), .B(new_n868), .C1(new_n871), .C2(new_n873), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT121), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n913), .A3(G162gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n883), .A2(new_n261), .A3(new_n862), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1347gat));
  NOR2_X1   g715(.A1(new_n904), .A2(new_n685), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n848), .A2(new_n411), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n816), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n744), .A2(new_n690), .A3(new_n480), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT122), .Z(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n330), .A3(new_n841), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n816), .A2(G169gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n923), .B2(new_n707), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n707), .A2(G176gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n917), .A2(new_n918), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(G1349gat));
  NAND4_X1  g731(.A1(new_n917), .A2(new_n368), .A3(new_n616), .A4(new_n918), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n923), .A2(new_n617), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n934), .B2(new_n351), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n933), .B(new_n937), .C1(new_n934), .C2(new_n351), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n352), .A3(new_n681), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n681), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(G190gat), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT61), .B(new_n352), .C1(new_n924), .C2(new_n681), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n745), .A2(new_n411), .A3(new_n733), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n907), .A2(new_n946), .A3(new_n816), .A4(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n816), .B(new_n947), .C1(new_n871), .C2(new_n873), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n948), .A2(new_n950), .A3(G197gat), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n733), .A2(new_n411), .A3(new_n330), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n917), .A2(new_n952), .ZN(new_n953));
  OR3_X1    g752(.A1(new_n953), .A2(G197gat), .A3(new_n257), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n954), .ZN(G1352gat));
  NAND4_X1  g754(.A1(new_n907), .A2(KEYINPUT125), .A3(new_n663), .A4(new_n947), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n663), .B(new_n947), .C1(new_n871), .C2(new_n873), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n956), .A2(new_n959), .A3(G204gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n707), .A2(G204gat), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT62), .B1(new_n953), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n917), .A2(new_n964), .A3(new_n952), .A4(new_n961), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n960), .A2(new_n966), .ZN(G1353gat));
  INV_X1    g766(.A(new_n953), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n286), .A3(new_n616), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n616), .B(new_n947), .C1(new_n871), .C2(new_n873), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n286), .B1(KEYINPUT126), .B2(new_n971), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n972), .B1(new_n970), .B2(new_n973), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  AOI21_X1  g775(.A(G218gat), .B1(new_n968), .B2(new_n681), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n907), .A2(new_n947), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n680), .A2(new_n287), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT127), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n977), .B1(new_n978), .B2(new_n980), .ZN(G1355gat));
endmodule


