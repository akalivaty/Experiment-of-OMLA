//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT64), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207));
  INV_X1    g006(.A(G120gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G113gat), .ZN(new_n209));
  INV_X1    g008(.A(G113gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G120gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT1), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT68), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G127gat), .B(G134gat), .Z(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n207), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n215), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT27), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT27), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(G190gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT28), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT28), .A4(new_n225), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  OR3_X1    g032(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n233), .A2(new_n234), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n230), .A2(KEYINPUT66), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT66), .B1(new_n230), .B2(new_n235), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT24), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(G183gat), .B(G190gat), .ZN(new_n241));
  OAI211_X1 g040(.A(KEYINPUT65), .B(new_n240), .C1(new_n241), .C2(new_n239), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n240), .B1(new_n241), .B2(new_n239), .ZN(new_n244));
  INV_X1    g043(.A(G169gat), .ZN(new_n245));
  INV_X1    g044(.A(G176gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT23), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n249), .A3(new_n232), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n242), .B(new_n243), .C1(new_n244), .C2(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n239), .A2(G183gat), .A3(G190gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n221), .A2(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n225), .A2(G183gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n255), .B2(KEYINPUT24), .ZN(new_n256));
  INV_X1    g055(.A(new_n250), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n256), .B(new_n257), .C1(KEYINPUT65), .C2(KEYINPUT25), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n220), .B1(new_n238), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT27), .B(G183gat), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT28), .B1(new_n262), .B2(new_n225), .ZN(new_n263));
  INV_X1    g062(.A(new_n229), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n234), .A2(new_n232), .A3(new_n231), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n266), .B1(new_n221), .B2(new_n225), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n261), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n230), .A2(KEYINPUT66), .A3(new_n235), .ZN(new_n269));
  AND4_X1   g068(.A1(new_n220), .A2(new_n259), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n206), .B1(new_n260), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n204), .B1(new_n271), .B2(KEYINPUT32), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n273));
  INV_X1    g072(.A(new_n206), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n268), .A3(new_n269), .ZN(new_n275));
  INV_X1    g074(.A(new_n220), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n220), .A2(new_n259), .A3(new_n268), .A4(new_n269), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n273), .B1(new_n279), .B2(KEYINPUT33), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT33), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n271), .A2(KEYINPUT69), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n272), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n271), .B(KEYINPUT32), .C1(new_n281), .C2(new_n204), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(new_n274), .A3(new_n278), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n287), .A2(KEYINPUT34), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n283), .A2(new_n284), .A3(new_n291), .A4(new_n289), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G22gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G141gat), .ZN(new_n302));
  INV_X1    g101(.A(G141gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(G148gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n297), .B(new_n300), .C1(new_n305), .C2(KEYINPUT2), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n297), .B1(new_n300), .B2(KEYINPUT2), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT75), .B1(new_n301), .B2(G141gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(new_n303), .B2(G148gat), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n301), .A2(KEYINPUT75), .A3(G141gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  INV_X1    g116(.A(G211gat), .ZN(new_n318));
  INV_X1    g117(.A(G218gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(KEYINPUT22), .B2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G211gat), .B(G218gat), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n321), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G228gat), .ZN(new_n326));
  INV_X1    g125(.A(G233gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n313), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n306), .A2(new_n311), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n325), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n321), .B(new_n322), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(new_n314), .B2(new_n315), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n330), .B(KEYINPUT76), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n315), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n313), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n296), .B(new_n332), .C1(new_n339), .C2(new_n328), .ZN(new_n340));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT31), .B(G50gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n335), .B1(new_n313), .B2(new_n337), .ZN(new_n346));
  OAI22_X1  g145(.A1(new_n346), .A2(new_n334), .B1(new_n326), .B2(new_n327), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n296), .B1(new_n347), .B2(new_n332), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT79), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n339), .A2(new_n328), .ZN(new_n350));
  INV_X1    g149(.A(new_n332), .ZN(new_n351));
  OAI21_X1  g150(.A(G22gat), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n344), .A4(new_n340), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n347), .A2(KEYINPUT78), .A3(new_n296), .A4(new_n332), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n352), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n343), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n355), .A2(KEYINPUT80), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT80), .B1(new_n355), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n295), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n335), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n364));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n276), .A2(new_n314), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n220), .A2(new_n312), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n364), .A2(new_n365), .A3(new_n367), .A4(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n220), .B(new_n312), .ZN(new_n373));
  INV_X1    g172(.A(new_n365), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n367), .A2(new_n372), .A3(new_n365), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n335), .A2(new_n369), .A3(new_n220), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n368), .A2(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT6), .ZN(new_n384));
  XOR2_X1   g183(.A(G1gat), .B(G29gat), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n383), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n388), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n384), .B1(new_n382), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT77), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OAI22_X1  g193(.A1(new_n392), .A2(KEYINPUT77), .B1(new_n388), .B2(new_n383), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n315), .ZN(new_n397));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n251), .A2(new_n258), .B1(new_n230), .B2(new_n235), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n275), .A2(new_n400), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n324), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n399), .A2(KEYINPUT29), .ZN(new_n404));
  OAI22_X1  g203(.A1(new_n275), .A2(new_n398), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n333), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G8gat), .B(G36gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n411), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n415));
  OR3_X1    g214(.A1(new_n407), .A2(KEYINPUT30), .A3(new_n413), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT35), .B1(new_n363), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n383), .A2(KEYINPUT84), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n382), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n388), .B(KEYINPUT82), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n392), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n389), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n417), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n427), .A2(KEYINPUT35), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n355), .A2(new_n360), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT80), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n293), .A2(KEYINPUT72), .A3(new_n294), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT72), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n285), .A2(new_n436), .A3(new_n292), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(new_n434), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n408), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n413), .B1(new_n407), .B2(KEYINPUT37), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT38), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n402), .B2(new_n333), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n405), .A2(new_n324), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT38), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n427), .A2(new_n412), .A3(new_n445), .A4(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n365), .B1(new_n380), .B2(new_n367), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT39), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n424), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n373), .A2(new_n374), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n455), .A2(KEYINPUT83), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n455), .B2(KEYINPUT83), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n454), .B1(new_n458), .B2(new_n452), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(KEYINPUT40), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n428), .A3(new_n425), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n451), .A2(new_n434), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n435), .A2(new_n463), .A3(new_n437), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT73), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n435), .A2(new_n466), .A3(new_n463), .A4(new_n437), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n293), .A2(KEYINPUT36), .A3(new_n294), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n293), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n294), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n383), .A2(new_n388), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT77), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n474), .B1(new_n426), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n389), .B1(new_n476), .B2(new_n393), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n432), .B(new_n433), .C1(new_n477), .C2(new_n428), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n462), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n478), .A3(KEYINPUT81), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n441), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n484));
  INV_X1    g283(.A(G8gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G1gat), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT16), .ZN(new_n489));
  INV_X1    g288(.A(G1gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT89), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G1gat), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n485), .B(new_n488), .C1(new_n498), .C2(new_n487), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n487), .B1(new_n496), .B2(new_n497), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n486), .A2(new_n490), .ZN(new_n501));
  OAI21_X1  g300(.A(G8gat), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT86), .B(G29gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(G36gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(KEYINPUT87), .A3(G36gat), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(G50gat), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT88), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(G50gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n512), .B2(new_n513), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT15), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n513), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n518), .A2(new_n516), .A3(new_n511), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT14), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT14), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n517), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n525), .B(KEYINPUT85), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n507), .A2(new_n508), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n519), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n531), .B1(new_n527), .B2(new_n530), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n484), .B(new_n503), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(new_n530), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT17), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n537), .A2(new_n532), .B1(new_n502), .B2(new_n499), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT91), .B1(new_n503), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n535), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G197gat), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT11), .B(G169gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n549), .B(KEYINPUT12), .Z(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n541), .A2(KEYINPUT18), .A3(new_n542), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n503), .B(new_n539), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n542), .B(KEYINPUT13), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n545), .A2(new_n551), .A3(new_n552), .A4(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n543), .A2(new_n544), .B1(new_n553), .B2(new_n554), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n551), .B1(new_n558), .B2(new_n552), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G57gat), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n568), .A2(KEYINPUT93), .ZN(new_n570));
  OR3_X1    g369(.A1(new_n565), .A2(KEYINPUT92), .A3(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(KEYINPUT92), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n572), .A3(new_n566), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(new_n568), .B2(KEYINPUT93), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT94), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n570), .A2(new_n575), .A3(new_n573), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n569), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n503), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G127gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n587), .A2(new_n588), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n584), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(new_n589), .A3(new_n583), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G155gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G183gat), .B(G211gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n592), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n592), .B2(new_n594), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G99gat), .B(G106gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT95), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(G85gat), .ZN(new_n607));
  INV_X1    g406(.A(G92gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n603), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n602), .A2(new_n612), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n605), .B(new_n609), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n611), .A2(KEYINPUT96), .A3(new_n615), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n603), .A2(KEYINPUT96), .A3(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n619), .B1(new_n533), .B2(new_n534), .ZN(new_n620));
  AND2_X1   g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n618), .A2(new_n536), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n624), .B(KEYINPUT97), .Z(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n625), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n620), .A2(new_n630), .A3(new_n622), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n626), .B2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT98), .B1(new_n601), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n636), .B(new_n637), .C1(new_n599), .C2(new_n600), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(G230gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(new_n327), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n611), .A2(KEYINPUT99), .A3(new_n615), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n603), .A2(new_n643), .A3(new_n610), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n580), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT100), .B(KEYINPUT10), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n646), .B(new_n647), .C1(new_n580), .C2(new_n618), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n618), .A2(new_n580), .A3(KEYINPUT10), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n641), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n641), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n619), .A2(new_n581), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n646), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n651), .B(new_n660), .C1(new_n659), .C2(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n655), .B1(new_n650), .B2(new_n658), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR4_X1    g462(.A1(new_n483), .A2(new_n561), .A3(new_n639), .A4(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n396), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(new_n490), .ZN(G1324gat));
  NOR2_X1   g465(.A1(new_n664), .A2(new_n417), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(new_n485), .B2(new_n667), .ZN(new_n670));
  MUX2_X1   g469(.A(new_n669), .B(new_n670), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n664), .B2(new_n473), .ZN(new_n672));
  INV_X1    g471(.A(new_n438), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n672), .B1(new_n664), .B2(new_n674), .ZN(G1326gat));
  OR3_X1    g474(.A1(new_n664), .A2(KEYINPUT102), .A3(new_n434), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT102), .B1(new_n664), .B2(new_n434), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  NAND2_X1  g479(.A1(new_n479), .A2(new_n480), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n451), .A2(new_n434), .A3(new_n461), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n482), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n636), .B1(new_n683), .B2(new_n440), .ZN(new_n684));
  INV_X1    g483(.A(new_n601), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(new_n561), .A3(new_n663), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n504), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n477), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT45), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n691), .B(KEYINPUT44), .C1(new_n483), .C2(new_n636), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n683), .A2(new_n440), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(new_n634), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n682), .A2(new_n473), .A3(new_n478), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n636), .B1(new_n440), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n691), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n692), .B(new_n686), .C1(new_n695), .C2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n698), .B1(new_n684), .B2(new_n693), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n702), .A2(new_n703), .A3(new_n692), .A4(new_n686), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n701), .A2(new_n477), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n701), .A2(KEYINPUT105), .A3(new_n477), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n504), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n690), .B1(new_n707), .B2(new_n709), .ZN(G1328gat));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n521), .A3(new_n428), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  AND3_X1   g511(.A1(new_n701), .A2(new_n428), .A3(new_n704), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n521), .B2(new_n713), .ZN(G1329gat));
  OAI21_X1  g513(.A(G43gat), .B1(new_n700), .B2(new_n473), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n687), .A2(new_n510), .A3(new_n438), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(KEYINPUT47), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n716), .ZN(new_n718));
  INV_X1    g517(.A(new_n473), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n701), .A2(new_n719), .A3(new_n704), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n720), .B2(G43gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n717), .B1(new_n721), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  INV_X1    g522(.A(new_n434), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n687), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n702), .A2(new_n724), .A3(new_n692), .A4(new_n686), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G50gat), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n726), .A2(new_n727), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT48), .B(new_n725), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n725), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n701), .A2(new_n724), .A3(new_n704), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n733), .B2(G50gat), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n731), .B1(new_n734), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g534(.A1(new_n440), .A2(new_n696), .ZN(new_n736));
  INV_X1    g535(.A(new_n663), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n639), .A2(new_n560), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n396), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(new_n563), .ZN(G1332gat));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n417), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n739), .B2(new_n473), .ZN(new_n747));
  INV_X1    g546(.A(G71gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n438), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g550(.A1(new_n739), .A2(new_n434), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g552(.A1(new_n697), .A2(KEYINPUT107), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n561), .A3(new_n601), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n697), .A2(KEYINPUT107), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT51), .B1(new_n755), .B2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n737), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n607), .A3(new_n477), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n702), .A2(new_n692), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n685), .A2(new_n560), .A3(new_n737), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n764), .A2(new_n477), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n607), .B2(new_n766), .ZN(G1336gat));
  NOR2_X1   g566(.A1(new_n417), .A2(G92gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n759), .A2(new_n663), .A3(new_n760), .A4(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n702), .A2(new_n428), .A3(new_n692), .A4(new_n765), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n770), .A2(new_n774), .A3(G92gat), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n770), .B2(G92gat), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n663), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n758), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n757), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n778), .B(new_n758), .C1(new_n755), .C2(new_n756), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n777), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n775), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n773), .B1(new_n783), .B2(new_n772), .ZN(G1337gat));
  INV_X1    g583(.A(G99gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n762), .A2(new_n785), .A3(new_n438), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n764), .A2(new_n719), .A3(new_n765), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n785), .B2(new_n787), .ZN(G1338gat));
  NAND4_X1  g587(.A1(new_n702), .A2(new_n724), .A3(new_n692), .A4(new_n765), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n789), .A2(G106gat), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n780), .A2(new_n781), .ZN(new_n791));
  OR3_X1    g590(.A1(new_n434), .A2(G106gat), .A3(new_n737), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT110), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n790), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n761), .B2(new_n792), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n794), .A2(new_n795), .B1(new_n797), .B2(new_n790), .ZN(G1339gat));
  AOI211_X1 g597(.A(KEYINPUT54), .B(new_n641), .C1(new_n648), .C2(new_n649), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT112), .B1(new_n799), .B2(new_n654), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n650), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n655), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n648), .A2(new_n641), .A3(new_n649), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n541), .A2(new_n542), .B1(new_n553), .B2(new_n554), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n549), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n556), .A2(new_n634), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n799), .A2(KEYINPUT112), .A3(new_n654), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n803), .B1(new_n802), .B2(new_n655), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT55), .B(new_n807), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n815), .A2(new_n661), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n812), .A2(new_n816), .A3(KEYINPUT113), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n808), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n560), .A2(new_n816), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n556), .A2(new_n663), .A3(new_n810), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n634), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n601), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n635), .A2(new_n561), .A3(new_n638), .A4(new_n737), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n396), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n363), .A2(new_n428), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n560), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n827), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n724), .A2(new_n673), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n477), .A2(new_n417), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n561), .A2(new_n210), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(G1340gat));
  AOI21_X1  g638(.A(new_n208), .B1(new_n837), .B2(new_n663), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT114), .Z(new_n841));
  NAND3_X1  g640(.A1(new_n831), .A2(new_n208), .A3(new_n663), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1341gat));
  NOR3_X1   g642(.A1(new_n830), .A2(KEYINPUT115), .A3(new_n601), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(G127gat), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT115), .B1(new_n830), .B2(new_n601), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n601), .A2(new_n588), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n845), .A2(new_n846), .B1(new_n837), .B2(new_n847), .ZN(G1342gat));
  NOR2_X1   g647(.A1(new_n636), .A2(G134gat), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n837), .A2(new_n634), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(G134gat), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT116), .B1(new_n850), .B2(KEYINPUT56), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n850), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n853), .B(KEYINPUT117), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n852), .A2(G134gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(KEYINPUT56), .B2(new_n850), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n861), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n719), .A2(new_n836), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n724), .A2(KEYINPUT57), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n661), .B(new_n815), .C1(new_n557), .C2(new_n559), .ZN(new_n865));
  XNOR2_X1  g664(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n866), .B1(new_n805), .B2(new_n807), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n824), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n636), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(KEYINPUT119), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n815), .A2(new_n661), .ZN(new_n872));
  NOR4_X1   g671(.A1(new_n872), .A2(new_n808), .A3(new_n811), .A4(new_n818), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT113), .B1(new_n812), .B2(new_n816), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n875), .B1(new_n870), .B2(KEYINPUT119), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n601), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n864), .B1(new_n877), .B2(new_n827), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n833), .B2(new_n724), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n863), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n561), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n828), .A2(new_n417), .A3(new_n724), .A4(new_n473), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n303), .A3(new_n560), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT58), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT58), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n301), .A2(KEYINPUT59), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n880), .B2(new_n737), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n824), .B1(new_n865), .B2(new_n808), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n636), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n685), .B1(new_n875), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n827), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT57), .B(new_n724), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT121), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT121), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n833), .A2(new_n898), .A3(KEYINPUT57), .A4(new_n724), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n685), .B1(new_n869), .B2(new_n817), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n724), .B1(new_n900), .B2(new_n895), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n899), .A3(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n719), .A2(new_n737), .A3(new_n836), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G148gat), .ZN(new_n907));
  XNOR2_X1  g706(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT122), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n301), .B1(new_n904), .B2(new_n905), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(new_n908), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n891), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n883), .A2(new_n301), .A3(new_n663), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n880), .B2(new_n601), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n883), .A2(new_n298), .A3(new_n685), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  AOI21_X1  g718(.A(G162gat), .B1(new_n883), .B2(new_n634), .ZN(new_n920));
  INV_X1    g719(.A(new_n880), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n636), .A2(new_n299), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(G1347gat));
  NOR2_X1   g722(.A1(new_n477), .A2(new_n417), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n833), .A2(new_n834), .A3(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n925), .A2(new_n245), .A3(new_n561), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n477), .B1(new_n826), .B2(new_n827), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(new_n428), .A3(new_n295), .A4(new_n434), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n560), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n926), .B1(new_n930), .B2(new_n245), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n925), .B2(new_n737), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n663), .A2(new_n246), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n928), .B2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n262), .A3(new_n685), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n925), .B2(new_n601), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n929), .A2(new_n225), .A3(new_n634), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  INV_X1    g739(.A(new_n925), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n634), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(G190gat), .ZN(new_n943));
  AOI211_X1 g742(.A(KEYINPUT61), .B(new_n225), .C1(new_n941), .C2(new_n634), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n939), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT123), .ZN(G1351gat));
  NAND3_X1  g745(.A1(new_n473), .A2(new_n428), .A3(new_n724), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n927), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(G197gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n560), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n473), .A2(new_n924), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT126), .Z(new_n957));
  AND2_X1   g756(.A1(new_n904), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(new_n560), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n955), .B1(new_n959), .B2(new_n953), .ZN(G1352gat));
  NOR3_X1   g759(.A1(new_n951), .A2(G204gat), .A3(new_n737), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT62), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n958), .A2(new_n663), .ZN(new_n963));
  INV_X1    g762(.A(G204gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(G1353gat));
  NAND3_X1  g764(.A1(new_n952), .A2(new_n318), .A3(new_n685), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n958), .A2(new_n685), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n967), .B2(G211gat), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT63), .ZN(new_n969));
  AOI211_X1 g768(.A(new_n969), .B(new_n318), .C1(new_n958), .C2(new_n685), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(G1354gat));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n958), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n634), .B1(new_n958), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g773(.A(G218gat), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n952), .A2(new_n319), .A3(new_n634), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


