//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(G355));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n203), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n215), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n215), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n213), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(new_n207), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n224), .B(new_n227), .C1(new_n229), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(G97), .B(G107), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G68), .Z(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n228), .ZN(new_n248));
  AOI21_X1  g0048(.A(new_n248), .B1(new_n212), .B2(G20), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G77), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n250), .B1(G77), .B2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n248), .ZN(new_n253));
  XOR2_X1   g0053(.A(KEYINPUT8), .B(G58), .Z(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n254), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT15), .B(G87), .Z(new_n257));
  NAND2_X1  g0057(.A1(new_n213), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n253), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n252), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT66), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G41), .ZN(new_n266));
  AOI21_X1  g0066(.A(G45), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n212), .A2(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G1), .A3(G13), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n212), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(new_n274), .A2(G244), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G232), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G107), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(G1698), .ZN(new_n280));
  OAI221_X1 g0080(.A(new_n278), .B1(new_n279), .B2(new_n276), .C1(new_n280), .C2(new_n218), .ZN(new_n281));
  INV_X1    g0081(.A(new_n271), .ZN(new_n282));
  AOI211_X1 g0082(.A(new_n269), .B(new_n275), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G200), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n262), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n283), .A2(G190), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n285), .A2(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n208), .A2(G20), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n254), .A2(new_n259), .B1(G150), .B2(new_n255), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n253), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n249), .A2(G50), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n295), .B1(G50), .B2(new_n251), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n276), .A2(G222), .A3(new_n277), .ZN(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  INV_X1    g0100(.A(G223), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n299), .B1(new_n300), .B2(new_n276), .C1(new_n280), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n282), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n269), .B1(G226), .B2(new_n274), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n298), .B1(new_n306), .B2(G169), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(G179), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(KEYINPUT67), .ZN(new_n311));
  OR2_X1    g0111(.A1(new_n283), .A2(G169), .ZN(new_n312));
  INV_X1    g0112(.A(new_n262), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n283), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  AND4_X1   g0116(.A1(new_n291), .A2(new_n310), .A3(new_n311), .A4(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT70), .B1(new_n305), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(G200), .B2(new_n305), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT69), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT9), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(KEYINPUT69), .A2(KEYINPUT9), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n298), .B2(new_n324), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n298), .A2(new_n324), .A3(new_n323), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n320), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT10), .ZN(new_n328));
  INV_X1    g0128(.A(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT3), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT7), .B1(new_n333), .B2(new_n213), .ZN(new_n336));
  OAI21_X1  g0136(.A(G68), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(KEYINPUT16), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT16), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n276), .B2(G20), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n203), .B1(new_n343), .B2(new_n334), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n202), .A2(new_n203), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n206), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n255), .A2(G159), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n341), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n340), .A2(new_n349), .A3(new_n248), .ZN(new_n350));
  INV_X1    g0150(.A(new_n254), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n251), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n249), .B2(new_n351), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n273), .A2(new_n217), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT77), .B1(new_n269), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n276), .A2(G226), .A3(G1698), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n330), .A2(new_n332), .A3(G223), .A4(new_n277), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G33), .A2(G87), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n282), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n362), .B1(new_n273), .B2(new_n217), .C1(new_n267), .C2(new_n268), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n356), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n269), .A2(new_n355), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n364), .A2(new_n314), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n354), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT18), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n284), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n356), .A2(new_n361), .A3(new_n363), .A4(new_n318), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(new_n350), .A3(new_n353), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT17), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n317), .A2(new_n328), .A3(new_n371), .A4(new_n376), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n258), .A2(new_n300), .B1(new_n213), .B2(G68), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(KEYINPUT74), .B1(G50), .B2(new_n255), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(KEYINPUT74), .B2(new_n378), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n248), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT11), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT75), .B1(new_n251), .B2(G68), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT12), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(G68), .B2(new_n249), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT76), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT13), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n330), .A2(new_n332), .A3(G232), .A4(G1698), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT71), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n276), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G97), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n276), .A2(G226), .A3(new_n277), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n282), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n267), .A2(new_n268), .B1(new_n273), .B2(new_n218), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n388), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AOI211_X1 g0199(.A(KEYINPUT13), .B(new_n397), .C1(new_n395), .C2(new_n282), .ZN(new_n400));
  OAI21_X1  g0200(.A(G169), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(G169), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n396), .A2(new_n388), .A3(new_n398), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT73), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n396), .A2(new_n398), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n388), .B1(new_n409), .B2(KEYINPUT72), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n397), .B1(new_n395), .B2(new_n282), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT72), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n408), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT13), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  AOI211_X1 g0215(.A(KEYINPUT72), .B(new_n397), .C1(new_n395), .C2(new_n282), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n415), .A2(new_n407), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(G179), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n387), .B1(new_n405), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n407), .B(new_n406), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n409), .A2(KEYINPUT72), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n421), .A2(KEYINPUT73), .A3(KEYINPUT13), .A4(new_n413), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n314), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n402), .A2(new_n404), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT76), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n386), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  OR2_X1    g0226(.A1(new_n399), .A2(new_n400), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n386), .B1(G200), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(G190), .B1(new_n414), .B2(new_n417), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT88), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n331), .A2(G33), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n329), .A2(KEYINPUT3), .ZN(new_n434));
  OAI21_X1  g0234(.A(G303), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n330), .A2(new_n332), .A3(G257), .A4(new_n277), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n330), .A2(new_n332), .A3(G264), .A4(G1698), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n282), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT5), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n264), .A2(new_n266), .A3(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n212), .B(G45), .C1(new_n441), .C2(G41), .ZN(new_n443));
  OAI211_X1 g0243(.A(G270), .B(new_n271), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT66), .B(G41), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n445), .B2(new_n441), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G274), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n432), .B1(new_n440), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n443), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n264), .A2(new_n266), .A3(new_n441), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n282), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(G270), .B1(new_n446), .B2(G274), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(KEYINPUT88), .A3(new_n439), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n365), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n213), .C1(G33), .C2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n248), .C1(new_n213), .C2(G116), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT20), .ZN(new_n460));
  INV_X1    g0260(.A(new_n251), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n329), .A2(KEYINPUT79), .A3(G1), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT79), .B1(new_n329), .B2(G1), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n253), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n463), .B1(new_n467), .B2(new_n462), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n460), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT21), .B1(new_n455), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT89), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n440), .A2(new_n448), .A3(new_n314), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n455), .B2(KEYINPUT21), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(new_n469), .ZN(new_n475));
  AND4_X1   g0275(.A1(KEYINPUT88), .A2(new_n439), .A3(new_n447), .A4(new_n444), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT88), .B1(new_n453), .B2(new_n439), .ZN(new_n477));
  OAI211_X1 g0277(.A(KEYINPUT21), .B(G169), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n473), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT89), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n471), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT78), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT6), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n241), .A2(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n484), .A2(new_n457), .A3(G107), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n213), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n255), .A2(G77), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n483), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n486), .B1(new_n484), .B2(new_n241), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT78), .B(new_n489), .C1(new_n492), .C2(new_n213), .ZN(new_n493));
  OAI21_X1  g0293(.A(G107), .B1(new_n335), .B2(new_n336), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n248), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n251), .A2(G97), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(G97), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n452), .A2(G257), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n500), .A2(new_n447), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n330), .A2(new_n332), .A3(G244), .A4(new_n277), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n276), .A2(KEYINPUT4), .A3(G244), .A4(new_n277), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n276), .A2(G250), .A3(G1698), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n504), .A2(new_n505), .A3(new_n456), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n282), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(G190), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n496), .A2(new_n499), .A3(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n507), .A2(KEYINPUT80), .A3(new_n282), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT80), .B1(new_n507), .B2(new_n282), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n501), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n284), .B1(new_n513), .B2(KEYINPUT81), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT81), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n515), .B(new_n501), .C1(new_n511), .C2(new_n512), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(G87), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT90), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(KEYINPUT22), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n276), .A2(new_n213), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n519), .B2(KEYINPUT22), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n276), .A2(new_n520), .A3(new_n213), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT91), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(G20), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n213), .A2(KEYINPUT91), .A3(G33), .A4(G116), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n213), .B2(G107), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n279), .A2(KEYINPUT23), .A3(G20), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n525), .A2(KEYINPUT24), .A3(new_n533), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n248), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n330), .A2(new_n332), .A3(G250), .A4(new_n277), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n330), .A2(new_n332), .A3(G257), .A4(G1698), .ZN(new_n540));
  INV_X1    g0340(.A(G294), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n540), .C1(new_n329), .C2(new_n541), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n282), .B1(new_n452), .B2(G264), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n543), .A2(G190), .A3(new_n447), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n251), .A2(G107), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT25), .ZN(new_n546));
  OR2_X1    g0346(.A1(new_n546), .A2(KEYINPUT92), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(KEYINPUT92), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n547), .B(new_n548), .C1(KEYINPUT25), .C2(new_n545), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n498), .A2(G107), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(new_n282), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n452), .A2(G264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n447), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(G200), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n538), .A2(new_n544), .A3(new_n551), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n496), .A2(new_n499), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n314), .B(new_n501), .C1(new_n511), .C2(new_n512), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n501), .A2(new_n508), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n365), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n517), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n554), .A2(new_n365), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n543), .A2(new_n314), .A3(new_n447), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n538), .B2(new_n551), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(G200), .B1(new_n476), .B2(new_n477), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n449), .A2(G190), .A3(new_n454), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n469), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n257), .A2(new_n251), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n276), .A2(KEYINPUT86), .A3(new_n213), .A4(G68), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n330), .A2(new_n332), .A3(new_n213), .A4(G68), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT86), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n213), .A2(G33), .A3(G97), .ZN(new_n577));
  NAND2_X1  g0377(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT87), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT87), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n577), .B(new_n583), .C1(new_n579), .C2(new_n580), .ZN(new_n584));
  AND4_X1   g0384(.A1(new_n573), .A2(new_n576), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  OR2_X1    g0385(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n586));
  AND2_X1   g0386(.A1(G33), .A2(G97), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n578), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n213), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT85), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n213), .ZN(new_n592));
  NOR3_X1   g0392(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n572), .B1(new_n596), .B2(new_n248), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n330), .A2(new_n332), .A3(G244), .A4(G1698), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT83), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n276), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n276), .A2(G238), .A3(new_n277), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n527), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n282), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n212), .A2(G45), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n605), .B(KEYINPUT82), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n271), .A2(G250), .ZN(new_n607));
  INV_X1    g0407(.A(G45), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n606), .A2(new_n607), .B1(new_n608), .B2(new_n268), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G200), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n609), .B1(new_n282), .B2(new_n603), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G190), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n498), .A2(G87), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n597), .A2(new_n612), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n588), .A2(KEYINPUT85), .A3(new_n213), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT85), .B1(new_n588), .B2(new_n213), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n617), .A2(new_n618), .A3(new_n593), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n576), .A2(new_n582), .A3(new_n573), .A4(new_n584), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n248), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n572), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n498), .A2(new_n257), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n611), .A2(new_n365), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n613), .A2(new_n314), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n571), .A2(new_n616), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n482), .A2(new_n563), .A3(new_n568), .A4(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n377), .A2(new_n431), .A3(new_n629), .ZN(G372));
  NAND2_X1  g0430(.A1(new_n310), .A2(new_n311), .ZN(new_n631));
  INV_X1    g0431(.A(new_n386), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n405), .A2(new_n418), .A3(new_n387), .ZN(new_n633));
  OAI21_X1  g0433(.A(KEYINPUT76), .B1(new_n423), .B2(new_n424), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n316), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n430), .A2(new_n376), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n371), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n631), .B1(new_n639), .B2(new_n328), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n377), .A2(new_n431), .ZN(new_n641));
  INV_X1    g0441(.A(new_n510), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n500), .A2(new_n447), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT80), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n508), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n507), .A2(KEYINPUT80), .A3(new_n282), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(G200), .B1(new_n647), .B2(new_n515), .ZN(new_n648));
  INV_X1    g0448(.A(new_n516), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n496), .A2(new_n499), .B1(new_n560), .B2(new_n365), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n559), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n556), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n480), .A2(new_n471), .A3(new_n567), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT93), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n621), .A2(new_n622), .A3(new_n615), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n613), .A2(new_n284), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n597), .A2(new_n612), .A3(KEYINPUT93), .A4(new_n615), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n614), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n627), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n653), .A2(new_n654), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n660), .A2(new_n663), .A3(new_n562), .A4(new_n627), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n651), .A2(new_n627), .A3(new_n616), .A4(new_n559), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n627), .A3(new_n666), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n641), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n640), .A2(new_n669), .ZN(G369));
  INV_X1    g0470(.A(G13), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(new_n212), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n538), .B2(new_n551), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n568), .B1(new_n557), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n567), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT95), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n482), .A2(new_n678), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n684), .A2(new_n685), .B1(new_n567), .B2(new_n679), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n469), .A2(new_n679), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT94), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n482), .A2(new_n571), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n480), .A2(new_n471), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n684), .A2(new_n691), .A3(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n686), .A2(new_n692), .ZN(G399));
  INV_X1    g0493(.A(new_n225), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(new_n445), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n594), .A2(G116), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(G1), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n230), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n696), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n668), .A2(new_n679), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n471), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n480), .A2(KEYINPUT89), .ZN(new_n706));
  AOI211_X1 g0506(.A(new_n472), .B(new_n469), .C1(new_n478), .C2(new_n479), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n705), .B(new_n568), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n661), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n563), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT26), .B1(new_n661), .B2(new_n652), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(new_n627), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT29), .B(new_n679), .C1(new_n711), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n704), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n501), .A2(new_n543), .A3(new_n508), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n473), .A3(KEYINPUT30), .A4(new_n613), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n613), .A2(G179), .A3(new_n439), .A4(new_n453), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n501), .A2(new_n543), .A3(new_n508), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT96), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n449), .A2(new_n454), .ZN(new_n725));
  AOI21_X1  g0525(.A(G179), .B1(new_n543), .B2(new_n447), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n611), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n724), .B1(new_n727), .B2(new_n647), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n726), .A2(new_n611), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n725), .A3(KEYINPUT96), .A4(new_n513), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n723), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT97), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n678), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI211_X1 g0533(.A(KEYINPUT97), .B(new_n723), .C1(new_n728), .C2(new_n730), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n628), .A2(new_n556), .A3(new_n650), .A4(new_n652), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n708), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n679), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n735), .B1(new_n738), .B2(KEYINPUT31), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  INV_X1    g0540(.A(new_n723), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n729), .A2(new_n725), .A3(new_n513), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n740), .B(new_n679), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(G330), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n716), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n701), .B1(new_n746), .B2(G1), .ZN(G364));
  AOI21_X1  g0547(.A(new_n212), .B1(new_n672), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n695), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n691), .B2(G330), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n691), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n228), .B1(G20), .B2(new_n365), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n213), .A2(new_n318), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n284), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n314), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G322), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n333), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n213), .A2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G179), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n760), .B(new_n764), .C1(G329), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n213), .B1(new_n766), .B2(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G294), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT98), .ZN(new_n773));
  AND3_X1   g0573(.A1(new_n761), .A2(new_n765), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n773), .B1(new_n761), .B2(new_n765), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G311), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n314), .A2(new_n284), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n765), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  NAND2_X1  g0581(.A1(new_n756), .A2(new_n779), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n765), .A2(new_n757), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n784), .B1(G283), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n769), .A2(new_n772), .A3(new_n778), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n777), .A2(G77), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n767), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT32), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n276), .B1(new_n762), .B2(new_n202), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(G97), .B2(new_n771), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n782), .A2(new_n207), .B1(new_n758), .B2(new_n518), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n780), .A2(new_n203), .B1(new_n785), .B2(new_n279), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n789), .A2(new_n792), .A3(new_n794), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n755), .B1(new_n788), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n754), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n694), .A2(new_n333), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n804), .A2(G355), .B1(new_n462), .B2(new_n694), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n694), .A2(new_n276), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n699), .B2(G45), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n245), .A2(new_n608), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n753), .B(new_n799), .C1(new_n803), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n802), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n691), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n752), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  NOR2_X1   g0614(.A1(new_n754), .A2(new_n800), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n753), .B1(new_n300), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n762), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G294), .A2(new_n817), .B1(new_n768), .B2(G311), .ZN(new_n818));
  INV_X1    g0618(.A(G283), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n780), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n786), .A2(G87), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n279), .B2(new_n758), .ZN(new_n822));
  INV_X1    g0622(.A(new_n782), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n276), .B(new_n822), .C1(G303), .C2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n457), .B2(new_n770), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n820), .B(new_n825), .C1(G116), .C2(new_n777), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G137), .A2(new_n823), .B1(new_n817), .B2(G143), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n828), .B2(new_n780), .C1(new_n790), .C2(new_n776), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n276), .B1(new_n758), .B2(new_n207), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n785), .A2(new_n203), .B1(new_n767), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(G58), .C2(new_n771), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n826), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n316), .A2(KEYINPUT99), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n316), .A2(KEYINPUT99), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(new_n837), .B1(new_n289), .B2(new_n290), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n313), .A2(new_n678), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n636), .A2(new_n678), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n816), .B1(new_n755), .B2(new_n835), .C1(new_n842), .C2(new_n801), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n668), .B2(new_n679), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n679), .B(new_n838), .C1(new_n662), .C2(new_n667), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(G330), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT31), .B1(new_n629), .B2(new_n678), .ZN(new_n849));
  INV_X1    g0649(.A(new_n735), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n743), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n753), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n744), .A2(new_n844), .A3(new_n846), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n843), .B1(new_n854), .B2(new_n855), .ZN(G384));
  INV_X1    g0656(.A(new_n492), .ZN(new_n857));
  OAI211_X1 g0657(.A(G116), .B(new_n229), .C1(new_n857), .C2(KEYINPUT35), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(KEYINPUT35), .B2(new_n857), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT36), .Z(new_n860));
  NOR3_X1   g0660(.A1(new_n699), .A2(new_n300), .A3(new_n345), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n861), .A2(KEYINPUT100), .B1(G50), .B2(new_n203), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(KEYINPUT100), .B2(new_n861), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n671), .A2(G1), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n836), .A2(new_n679), .A3(new_n837), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n845), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT101), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n845), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n430), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n386), .A2(new_n678), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n635), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n632), .B(new_n679), .C1(new_n633), .C2(new_n634), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n349), .A2(new_n248), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT102), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n349), .A2(new_n880), .A3(new_n248), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n879), .A2(new_n340), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n353), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT103), .ZN(new_n884));
  INV_X1    g0684(.A(new_n676), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n353), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n344), .A2(new_n348), .A3(new_n341), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n878), .B2(KEYINPUT102), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n889), .B2(new_n881), .ZN(new_n890));
  OAI21_X1  g0690(.A(KEYINPUT103), .B1(new_n890), .B2(new_n676), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n371), .A2(new_n376), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n375), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n883), .B2(new_n368), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n886), .A3(new_n891), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n354), .B1(new_n368), .B2(new_n885), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n899), .A2(KEYINPUT37), .A3(new_n894), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT38), .B(new_n893), .C1(new_n897), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n900), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n902), .B1(new_n903), .B2(new_n892), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n870), .A2(new_n877), .A3(new_n905), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n371), .A2(new_n885), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n375), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n374), .A2(KEYINPUT104), .A3(new_n350), .A4(new_n353), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n898), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT105), .ZN(new_n913));
  INV_X1    g0713(.A(new_n900), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT105), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n915), .A3(KEYINPUT37), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n371), .A2(new_n376), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n354), .A3(new_n885), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n901), .B(new_n904), .C1(new_n920), .C2(KEYINPUT106), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n903), .A2(new_n902), .A3(new_n892), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(new_n920), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT106), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n924), .A2(KEYINPUT39), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n921), .A2(KEYINPUT39), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n635), .A2(new_n679), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n906), .B(new_n907), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n704), .A2(new_n715), .A3(new_n641), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n640), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n928), .B(new_n930), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n735), .A2(KEYINPUT31), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n740), .B1(new_n737), .B2(new_n679), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n933), .B2(new_n735), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G330), .A3(new_n641), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n838), .A2(new_n839), .B1(new_n636), .B2(new_n678), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n426), .A2(new_n430), .A3(new_n872), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n635), .A2(new_n678), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n934), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n905), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n733), .A2(new_n734), .A3(new_n740), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n849), .B2(new_n850), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n842), .B1(new_n874), .B2(new_n875), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT107), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n923), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n947), .A2(new_n941), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n943), .B1(new_n949), .B2(KEYINPUT40), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n935), .B1(new_n950), .B2(new_n848), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n934), .A2(new_n939), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n923), .B1(new_n953), .B2(KEYINPUT107), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n952), .B1(new_n954), .B2(new_n941), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n641), .B(new_n934), .C1(new_n955), .C2(new_n943), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n931), .A2(new_n951), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n212), .B2(new_n672), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n931), .B1(new_n951), .B2(new_n956), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n860), .B1(new_n863), .B2(new_n864), .C1(new_n958), .C2(new_n959), .ZN(G367));
  NAND2_X1  g0760(.A1(new_n656), .A2(new_n678), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n709), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n627), .B2(new_n961), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT108), .Z(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n684), .A2(new_n685), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n652), .A2(new_n679), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n558), .A2(new_n678), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n650), .A2(new_n652), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n969), .A2(KEYINPUT42), .A3(new_n568), .A4(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT42), .ZN(new_n976));
  INV_X1    g0776(.A(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n976), .B1(new_n686), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n652), .A2(new_n678), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n966), .B(new_n967), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n975), .A2(new_n978), .B1(new_n562), .B2(new_n679), .ZN(new_n982));
  INV_X1    g0782(.A(new_n967), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n965), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n692), .A2(new_n977), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n981), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n985), .B1(new_n981), .B2(new_n984), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n695), .B(KEYINPUT41), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n692), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n968), .A2(new_n682), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n992), .A2(KEYINPUT111), .A3(new_n977), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT111), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n686), .B2(new_n974), .ZN(new_n995));
  XOR2_X1   g0795(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n996));
  NAND3_X1  g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT45), .B1(new_n992), .B2(new_n977), .ZN(new_n999));
  INV_X1    g0799(.A(new_n996), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n994), .B(new_n1000), .C1(new_n686), .C2(new_n974), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT45), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n686), .A2(new_n1002), .A3(new_n974), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n991), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n999), .A2(new_n1003), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1006), .A2(new_n692), .A3(new_n997), .A4(new_n1001), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n684), .B(new_n685), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n691), .A2(G330), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1010), .A2(new_n745), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1005), .A2(new_n1007), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n990), .B1(new_n1012), .B2(new_n746), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n988), .B1(new_n1013), .B2(new_n749), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n806), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n238), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n257), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n803), .B1(new_n225), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n750), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(G143), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n276), .B1(new_n782), .B2(new_n1020), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n762), .A2(new_n828), .B1(new_n785), .B2(new_n300), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G68), .C2(new_n771), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n202), .A2(new_n758), .B1(new_n780), .B2(new_n790), .ZN(new_n1024));
  XOR2_X1   g0824(.A(KEYINPUT113), .B(G137), .Z(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(new_n768), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1023), .B(new_n1026), .C1(new_n207), .C2(new_n776), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n758), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(G116), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT46), .ZN(new_n1030));
  INV_X1    g0830(.A(G311), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n782), .A2(new_n1031), .B1(new_n780), .B2(new_n541), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n762), .A2(new_n759), .B1(new_n785), .B2(new_n457), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n770), .A2(new_n279), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(KEYINPUT112), .B(G317), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n276), .B(new_n1035), .C1(new_n768), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n777), .A2(G283), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1030), .A2(new_n1034), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT47), .B1(new_n1027), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1040), .A2(new_n755), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1027), .A2(KEYINPUT47), .A3(new_n1039), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1019), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n963), .B2(new_n811), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1014), .A2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT114), .Z(G387));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n254), .A2(new_n207), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n697), .B(new_n1047), .C1(new_n1048), .C2(KEYINPUT50), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(KEYINPUT50), .B2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n806), .B1(new_n235), .B2(new_n608), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n804), .B1(G116), .B2(new_n594), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n225), .A2(G107), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n803), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n750), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n762), .A2(new_n207), .B1(new_n767), .B2(new_n828), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n333), .B(new_n1057), .C1(G97), .C2(new_n786), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1017), .A2(new_n770), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n777), .A2(G68), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n351), .A2(new_n780), .B1(new_n300), .B2(new_n758), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G159), .B2(new_n823), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n276), .B1(new_n768), .B2(G326), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n780), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n817), .A2(new_n1036), .B1(new_n1066), .B2(G311), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n763), .B2(new_n782), .C1(new_n776), .C2(new_n759), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT48), .Z(new_n1069));
  OAI22_X1  g0869(.A1(new_n758), .A2(new_n541), .B1(new_n770), .B2(new_n819), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1065), .B1(new_n462), .B2(new_n785), .C1(new_n1071), .C2(KEYINPUT49), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1064), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1056), .B1(new_n1074), .B2(new_n754), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n684), .B2(new_n811), .ZN(new_n1076));
  AND2_X1   g0876(.A1(new_n1010), .A2(new_n745), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n695), .B1(new_n1010), .B2(new_n745), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1076), .B1(new_n748), .B2(new_n1010), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  NAND3_X1  g0879(.A1(new_n1005), .A2(new_n1007), .A3(new_n749), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1015), .A2(new_n242), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n803), .B1(new_n457), .B2(new_n225), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n750), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n758), .A2(new_n819), .B1(new_n767), .B2(new_n763), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n333), .B1(new_n770), .B2(new_n462), .C1(new_n279), .C2(new_n785), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(G303), .C2(new_n1066), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT52), .ZN(new_n1087));
  INV_X1    g0887(.A(G317), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n782), .A2(new_n1088), .B1(new_n762), .B2(new_n1031), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n777), .A2(G294), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1086), .B(new_n1090), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n776), .A2(new_n351), .B1(new_n207), .B2(new_n780), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT115), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n782), .A2(new_n828), .B1(new_n762), .B2(new_n790), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT51), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n771), .A2(G77), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n333), .B1(new_n786), .B2(G87), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G68), .A2(new_n1028), .B1(new_n768), .B2(G143), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1091), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1083), .B1(new_n1100), .B2(new_n754), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n974), .B2(new_n811), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1012), .A2(new_n695), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1011), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1080), .B(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(G390));
  OAI211_X1 g0905(.A(new_n679), .B(new_n838), .C1(new_n711), .C2(new_n714), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1106), .A2(new_n865), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n948), .B(new_n927), .C1(new_n1107), .C2(new_n876), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n853), .A2(new_n939), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n927), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n870), .B2(new_n877), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n917), .A2(new_n919), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT106), .B1(new_n1112), .B2(new_n902), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT39), .B1(new_n905), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n923), .A2(new_n925), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1108), .B(new_n1109), .C1(new_n1111), .C2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n848), .B1(new_n851), .B2(new_n932), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1119), .A2(new_n946), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n927), .B1(new_n922), .B2(new_n920), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1106), .A2(new_n865), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n877), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n845), .A2(new_n868), .A3(new_n865), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n868), .B1(new_n845), .B2(new_n865), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n877), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n927), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1124), .B1(new_n1128), .B2(new_n926), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1117), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n842), .C1(new_n739), .C2(new_n743), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1131), .A2(new_n876), .B1(new_n1118), .B2(new_n939), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n870), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1107), .B1(new_n744), .B2(new_n946), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n877), .B1(new_n1118), .B2(new_n842), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1132), .A2(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n935), .A2(KEYINPUT116), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT116), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n934), .A2(new_n641), .A3(new_n1138), .A4(G330), .ZN(new_n1139));
  AND4_X1   g0939(.A1(new_n640), .A2(new_n1137), .A3(new_n929), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n1130), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1130), .A2(new_n1141), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n695), .A3(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1117), .B(new_n749), .C1(new_n1121), .C2(new_n1129), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n753), .B1(new_n351), .B2(new_n815), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT117), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n276), .B1(new_n1028), .B2(G87), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G68), .A2(new_n786), .B1(new_n768), .B2(G294), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n279), .B2(new_n780), .C1(new_n819), .C2(new_n782), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(G97), .C2(new_n777), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1096), .B1(new_n462), .B2(new_n762), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT119), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n276), .B1(new_n770), .B2(new_n790), .C1(new_n207), .C2(new_n785), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1025), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1157), .A2(new_n780), .B1(new_n1158), .B2(new_n767), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n782), .A2(new_n1160), .B1(new_n762), .B2(new_n832), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1156), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT54), .B(G143), .Z(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1028), .A3(G150), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1164), .B1(new_n758), .B2(new_n828), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n777), .A2(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1152), .A2(new_n1155), .B1(new_n1162), .B2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1147), .B1(new_n755), .B2(new_n1169), .C1(new_n1116), .C2(new_n801), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1145), .A2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(KEYINPUT120), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(KEYINPUT120), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1144), .B1(new_n1172), .B2(new_n1173), .ZN(G378));
  OAI22_X1  g0974(.A1(new_n782), .A2(new_n462), .B1(new_n785), .B2(new_n202), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G107), .A2(new_n817), .B1(new_n768), .B2(G283), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n457), .B2(new_n780), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1175), .B(new_n1177), .C1(G68), .C2(new_n771), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n276), .A2(new_n445), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n300), .B2(new_n758), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT121), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n777), .A2(new_n257), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1178), .B(new_n1182), .C1(new_n1181), .C2(new_n1180), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT58), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1185), .B(new_n1186), .C1(new_n1179), .C2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G132), .A2(new_n1066), .B1(new_n1028), .B2(new_n1163), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1160), .B2(new_n762), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G137), .B2(new_n777), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n782), .A2(new_n1158), .B1(new_n770), .B2(new_n828), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT122), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n768), .C2(G124), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n790), .B2(new_n785), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n754), .B1(new_n1188), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n753), .B1(new_n207), .B2(new_n815), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n328), .B1(new_n308), .B2(new_n307), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT56), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n297), .A2(new_n676), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT55), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT123), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1203), .B(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1200), .B(new_n1201), .C1(new_n1207), .C2(new_n801), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n950), .B2(new_n848), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1207), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G330), .B(new_n1211), .C1(new_n955), .C2(new_n943), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n928), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1209), .B1(new_n1216), .B2(new_n749), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1140), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT57), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1210), .A2(new_n1212), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n928), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(KEYINPUT57), .A3(new_n1222), .A4(new_n1218), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n695), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1219), .B2(new_n1224), .ZN(G375));
  AOI21_X1  g1025(.A(new_n753), .B1(new_n203), .B2(new_n815), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n817), .A2(new_n1025), .B1(new_n1066), .B2(new_n1163), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n832), .B2(new_n782), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G150), .B2(new_n777), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n276), .B1(new_n785), .B2(new_n202), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n758), .A2(new_n790), .B1(new_n767), .B2(new_n1160), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(G50), .C2(new_n771), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(G97), .A2(new_n1028), .B1(new_n768), .B2(G303), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n541), .B2(new_n782), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G107), .B2(new_n777), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n762), .A2(new_n819), .B1(new_n780), .B2(new_n462), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n333), .B1(new_n785), .B2(new_n300), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1059), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1229), .A2(new_n1232), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1226), .B1(new_n755), .B2(new_n1239), .C1(new_n877), .C2(new_n801), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1136), .B2(new_n749), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1141), .A2(new_n989), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(G381));
  INV_X1    g1045(.A(G375), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1171), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1144), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  OR4_X1    g1050(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1251));
  OR4_X1    g1051(.A1(G387), .A2(new_n1250), .A3(G381), .A4(new_n1251), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1250), .ZN(G409));
  INV_X1    g1053(.A(KEYINPUT62), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n677), .A2(G213), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n696), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1244), .B2(KEYINPUT60), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT124), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1244), .A2(new_n1260), .A3(KEYINPUT60), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1137), .A2(new_n929), .A3(new_n640), .A4(new_n1139), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .A4(KEYINPUT60), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT124), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1259), .B1(new_n1261), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1242), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1257), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1266), .A2(new_n1261), .ZN(new_n1270));
  OAI211_X1 g1070(.A(G384), .B(new_n1242), .C1(new_n1270), .C2(new_n1259), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  OAI211_X1 g1072(.A(G378), .B(new_n1217), .C1(new_n1219), .C2(new_n1224), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1221), .A2(new_n989), .A3(new_n1222), .A4(new_n1218), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1221), .A2(new_n749), .A3(new_n1222), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1208), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1249), .A2(new_n1276), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1256), .B(new_n1272), .C1(new_n1273), .C2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1254), .B1(new_n1278), .B2(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1272), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1255), .A3(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT127), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(new_n1283), .A3(KEYINPUT62), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1255), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1256), .A2(G2897), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1272), .B(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT61), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1279), .A2(new_n1284), .A3(new_n1288), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(G393), .B(new_n813), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1014), .A2(new_n1044), .A3(G390), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G390), .B1(new_n1014), .B2(new_n1044), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(G390), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1045), .A2(KEYINPUT125), .A3(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1290), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT126), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT126), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1298), .B(new_n1290), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1294), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1290), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1301), .A2(new_n1291), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1297), .A2(new_n1299), .B1(new_n1300), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1289), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1278), .A2(KEYINPUT63), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1278), .A2(KEYINPUT63), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1288), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1304), .A2(new_n1310), .ZN(G405));
  OAI21_X1  g1111(.A(new_n1273), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1281), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1273), .B(new_n1272), .C1(new_n1246), .C2(new_n1248), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(new_n1303), .B(new_n1315), .ZN(G402));
endmodule


