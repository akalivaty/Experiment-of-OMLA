//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT71), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n203), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  NAND4_X1  g009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G127gat), .B(G134gat), .Z(new_n212));
  XNOR2_X1  g011(.A(G113gat), .B(G120gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(KEYINPUT1), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT27), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G183gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT27), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n217), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(KEYINPUT27), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(G183gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT69), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G190gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n226), .ZN(new_n231));
  AND3_X1   g030(.A1(new_n228), .A2(KEYINPUT70), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT70), .B1(new_n228), .B2(new_n231), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT26), .ZN(new_n237));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n236), .A2(KEYINPUT26), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n232), .A2(new_n233), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G169gat), .ZN(new_n244));
  INV_X1    g043(.A(G176gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT23), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n236), .B2(KEYINPUT23), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n250), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n220), .A2(new_n229), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT24), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT68), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n246), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n249), .B2(new_n251), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(new_n254), .A3(new_n255), .A4(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n265), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n255), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT65), .B1(new_n272), .B2(new_n256), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n259), .A2(new_n254), .A3(new_n274), .A4(new_n255), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n235), .B1(KEYINPUT23), .B2(new_n236), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n273), .A2(new_n275), .A3(new_n252), .A4(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n263), .A2(new_n270), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n216), .B1(new_n243), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT64), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n271), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n253), .A2(new_n262), .A3(KEYINPUT68), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n266), .B1(new_n265), .B2(new_n269), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n228), .A2(new_n231), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n228), .A2(new_n231), .A3(KEYINPUT70), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n241), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n290), .A3(new_n215), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n279), .A2(new_n281), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT33), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G71gat), .B(G99gat), .Z(new_n296));
  XNOR2_X1  g095(.A(G15gat), .B(G43gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n293), .B1(new_n298), .B2(KEYINPUT33), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n292), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT72), .B1(new_n292), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT34), .ZN(new_n304));
  INV_X1    g103(.A(new_n281), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(KEYINPUT73), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n279), .A2(new_n291), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n307), .B1(new_n308), .B2(new_n305), .ZN(new_n309));
  AOI211_X1 g108(.A(new_n281), .B(new_n306), .C1(new_n279), .C2(new_n291), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n303), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n292), .A2(new_n300), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n292), .A2(KEYINPUT72), .A3(new_n300), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n311), .B1(new_n318), .B2(new_n299), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n202), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n312), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n311), .A3(new_n299), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT36), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G8gat), .B(G36gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n325), .B(new_n326), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(G197gat), .A2(G204gat), .ZN(new_n329));
  AND2_X1   g128(.A1(G197gat), .A2(G204gat), .ZN(new_n330));
  AND2_X1   g129(.A1(G211gat), .A2(G218gat), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n329), .A2(new_n330), .B1(new_n331), .B2(KEYINPUT22), .ZN(new_n332));
  XOR2_X1   g131(.A(G211gat), .B(G218gat), .Z(new_n333));
  OR2_X1    g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n333), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n243), .B2(new_n278), .ZN(new_n340));
  NAND2_X1  g139(.A1(G226gat), .A2(G233gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n243), .B2(new_n278), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n338), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n285), .B2(new_n290), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n344), .B(new_n338), .C1(new_n346), .C2(new_n343), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n328), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n344), .B1(new_n346), .B2(new_n343), .ZN(new_n350));
  INV_X1    g149(.A(new_n338), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n347), .A3(new_n327), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(KEYINPUT30), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n352), .A2(new_n355), .A3(new_n347), .A4(new_n327), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G1gat), .B(G29gat), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT0), .ZN(new_n359));
  XOR2_X1   g158(.A(G57gat), .B(G85gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT5), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G162gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G155gat), .ZN(new_n367));
  INV_X1    g166(.A(G155gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G162gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G141gat), .B(G148gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(KEYINPUT2), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(G141gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT75), .B(G148gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(G141gat), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT2), .B1(new_n366), .B2(KEYINPUT76), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(new_n367), .A3(new_n369), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(KEYINPUT75), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT75), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G148gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n383), .A3(G141gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G141gat), .B2(new_n373), .ZN(new_n385));
  INV_X1    g184(.A(new_n378), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n372), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n380), .A2(new_n389), .A3(new_n215), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n211), .A2(new_n214), .A3(new_n372), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n378), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT4), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n393), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT77), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT77), .B(KEYINPUT4), .C1(new_n392), .C2(new_n393), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n365), .B(new_n391), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n214), .A2(new_n372), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n387), .A4(new_n211), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n394), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n390), .A3(new_n362), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  INV_X1    g204(.A(new_n379), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n406), .A2(new_n216), .B1(new_n392), .B2(new_n393), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(new_n363), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(KEYINPUT6), .B(new_n361), .C1(new_n399), .C2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n361), .B1(new_n399), .B2(new_n409), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n364), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n361), .B1(new_n404), .B2(new_n408), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT6), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n415), .B2(KEYINPUT78), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  AOI211_X1 g216(.A(new_n417), .B(KEYINPUT6), .C1(new_n413), .C2(new_n414), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n410), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n357), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n334), .B(KEYINPUT74), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n337), .B(KEYINPUT79), .Z(new_n422));
  OAI21_X1  g221(.A(new_n339), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n406), .B1(new_n423), .B2(new_n388), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n338), .B1(new_n339), .B2(new_n389), .ZN(new_n425));
  INV_X1    g224(.A(G228gat), .ZN(new_n426));
  INV_X1    g225(.A(G233gat), .ZN(new_n427));
  OAI22_X1  g226(.A1(new_n424), .A2(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n389), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n351), .B1(KEYINPUT29), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n338), .A2(new_n339), .A3(new_n379), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n426), .A2(new_n427), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n430), .A2(new_n380), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(KEYINPUT80), .A2(G22gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(G78gat), .B(G106gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT31), .B(G50gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  MUX2_X1   g236(.A(G22gat), .B(new_n434), .S(new_n437), .Z(new_n438));
  AND3_X1   g237(.A1(new_n428), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n438), .B1(new_n428), .B2(new_n433), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n420), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n413), .A2(new_n414), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT6), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n361), .B(KEYINPUT81), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n404), .A2(new_n408), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(new_n413), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n410), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n353), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT37), .B1(new_n345), .B2(new_n348), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT37), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n352), .A2(new_n454), .A3(new_n347), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n453), .A2(new_n455), .A3(new_n328), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT38), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT38), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n453), .A2(new_n458), .A3(new_n455), .A4(new_n328), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT82), .B(KEYINPUT39), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n397), .A2(new_n398), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n363), .B(new_n461), .C1(new_n462), .C2(new_n391), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n407), .A2(new_n363), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n412), .B2(new_n362), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n447), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n449), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n463), .A2(new_n467), .A3(KEYINPUT40), .A4(new_n447), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n354), .A2(new_n470), .A3(new_n356), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n441), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n324), .B(new_n443), .C1(new_n460), .C2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n321), .A2(new_n441), .A3(new_n322), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT35), .B1(new_n420), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n313), .A2(new_n319), .ZN(new_n477));
  XOR2_X1   g276(.A(KEYINPUT83), .B(KEYINPUT35), .Z(new_n478));
  AND2_X1   g277(.A1(new_n450), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n477), .A2(new_n357), .A3(new_n441), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT84), .B1(new_n474), .B2(new_n481), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT98), .ZN(new_n485));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G71gat), .B(G78gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n490), .A2(KEYINPUT21), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT94), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G183gat), .B(G211gat), .Z(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT16), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(G1gat), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n499), .B(KEYINPUT92), .C1(G1gat), .C2(new_n497), .ZN(new_n500));
  INV_X1    g299(.A(G8gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT93), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n500), .B(G8gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n490), .A2(KEYINPUT21), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(G127gat), .B(G155gat), .Z(new_n509));
  NAND2_X1  g308(.A1(G231gat), .A2(G233gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n508), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n496), .B(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  INV_X1    g315(.A(G36gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(KEYINPUT89), .ZN(new_n519));
  NOR3_X1   g318(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT89), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n514), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT90), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g324(.A1(G43gat), .A2(G50gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G43gat), .A2(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT86), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n526), .A2(new_n530), .A3(new_n527), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(KEYINPUT15), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT90), .B(new_n514), .C1(new_n519), .C2(new_n522), .ZN(new_n533));
  INV_X1    g332(.A(new_n528), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT88), .B(G36gat), .Z(new_n536));
  AOI22_X1  g335(.A1(new_n534), .A2(new_n535), .B1(new_n536), .B2(G29gat), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n525), .A2(new_n532), .A3(new_n533), .A4(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n536), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n514), .B1(new_n520), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n542));
  OAI22_X1  g341(.A1(new_n539), .A2(new_n516), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(KEYINPUT15), .A3(new_n531), .A4(new_n529), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n538), .A2(new_n544), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI211_X1 g349(.A(KEYINPUT91), .B(KEYINPUT17), .C1(new_n538), .C2(new_n544), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n502), .B(new_n546), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n503), .A2(new_n506), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n548), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n552), .A2(KEYINPUT18), .A3(new_n553), .A4(new_n555), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n503), .A2(new_n506), .A3(new_n545), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n553), .B(KEYINPUT13), .Z(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n559), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G113gat), .B(G141gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G197gat), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT11), .B(G169gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT12), .Z(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n564), .A2(KEYINPUT85), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n570), .B1(new_n564), .B2(KEYINPUT85), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n579), .A2(KEYINPUT97), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n581), .A2(new_n582), .B1(G85gat), .B2(G92gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(KEYINPUT96), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n586), .B1(new_n583), .B2(new_n584), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G99gat), .B(G106gat), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n595), .A2(new_n603), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n545), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n606), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n546), .B(new_n605), .C1(new_n550), .C2(new_n551), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n607), .A2(new_n612), .A3(new_n608), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n580), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n578), .B(KEYINPUT97), .Z(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n613), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n490), .A3(new_n604), .ZN(new_n619));
  INV_X1    g418(.A(new_n490), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n603), .B1(new_n595), .B2(new_n599), .ZN(new_n621));
  INV_X1    g420(.A(new_n599), .ZN(new_n622));
  AOI211_X1 g421(.A(new_n601), .B(new_n622), .C1(new_n591), .C2(new_n594), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n490), .A4(new_n604), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G230gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n427), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n619), .A2(new_n624), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n630), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n632), .A2(new_n634), .A3(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR4_X1   g441(.A1(new_n513), .A2(new_n574), .A3(new_n618), .A4(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n484), .A2(new_n485), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n474), .A2(new_n481), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT84), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n474), .A2(KEYINPUT84), .A3(new_n481), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n647), .A2(new_n643), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n419), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT99), .B(G1gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1324gat));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  INV_X1    g455(.A(new_n357), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n485), .B1(new_n484), .B2(new_n643), .ZN(new_n658));
  AND4_X1   g457(.A1(new_n485), .A2(new_n647), .A3(new_n648), .A4(new_n643), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G8gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT16), .B(G8gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n651), .A2(new_n657), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n656), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  AOI211_X1 g464(.A(new_n357), .B(new_n662), .C1(new_n644), .C2(new_n650), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT100), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n501), .B1(new_n651), .B2(new_n657), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n669), .B2(new_n666), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n664), .A2(new_n656), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(new_n651), .ZN(new_n675));
  INV_X1    g474(.A(new_n477), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n675), .A2(G15gat), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n675), .B2(new_n324), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(G1326gat));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n651), .A2(new_n442), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n683), .A3(new_n680), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1327gat));
  NAND2_X1  g488(.A1(new_n481), .A2(KEYINPUT104), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n476), .A2(new_n691), .A3(new_n480), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n446), .A2(new_n417), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n415), .A2(KEYINPUT78), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n411), .A3(new_n695), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n696), .A2(new_n410), .B1(new_n354), .B2(new_n356), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT102), .B1(new_n697), .B2(new_n441), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n452), .A2(new_n457), .A3(new_n459), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n472), .A3(new_n441), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT102), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n420), .A2(new_n701), .A3(new_n442), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n698), .A2(new_n700), .A3(new_n324), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n420), .B2(new_n442), .ZN(new_n706));
  AOI211_X1 g505(.A(KEYINPUT102), .B(new_n441), .C1(new_n357), .C2(new_n419), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n472), .A2(new_n441), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n709), .A2(new_n699), .B1(new_n323), .B2(new_n320), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n705), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n693), .B1(new_n704), .B2(new_n711), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n618), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n647), .A2(new_n648), .A3(new_n618), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n642), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n513), .A2(new_n573), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n721), .B2(new_n419), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723));
  INV_X1    g522(.A(new_n618), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n482), .A2(new_n483), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n720), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n652), .A2(new_n516), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OR3_X1    g527(.A1(new_n726), .A2(new_n723), .A3(new_n727), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n722), .A2(new_n728), .A3(new_n729), .ZN(G1328gat));
  OAI21_X1  g529(.A(new_n536), .B1(new_n721), .B2(new_n357), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n657), .A2(new_n539), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT46), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n732), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n731), .A2(new_n733), .A3(new_n734), .ZN(G1329gat));
  NOR2_X1   g534(.A1(new_n676), .A2(G43gat), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n726), .A2(new_n737), .B1(KEYINPUT106), .B2(KEYINPUT47), .ZN(new_n738));
  INV_X1    g537(.A(new_n324), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n717), .A2(new_n739), .A3(new_n720), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(G43gat), .ZN(new_n741));
  AND2_X1   g540(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1330gat));
  NAND2_X1  g542(.A1(new_n442), .A2(G50gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n721), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n726), .ZN(new_n746));
  AOI21_X1  g545(.A(G50gat), .B1(new_n746), .B2(new_n442), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT48), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n747), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n749), .B(new_n750), .C1(new_n721), .C2(new_n744), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1331gat));
  INV_X1    g551(.A(new_n513), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n753), .A2(new_n574), .A3(new_n724), .A4(new_n642), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n703), .A2(KEYINPUT103), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n708), .A2(new_n710), .A3(new_n705), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(new_n693), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n652), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT107), .B(G57gat), .Z(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1332gat));
  AOI21_X1  g560(.A(new_n357), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT108), .Z(new_n763));
  NAND2_X1  g562(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT109), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(G1333gat));
  NAND2_X1  g566(.A1(new_n758), .A2(new_n739), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n676), .A2(G71gat), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n768), .A2(G71gat), .B1(new_n758), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g570(.A1(new_n758), .A2(new_n442), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT110), .B(G78gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n753), .A2(new_n573), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n642), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n717), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n419), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n712), .A2(new_n618), .A3(new_n775), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n712), .A2(new_n782), .A3(new_n618), .A4(new_n775), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n642), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n652), .A2(new_n597), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(G1336gat));
  INV_X1    g585(.A(new_n713), .ZN(new_n787));
  AOI211_X1 g586(.A(new_n724), .B(new_n787), .C1(new_n757), .C2(new_n693), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n725), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n657), .B(new_n777), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n776), .B1(new_n714), .B2(new_n716), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(KEYINPUT111), .A3(new_n657), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(G92gat), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n357), .A2(G92gat), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n642), .A3(new_n783), .A4(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n798), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n598), .B1(new_n794), .B2(new_n657), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT52), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n778), .B2(new_n324), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n676), .A2(G99gat), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n784), .B2(new_n807), .ZN(G1338gat));
  OAI21_X1  g607(.A(G106gat), .B1(new_n778), .B2(new_n441), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n442), .A2(new_n811), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n809), .B(new_n810), .C1(new_n784), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n784), .A2(new_n812), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n811), .B1(new_n794), .B2(new_n442), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT53), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n564), .A2(KEYINPUT85), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n569), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n626), .A2(new_n627), .A3(new_n630), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n632), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n630), .B1(new_n626), .B2(new_n627), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n638), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(KEYINPUT55), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n641), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(new_n821), .B2(new_n824), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n564), .A2(KEYINPUT85), .A3(new_n570), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n819), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT112), .B1(new_n561), .B2(new_n562), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  INV_X1    g631(.A(new_n562), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n555), .A2(new_n832), .A3(new_n560), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n553), .B1(new_n552), .B2(new_n555), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n568), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n558), .A2(new_n570), .A3(new_n563), .A4(new_n559), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n642), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n618), .B1(new_n830), .B2(new_n839), .ZN(new_n840));
  AND4_X1   g639(.A1(new_n618), .A2(new_n828), .A3(new_n838), .A4(new_n837), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n513), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n753), .A2(new_n574), .A3(new_n724), .A4(new_n718), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n475), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n652), .A3(new_n357), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n574), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(KEYINPUT113), .B2(new_n205), .ZN(new_n848));
  XNOR2_X1  g647(.A(KEYINPUT113), .B(G113gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(G1340gat));
  NOR2_X1   g649(.A1(new_n846), .A2(new_n718), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(new_n203), .ZN(G1341gat));
  NOR2_X1   g651(.A1(new_n846), .A2(new_n513), .ZN(new_n853));
  XOR2_X1   g652(.A(new_n853), .B(G127gat), .Z(G1342gat));
  NOR3_X1   g653(.A1(new_n724), .A2(new_n657), .A3(KEYINPUT114), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT114), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n618), .B2(new_n357), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n652), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n844), .A2(G134gat), .A3(new_n475), .A4(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n846), .B2(new_n724), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n324), .A2(new_n652), .A3(new_n357), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n442), .A2(KEYINPUT57), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n573), .A2(new_n828), .B1(KEYINPUT115), .B2(new_n839), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n839), .A2(KEYINPUT115), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n618), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n513), .B1(new_n869), .B2(new_n841), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n866), .B1(new_n870), .B2(new_n843), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n842), .A2(new_n843), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n872), .B2(new_n442), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n573), .B(new_n865), .C1(new_n871), .C2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n863), .B1(new_n874), .B2(G141gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n442), .ZN(new_n876));
  NOR4_X1   g675(.A1(new_n876), .A2(G141gat), .A3(new_n574), .A4(new_n864), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n877), .B1(new_n874), .B2(G141gat), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n875), .A2(new_n878), .A3(KEYINPUT58), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  AOI221_X4 g679(.A(new_n877), .B1(new_n863), .B2(new_n880), .C1(new_n874), .C2(G141gat), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n881), .ZN(G1344gat));
  NOR2_X1   g681(.A1(new_n871), .A2(new_n873), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n864), .ZN(new_n884));
  AOI211_X1 g683(.A(KEYINPUT59), .B(new_n375), .C1(new_n884), .C2(new_n642), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n843), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n442), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n844), .A2(new_n866), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n642), .B(new_n865), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n886), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  INV_X1    g690(.A(new_n876), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n865), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n642), .A2(new_n375), .ZN(new_n894));
  OAI22_X1  g693(.A1(new_n885), .A2(new_n891), .B1(new_n893), .B2(new_n894), .ZN(G1345gat));
  NOR2_X1   g694(.A1(new_n893), .A2(new_n513), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT117), .ZN(new_n897));
  AOI21_X1  g696(.A(G155gat), .B1(new_n896), .B2(KEYINPUT117), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n513), .A2(new_n368), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n897), .A2(new_n898), .B1(new_n884), .B2(new_n899), .ZN(G1346gat));
  XNOR2_X1  g699(.A(KEYINPUT76), .B(G162gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n324), .A2(new_n901), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n876), .A2(new_n858), .A3(new_n902), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n883), .A2(new_n724), .A3(new_n864), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n901), .ZN(G1347gat));
  NOR2_X1   g704(.A1(new_n652), .A2(new_n357), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n676), .ZN(new_n908));
  OR2_X1    g707(.A1(new_n908), .A2(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(KEYINPUT118), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n872), .A2(new_n441), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n244), .A3(new_n574), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n844), .A2(new_n475), .A3(new_n907), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n573), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(new_n244), .ZN(G1348gat));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n245), .A3(new_n642), .ZN(new_n916));
  OAI21_X1  g715(.A(G176gat), .B1(new_n911), .B2(new_n718), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1349gat));
  NOR2_X1   g717(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n919));
  AND2_X1   g718(.A1(KEYINPUT120), .A2(KEYINPUT60), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n909), .A2(new_n441), .A3(new_n910), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n844), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n923), .A3(new_n753), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT119), .B1(new_n911), .B2(new_n513), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(G183gat), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n913), .A2(new_n222), .A3(new_n225), .A4(new_n753), .ZN(new_n927));
  AOI211_X1 g726(.A(new_n919), .B(new_n920), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  AND4_X1   g727(.A1(KEYINPUT120), .A2(new_n926), .A3(KEYINPUT60), .A4(new_n927), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n229), .A3(new_n618), .ZN(new_n931));
  XOR2_X1   g730(.A(new_n931), .B(KEYINPUT121), .Z(new_n932));
  AOI21_X1  g731(.A(new_n229), .B1(new_n922), .B2(new_n618), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  OR3_X1    g733(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT61), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT61), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n933), .A2(new_n934), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n932), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n739), .A2(new_n907), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n892), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n573), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n939), .B(KEYINPUT123), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT124), .Z(new_n944));
  AND3_X1   g743(.A1(new_n944), .A2(G197gat), .A3(new_n573), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n888), .A2(new_n889), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n942), .B1(new_n945), .B2(new_n947), .ZN(G1352gat));
  NAND3_X1  g747(.A1(new_n947), .A2(new_n642), .A3(new_n944), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G204gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n940), .A2(G204gat), .A3(new_n718), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1353gat));
  NOR3_X1   g752(.A1(new_n940), .A2(G211gat), .A3(new_n513), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT125), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n943), .A2(new_n513), .ZN(new_n956));
  OAI21_X1  g755(.A(G211gat), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT63), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n959), .B(G211gat), .C1(new_n946), .C2(new_n956), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(new_n958), .A3(new_n960), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n941), .B2(new_n618), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n618), .A2(G218gat), .ZN(new_n963));
  XOR2_X1   g762(.A(new_n963), .B(KEYINPUT126), .Z(new_n964));
  AND2_X1   g763(.A1(new_n944), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n965), .B2(new_n947), .ZN(G1355gat));
endmodule


