

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U547 ( .A1(G2104), .A2(G2105), .ZN(n538) );
  NOR2_X1 U548 ( .A1(n933), .A2(n725), .ZN(n727) );
  OR2_X1 U549 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U550 ( .A1(n718), .A2(n719), .ZN(n761) );
  NAND2_X1 U551 ( .A1(n889), .A2(G137), .ZN(n541) );
  XNOR2_X1 U552 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n532) );
  NOR2_X1 U553 ( .A1(G164), .A2(G1384), .ZN(n719) );
  NOR2_X1 U554 ( .A1(G651), .A2(n645), .ZN(n651) );
  NOR2_X2 U555 ( .A1(n544), .A2(n543), .ZN(G160) );
  XOR2_X1 U556 ( .A(KEYINPUT75), .B(n525), .Z(n517) );
  XOR2_X1 U557 ( .A(n741), .B(KEYINPUT28), .Z(n518) );
  OR2_X1 U558 ( .A1(n761), .A2(n734), .ZN(n735) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n743) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n756) );
  NAND2_X1 U561 ( .A1(G160), .A2(G40), .ZN(n721) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n807) );
  NOR2_X1 U563 ( .A1(n645), .A2(n523), .ZN(n657) );
  INV_X1 U564 ( .A(KEYINPUT17), .ZN(n537) );
  INV_X1 U565 ( .A(G2105), .ZN(n539) );
  AND2_X1 U566 ( .A1(n539), .A2(G2104), .ZN(n888) );
  XNOR2_X1 U567 ( .A(n533), .B(n532), .ZN(n536) );
  XNOR2_X1 U568 ( .A(n531), .B(n530), .ZN(G168) );
  XNOR2_X1 U569 ( .A(KEYINPUT7), .B(KEYINPUT76), .ZN(n531) );
  NOR2_X2 U570 ( .A1(G543), .A2(G651), .ZN(n652) );
  NAND2_X1 U571 ( .A1(n652), .A2(G89), .ZN(n519) );
  XNOR2_X1 U572 ( .A(n519), .B(KEYINPUT4), .ZN(n521) );
  XOR2_X1 U573 ( .A(G543), .B(KEYINPUT0), .Z(n645) );
  XNOR2_X1 U574 ( .A(G651), .B(KEYINPUT67), .ZN(n523) );
  NAND2_X1 U575 ( .A1(G76), .A2(n657), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U577 ( .A(KEYINPUT5), .B(n522), .ZN(n529) );
  NOR2_X1 U578 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X2 U579 ( .A(KEYINPUT1), .B(n524), .Z(n655) );
  NAND2_X1 U580 ( .A1(G63), .A2(n655), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n651), .A2(G51), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n517), .A2(n526), .ZN(n527) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(n527), .Z(n528) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U585 ( .A1(G101), .A2(n888), .ZN(n533) );
  NOR2_X1 U586 ( .A1(n539), .A2(G2104), .ZN(n534) );
  XNOR2_X2 U587 ( .A(n534), .B(KEYINPUT64), .ZN(n893) );
  NAND2_X1 U588 ( .A1(G125), .A2(n893), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n544) );
  XNOR2_X2 U590 ( .A(n538), .B(n537), .ZN(n889) );
  AND2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U592 ( .A1(G113), .A2(n892), .ZN(n540) );
  NAND2_X1 U593 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U594 ( .A(n542), .B(KEYINPUT66), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G102), .A2(n888), .ZN(n545) );
  XNOR2_X1 U596 ( .A(n545), .B(KEYINPUT92), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G114), .A2(n892), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT91), .B(n546), .Z(n547) );
  NAND2_X1 U599 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U600 ( .A1(n889), .A2(G138), .ZN(n550) );
  NAND2_X1 U601 ( .A1(G126), .A2(n893), .ZN(n549) );
  NAND2_X1 U602 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U603 ( .A1(n552), .A2(n551), .ZN(G164) );
  XOR2_X1 U604 ( .A(G2446), .B(KEYINPUT104), .Z(n554) );
  XNOR2_X1 U605 ( .A(G2451), .B(G2430), .ZN(n553) );
  XNOR2_X1 U606 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U607 ( .A(n555), .B(G2427), .Z(n557) );
  XNOR2_X1 U608 ( .A(G1348), .B(G1341), .ZN(n556) );
  XNOR2_X1 U609 ( .A(n557), .B(n556), .ZN(n561) );
  XOR2_X1 U610 ( .A(G2443), .B(G2435), .Z(n559) );
  XNOR2_X1 U611 ( .A(G2438), .B(G2454), .ZN(n558) );
  XNOR2_X1 U612 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U613 ( .A(n561), .B(n560), .Z(n562) );
  AND2_X1 U614 ( .A1(G14), .A2(n562), .ZN(G401) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U616 ( .A1(G123), .A2(n893), .ZN(n564) );
  XNOR2_X1 U617 ( .A(KEYINPUT80), .B(KEYINPUT18), .ZN(n563) );
  XNOR2_X1 U618 ( .A(n564), .B(n563), .ZN(n571) );
  NAND2_X1 U619 ( .A1(G99), .A2(n888), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G135), .A2(n889), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G111), .A2(n892), .ZN(n567) );
  XNOR2_X1 U623 ( .A(KEYINPUT81), .B(n567), .ZN(n568) );
  NOR2_X1 U624 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n571), .A2(n570), .ZN(n992) );
  XNOR2_X1 U626 ( .A(G2096), .B(n992), .ZN(n572) );
  OR2_X1 U627 ( .A1(G2100), .A2(n572), .ZN(G156) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G69), .ZN(G235) );
  INV_X1 U630 ( .A(G108), .ZN(G238) );
  INV_X1 U631 ( .A(G120), .ZN(G236) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U634 ( .A(G223), .B(KEYINPUT71), .ZN(n827) );
  NAND2_X1 U635 ( .A1(n827), .A2(G567), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U637 ( .A1(n655), .A2(G56), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n575), .Z(n582) );
  NAND2_X1 U639 ( .A1(G81), .A2(n652), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT12), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT72), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G68), .A2(n657), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n651), .A2(G43), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n933) );
  XNOR2_X1 U648 ( .A(G860), .B(KEYINPUT73), .ZN(n611) );
  OR2_X1 U649 ( .A1(n933), .A2(n611), .ZN(G153) );
  NAND2_X1 U650 ( .A1(G52), .A2(n651), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G64), .A2(n655), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n591) );
  NAND2_X1 U653 ( .A1(n652), .A2(G90), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G77), .A2(n657), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U656 ( .A(KEYINPUT9), .B(n589), .Z(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U658 ( .A(KEYINPUT70), .B(n592), .ZN(G171) );
  INV_X1 U659 ( .A(G171), .ZN(G301) );
  NAND2_X1 U660 ( .A1(G301), .A2(G868), .ZN(n602) );
  NAND2_X1 U661 ( .A1(G92), .A2(n652), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G54), .A2(n651), .ZN(n594) );
  NAND2_X1 U663 ( .A1(G66), .A2(n655), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n657), .A2(G79), .ZN(n595) );
  XOR2_X1 U666 ( .A(KEYINPUT74), .B(n595), .Z(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X2 U669 ( .A(n600), .B(KEYINPUT15), .ZN(n936) );
  OR2_X1 U670 ( .A1(n936), .A2(G868), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n602), .A2(n601), .ZN(G284) );
  XOR2_X1 U672 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U673 ( .A1(G53), .A2(n651), .ZN(n604) );
  NAND2_X1 U674 ( .A1(G65), .A2(n655), .ZN(n603) );
  NAND2_X1 U675 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U676 ( .A1(n652), .A2(G91), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G78), .A2(n657), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n930) );
  INV_X1 U680 ( .A(n930), .ZN(G299) );
  NAND2_X1 U681 ( .A1(G868), .A2(G286), .ZN(n610) );
  INV_X1 U682 ( .A(G868), .ZN(n673) );
  NAND2_X1 U683 ( .A1(G299), .A2(n673), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U685 ( .A1(G559), .A2(n611), .ZN(n612) );
  XOR2_X1 U686 ( .A(KEYINPUT77), .B(n612), .Z(n613) );
  NAND2_X1 U687 ( .A1(n613), .A2(n936), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U689 ( .A1(n936), .A2(G868), .ZN(n615) );
  XOR2_X1 U690 ( .A(KEYINPUT79), .B(n615), .Z(n616) );
  NOR2_X1 U691 ( .A1(G559), .A2(n616), .ZN(n619) );
  NOR2_X1 U692 ( .A1(G868), .A2(n933), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT78), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G559), .A2(n936), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n620), .B(n933), .ZN(n671) );
  NOR2_X1 U697 ( .A1(n671), .A2(G860), .ZN(n629) );
  NAND2_X1 U698 ( .A1(n652), .A2(G93), .ZN(n622) );
  NAND2_X1 U699 ( .A1(G80), .A2(n657), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT82), .B(n623), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G55), .A2(n651), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G67), .A2(n655), .ZN(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U705 ( .A(KEYINPUT83), .B(n626), .Z(n627) );
  OR2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n674) );
  XOR2_X1 U707 ( .A(n629), .B(n674), .Z(G145) );
  NAND2_X1 U708 ( .A1(G50), .A2(n651), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G62), .A2(n655), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U711 ( .A(KEYINPUT84), .B(n632), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G75), .A2(n657), .ZN(n633) );
  XNOR2_X1 U713 ( .A(KEYINPUT85), .B(n633), .ZN(n634) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n652), .A2(G88), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(G303) );
  INV_X1 U717 ( .A(G303), .ZN(G166) );
  NAND2_X1 U718 ( .A1(G48), .A2(n651), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G86), .A2(n652), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n657), .A2(G73), .ZN(n640) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n640), .Z(n641) );
  NOR2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G61), .A2(n655), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G87), .A2(n645), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U729 ( .A1(n655), .A2(n648), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(G49), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U732 ( .A1(G47), .A2(n651), .ZN(n654) );
  NAND2_X1 U733 ( .A1(G85), .A2(n652), .ZN(n653) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n655), .A2(G60), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(KEYINPUT68), .ZN(n659) );
  NAND2_X1 U737 ( .A1(G72), .A2(n657), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U739 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U740 ( .A(KEYINPUT69), .B(n662), .ZN(G290) );
  XOR2_X1 U741 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n664) );
  XNOR2_X1 U742 ( .A(KEYINPUT88), .B(KEYINPUT86), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n664), .B(n663), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n930), .B(G305), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(G288), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n669) );
  XOR2_X1 U747 ( .A(G290), .B(n674), .Z(n668) );
  XNOR2_X1 U748 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U749 ( .A(G166), .B(n670), .ZN(n833) );
  XNOR2_X1 U750 ( .A(n671), .B(n833), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n672), .A2(G868), .ZN(n676) );
  NAND2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U759 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U760 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n682) );
  NAND2_X1 U761 ( .A1(G132), .A2(G82), .ZN(n681) );
  XNOR2_X1 U762 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U763 ( .A1(n683), .A2(G218), .ZN(n684) );
  NAND2_X1 U764 ( .A1(G96), .A2(n684), .ZN(n831) );
  NAND2_X1 U765 ( .A1(n831), .A2(G2106), .ZN(n689) );
  NOR2_X1 U766 ( .A1(G236), .A2(G238), .ZN(n686) );
  NOR2_X1 U767 ( .A1(G235), .A2(G237), .ZN(n685) );
  NAND2_X1 U768 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U769 ( .A(KEYINPUT90), .B(n687), .ZN(n832) );
  NAND2_X1 U770 ( .A1(n832), .A2(G567), .ZN(n688) );
  NAND2_X1 U771 ( .A1(n689), .A2(n688), .ZN(n908) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U773 ( .A1(n908), .A2(n690), .ZN(n830) );
  NAND2_X1 U774 ( .A1(n830), .A2(G36), .ZN(G176) );
  NOR2_X1 U775 ( .A1(n719), .A2(n721), .ZN(n822) );
  XNOR2_X1 U776 ( .A(KEYINPUT37), .B(G2067), .ZN(n820) );
  NAND2_X1 U777 ( .A1(G104), .A2(n888), .ZN(n692) );
  NAND2_X1 U778 ( .A1(G140), .A2(n889), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n694) );
  XOR2_X1 U780 ( .A(KEYINPUT34), .B(KEYINPUT93), .Z(n693) );
  XNOR2_X1 U781 ( .A(n694), .B(n693), .ZN(n699) );
  NAND2_X1 U782 ( .A1(G116), .A2(n892), .ZN(n696) );
  NAND2_X1 U783 ( .A1(G128), .A2(n893), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U785 ( .A(KEYINPUT35), .B(n697), .Z(n698) );
  NOR2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U787 ( .A(KEYINPUT36), .B(n700), .ZN(n866) );
  NOR2_X1 U788 ( .A1(n820), .A2(n866), .ZN(n1001) );
  NAND2_X1 U789 ( .A1(n822), .A2(n1001), .ZN(n818) );
  NAND2_X1 U790 ( .A1(G105), .A2(n888), .ZN(n701) );
  XNOR2_X1 U791 ( .A(n701), .B(KEYINPUT38), .ZN(n708) );
  NAND2_X1 U792 ( .A1(n889), .A2(G141), .ZN(n703) );
  NAND2_X1 U793 ( .A1(G129), .A2(n893), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n892), .A2(G117), .ZN(n704) );
  XOR2_X1 U796 ( .A(KEYINPUT94), .B(n704), .Z(n705) );
  NOR2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U799 ( .A(KEYINPUT95), .B(n709), .Z(n867) );
  NAND2_X1 U800 ( .A1(G1996), .A2(n867), .ZN(n717) );
  NAND2_X1 U801 ( .A1(G95), .A2(n888), .ZN(n711) );
  NAND2_X1 U802 ( .A1(G119), .A2(n893), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U804 ( .A1(G107), .A2(n892), .ZN(n713) );
  NAND2_X1 U805 ( .A1(G131), .A2(n889), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n879) );
  NAND2_X1 U808 ( .A1(G1991), .A2(n879), .ZN(n716) );
  NAND2_X1 U809 ( .A1(n717), .A2(n716), .ZN(n990) );
  NAND2_X1 U810 ( .A1(n822), .A2(n990), .ZN(n813) );
  NAND2_X1 U811 ( .A1(n818), .A2(n813), .ZN(n806) );
  INV_X1 U812 ( .A(n721), .ZN(n718) );
  AND2_X1 U813 ( .A1(n761), .A2(G1341), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n719), .A2(G1996), .ZN(n720) );
  NOR2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U816 ( .A(n722), .B(KEYINPUT26), .ZN(n723) );
  NOR2_X1 U817 ( .A1(n727), .A2(n936), .ZN(n726) );
  XNOR2_X1 U818 ( .A(n726), .B(KEYINPUT97), .ZN(n733) );
  NAND2_X1 U819 ( .A1(n727), .A2(n936), .ZN(n731) );
  INV_X1 U820 ( .A(n761), .ZN(n745) );
  NOR2_X1 U821 ( .A1(n745), .A2(G1348), .ZN(n729) );
  NOR2_X1 U822 ( .A1(G2067), .A2(n761), .ZN(n728) );
  NOR2_X1 U823 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n739) );
  INV_X1 U826 ( .A(G2072), .ZN(n734) );
  XNOR2_X1 U827 ( .A(n735), .B(KEYINPUT27), .ZN(n737) );
  INV_X1 U828 ( .A(G1956), .ZN(n963) );
  NOR2_X1 U829 ( .A1(n963), .A2(n745), .ZN(n736) );
  NOR2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n930), .A2(n740), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n930), .A2(n740), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n518), .ZN(n744) );
  XNOR2_X1 U835 ( .A(n744), .B(n743), .ZN(n749) );
  INV_X1 U836 ( .A(G1961), .ZN(n973) );
  NAND2_X1 U837 ( .A1(n761), .A2(n973), .ZN(n747) );
  XNOR2_X1 U838 ( .A(G2078), .B(KEYINPUT25), .ZN(n913) );
  NAND2_X1 U839 ( .A1(n745), .A2(n913), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n747), .A2(n746), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n753), .A2(G171), .ZN(n748) );
  NAND2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n759) );
  NAND2_X1 U843 ( .A1(G8), .A2(n761), .ZN(n760) );
  NOR2_X1 U844 ( .A1(G1966), .A2(n760), .ZN(n774) );
  NOR2_X1 U845 ( .A1(G2084), .A2(n761), .ZN(n771) );
  NOR2_X1 U846 ( .A1(n774), .A2(n771), .ZN(n750) );
  NAND2_X1 U847 ( .A1(G8), .A2(n750), .ZN(n751) );
  XNOR2_X1 U848 ( .A(KEYINPUT30), .B(n751), .ZN(n752) );
  NOR2_X1 U849 ( .A1(G168), .A2(n752), .ZN(n755) );
  NOR2_X1 U850 ( .A1(n753), .A2(G171), .ZN(n754) );
  NOR2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n757) );
  XNOR2_X1 U852 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U853 ( .A1(n759), .A2(n758), .ZN(n772) );
  NAND2_X1 U854 ( .A1(n772), .A2(G286), .ZN(n766) );
  NOR2_X1 U855 ( .A1(G1971), .A2(n760), .ZN(n763) );
  NOR2_X1 U856 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U857 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n764), .A2(G303), .ZN(n765) );
  NAND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U860 ( .A(n767), .B(KEYINPUT98), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n768), .A2(G8), .ZN(n770) );
  XOR2_X1 U862 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n769) );
  XNOR2_X1 U863 ( .A(n770), .B(n769), .ZN(n792) );
  NAND2_X1 U864 ( .A1(G8), .A2(n771), .ZN(n776) );
  INV_X1 U865 ( .A(n772), .ZN(n773) );
  NOR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n793) );
  NAND2_X1 U868 ( .A1(G1976), .A2(G288), .ZN(n940) );
  INV_X1 U869 ( .A(n940), .ZN(n777) );
  OR2_X1 U870 ( .A1(n760), .A2(n777), .ZN(n781) );
  INV_X1 U871 ( .A(n781), .ZN(n778) );
  AND2_X1 U872 ( .A1(n793), .A2(n778), .ZN(n779) );
  AND2_X1 U873 ( .A1(n792), .A2(n779), .ZN(n785) );
  NOR2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n787) );
  NOR2_X1 U875 ( .A1(G1971), .A2(G303), .ZN(n780) );
  NOR2_X1 U876 ( .A1(n787), .A2(n780), .ZN(n941) );
  OR2_X1 U877 ( .A1(n781), .A2(n941), .ZN(n783) );
  INV_X1 U878 ( .A(KEYINPUT33), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U880 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U881 ( .A(n786), .B(KEYINPUT100), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n787), .A2(KEYINPUT33), .ZN(n788) );
  NOR2_X1 U883 ( .A1(n760), .A2(n788), .ZN(n789) );
  NOR2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U885 ( .A(G1981), .B(G305), .Z(n947) );
  NAND2_X1 U886 ( .A1(n791), .A2(n947), .ZN(n799) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n796) );
  NOR2_X1 U888 ( .A1(G2090), .A2(G303), .ZN(n794) );
  NAND2_X1 U889 ( .A1(G8), .A2(n794), .ZN(n795) );
  NAND2_X1 U890 ( .A1(n796), .A2(n795), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n797), .A2(n760), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n804) );
  NOR2_X1 U893 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U894 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  XNOR2_X1 U895 ( .A(KEYINPUT96), .B(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n760), .A2(n802), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n808), .B(n807), .ZN(n810) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n938) );
  NAND2_X1 U901 ( .A1(n938), .A2(n822), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n825) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n867), .ZN(n996) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n879), .ZN(n991) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n991), .A2(n811), .ZN(n812) );
  XOR2_X1 U907 ( .A(KEYINPUT102), .B(n812), .Z(n814) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U909 ( .A(KEYINPUT103), .B(n815), .ZN(n816) );
  NOR2_X1 U910 ( .A1(n996), .A2(n816), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n820), .A2(n866), .ZN(n1005) );
  NAND2_X1 U914 ( .A1(n821), .A2(n1005), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U917 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U920 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U924 ( .A(G132), .ZN(G219) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U929 ( .A(n936), .B(n933), .ZN(n834) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n836) );
  XNOR2_X1 U931 ( .A(G286), .B(G301), .ZN(n835) );
  XNOR2_X1 U932 ( .A(n836), .B(n835), .ZN(n837) );
  NOR2_X1 U933 ( .A1(G37), .A2(n837), .ZN(G397) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1971), .B(G1956), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n857) );
  XOR2_X1 U946 ( .A(KEYINPUT105), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1961), .B(KEYINPUT106), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(G1976), .B(G1981), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1966), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT107), .B(G2474), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(G229) );
  NAND2_X1 U956 ( .A1(G100), .A2(n888), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G112), .A2(n892), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U959 ( .A1(G136), .A2(n889), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT108), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n893), .A2(G124), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n861), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U964 ( .A1(n865), .A2(n864), .ZN(G162) );
  XNOR2_X1 U965 ( .A(G162), .B(n866), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n878) );
  NAND2_X1 U967 ( .A1(G118), .A2(n892), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G130), .A2(n893), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U970 ( .A1(G106), .A2(n888), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G142), .A2(n889), .ZN(n871) );
  NAND2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U973 ( .A(n873), .B(KEYINPUT45), .Z(n874) );
  NOR2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n876), .B(n992), .ZN(n877) );
  XOR2_X1 U976 ( .A(n878), .B(n877), .Z(n887) );
  XNOR2_X1 U977 ( .A(KEYINPUT109), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n879), .B(KEYINPUT48), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(n882), .B(KEYINPUT111), .Z(n884) );
  XNOR2_X1 U981 ( .A(G160), .B(KEYINPUT112), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U983 ( .A(G164), .B(n885), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n900) );
  NAND2_X1 U985 ( .A1(G103), .A2(n888), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G139), .A2(n889), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n898) );
  NAND2_X1 U988 ( .A1(G115), .A2(n892), .ZN(n895) );
  NAND2_X1 U989 ( .A1(G127), .A2(n893), .ZN(n894) );
  NAND2_X1 U990 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U992 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U993 ( .A(KEYINPUT110), .B(n899), .Z(n1007) );
  XNOR2_X1 U994 ( .A(n900), .B(n1007), .ZN(n901) );
  NOR2_X1 U995 ( .A1(G37), .A2(n901), .ZN(G395) );
  NOR2_X1 U996 ( .A1(G401), .A2(n908), .ZN(n905) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n902) );
  XNOR2_X1 U998 ( .A(KEYINPUT49), .B(n902), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G397), .A2(n903), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n906) );
  NOR2_X1 U1001 ( .A1(n906), .A2(G395), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n907), .B(KEYINPUT113), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(n908), .ZN(G319) );
  XOR2_X1 U1005 ( .A(G2084), .B(G34), .Z(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT54), .B(n909), .ZN(n926) );
  XNOR2_X1 U1007 ( .A(G2090), .B(G35), .ZN(n924) );
  XOR2_X1 U1008 ( .A(G1991), .B(G25), .Z(n910) );
  NAND2_X1 U1009 ( .A1(n910), .A2(G28), .ZN(n920) );
  XNOR2_X1 U1010 ( .A(G2067), .B(G26), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(G33), .B(G2072), .ZN(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n918) );
  XOR2_X1 U1013 ( .A(n913), .B(G27), .Z(n916) );
  INV_X1 U1014 ( .A(G1996), .ZN(n914) );
  XOR2_X1 U1015 ( .A(n914), .B(G32), .Z(n915) );
  NOR2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1019 ( .A(KEYINPUT117), .B(n921), .Z(n922) );
  XNOR2_X1 U1020 ( .A(n922), .B(KEYINPUT53), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(KEYINPUT118), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n928), .B(KEYINPUT55), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(G29), .A2(n929), .ZN(n987) );
  XNOR2_X1 U1026 ( .A(G16), .B(KEYINPUT56), .ZN(n955) );
  XNOR2_X1 U1027 ( .A(n930), .B(G1956), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(G171), .B(G1961), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(G1341), .B(n933), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n953) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n936), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n937), .B(KEYINPUT119), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n946) );
  AND2_X1 U1035 ( .A1(G303), .A2(G1971), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(KEYINPUT120), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n951) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G168), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1042 ( .A(KEYINPUT57), .B(n949), .Z(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1045 ( .A1(n955), .A2(n954), .ZN(n985) );
  INV_X1 U1046 ( .A(G16), .ZN(n983) );
  XNOR2_X1 U1047 ( .A(G1986), .B(G24), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(G1971), .B(G22), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(G23), .B(G1976), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(KEYINPUT123), .B(n958), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1053 ( .A(n961), .B(KEYINPUT124), .Z(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT58), .B(n962), .ZN(n980) );
  XOR2_X1 U1055 ( .A(G1341), .B(G19), .Z(n965) );
  XNOR2_X1 U1056 ( .A(n963), .B(G20), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n971) );
  XOR2_X1 U1058 ( .A(G1981), .B(G6), .Z(n969) );
  XOR2_X1 U1059 ( .A(G1348), .B(G4), .Z(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT121), .B(n966), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(n967), .B(KEYINPUT59), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT60), .B(n972), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(n973), .B(G5), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G21), .B(G1966), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT122), .B(n978), .Z(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(KEYINPUT61), .B(n981), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1073 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1074 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1075 ( .A1(G11), .A2(n988), .ZN(n989) );
  XOR2_X1 U1076 ( .A(KEYINPUT125), .B(n989), .Z(n1019) );
  NOR2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n993) );
  NAND2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n999) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n994) );
  XNOR2_X1 U1080 ( .A(KEYINPUT114), .B(n994), .ZN(n995) );
  NOR2_X1 U1081 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1082 ( .A(KEYINPUT51), .B(n997), .ZN(n998) );
  NOR2_X1 U1083 ( .A1(n999), .A2(n998), .ZN(n1003) );
  XOR2_X1 U1084 ( .A(G160), .B(G2084), .Z(n1000) );
  NOR2_X1 U1085 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1086 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1087 ( .A(n1004), .B(KEYINPUT115), .ZN(n1006) );
  NAND2_X1 U1088 ( .A1(n1006), .A2(n1005), .ZN(n1012) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n1009) );
  XNOR2_X1 U1090 ( .A(G2072), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1091 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1092 ( .A(KEYINPUT50), .B(n1010), .Z(n1011) );
  NOR2_X1 U1093 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1094 ( .A(KEYINPUT52), .B(n1013), .ZN(n1015) );
  INV_X1 U1095 ( .A(KEYINPUT55), .ZN(n1014) );
  NAND2_X1 U1096 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1097 ( .A1(n1016), .A2(G29), .ZN(n1017) );
  XOR2_X1 U1098 ( .A(n1017), .B(KEYINPUT116), .Z(n1018) );
  NOR2_X1 U1099 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1100 ( .A(KEYINPUT62), .B(n1020), .Z(n1021) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1021), .Z(G311) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

