//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT26), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n210), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n219), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n217), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n215), .A2(new_n216), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT23), .B1(new_n208), .B2(new_n209), .ZN(new_n225));
  OR3_X1    g024(.A1(new_n216), .A2(KEYINPUT66), .A3(KEYINPUT24), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(new_n219), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n230), .B(new_n216), .C1(KEYINPUT66), .C2(KEYINPUT24), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n225), .A2(new_n226), .A3(new_n228), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT25), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n211), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n216), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n230), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n238), .A2(new_n239), .A3(new_n228), .A4(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n233), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n246));
  INV_X1    g045(.A(G120gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n247), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n249), .A2(G120gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n246), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(G127gat), .A2(G134gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G127gat), .A2(G134gat), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT1), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n251), .ZN(new_n258));
  NOR2_X1   g057(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n259));
  OAI21_X1  g058(.A(G120gat), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n253), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264));
  INV_X1    g063(.A(G134gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(G127gat), .ZN(new_n266));
  OAI221_X1 g065(.A(new_n255), .B1(new_n264), .B2(KEYINPUT1), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n245), .A2(new_n268), .ZN(new_n269));
  AND4_X1   g068(.A1(new_n239), .A2(new_n236), .A3(new_n243), .A4(new_n237), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n228), .A2(new_n270), .B1(new_n232), .B2(KEYINPUT25), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n271), .A2(new_n224), .B1(new_n263), .B2(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n205), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT33), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT32), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n245), .A2(new_n268), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n263), .A2(new_n267), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n271), .A3(new_n224), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n281), .B2(new_n205), .ZN(new_n282));
  XOR2_X1   g081(.A(G15gat), .B(G43gat), .Z(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n275), .A2(new_n276), .A3(new_n282), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n205), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n287), .B1(new_n278), .B2(new_n280), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n276), .B(new_n285), .C1(new_n288), .C2(KEYINPUT33), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n273), .A2(KEYINPUT32), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n281), .B2(new_n205), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT34), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(KEYINPUT72), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n278), .A2(new_n280), .A3(new_n287), .A4(new_n295), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n286), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n286), .B2(new_n291), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n300), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n202), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G211gat), .ZN(new_n305));
  INV_X1    g104(.A(G218gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G211gat), .A2(G218gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n315));
  XNOR2_X1  g114(.A(G197gat), .B(G204gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n314), .B(new_n320), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(new_n316), .A3(new_n310), .A4(new_n312), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT76), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT76), .B1(new_n319), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G141gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n326), .A2(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(G141gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT79), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(G141gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(G148gat), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT79), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G155gat), .B(G162gat), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G155gat), .ZN(new_n339));
  INV_X1    g138(.A(G162gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n331), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n342), .B1(new_n332), .B2(new_n333), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n347));
  OAI21_X1  g146(.A(new_n325), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G228gat), .A2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n319), .A2(new_n322), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(KEYINPUT29), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n345), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G22gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n351), .B1(new_n352), .B2(new_n347), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n345), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n348), .A2(new_n365), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n349), .B(KEYINPUT83), .Z(new_n367));
  OAI211_X1 g166(.A(new_n355), .B(new_n363), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n348), .A2(new_n350), .A3(new_n354), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n348), .B2(new_n365), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n362), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n286), .A2(new_n291), .ZN(new_n373));
  INV_X1    g172(.A(new_n297), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n286), .A2(new_n291), .A3(new_n297), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(KEYINPUT73), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(KEYINPUT89), .A3(new_n302), .ZN(new_n378));
  INV_X1    g177(.A(new_n325), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT77), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n245), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n383), .B1(new_n245), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n379), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n245), .A2(new_n383), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n347), .B1(new_n271), .B2(new_n224), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n325), .B(new_n387), .C1(new_n388), .C2(new_n381), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT30), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  INV_X1    g191(.A(G64gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G92gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n390), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n390), .A2(new_n397), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n386), .A2(new_n389), .A3(new_n396), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n343), .B1(new_n336), .B2(new_n337), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n404), .A2(new_n263), .A3(new_n267), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n263), .A2(new_n267), .B1(new_n338), .B2(new_n344), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n404), .A2(new_n351), .B1(new_n263), .B2(new_n267), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n345), .A2(KEYINPUT3), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n413), .B1(new_n268), .B2(new_n345), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n404), .A2(KEYINPUT4), .A3(new_n263), .A4(new_n267), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n412), .A2(new_n402), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT5), .ZN(new_n417));
  OAI211_X1 g216(.A(KEYINPUT80), .B(new_n403), .C1(new_n405), .C2(new_n406), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n409), .A2(new_n416), .A3(new_n417), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n414), .A2(new_n415), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n417), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n402), .A3(new_n412), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G1gat), .B(G29gat), .Z(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G57gat), .B(G85gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n419), .A2(new_n429), .A3(new_n423), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n435));
  AOI221_X4 g234(.A(KEYINPUT35), .B1(new_n398), .B2(new_n401), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n304), .A2(new_n372), .A3(new_n378), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n401), .A2(new_n398), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n432), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n429), .B1(new_n419), .B2(new_n423), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n435), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n375), .A2(new_n372), .A3(new_n376), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT35), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(KEYINPUT90), .B(KEYINPUT35), .C1(new_n443), .C2(new_n444), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n437), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n377), .A2(new_n450), .A3(new_n302), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n298), .A2(new_n299), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT36), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n372), .B(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n451), .A2(new_n453), .B1(new_n443), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n404), .A2(new_n351), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n268), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n404), .A2(new_n351), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n403), .B1(new_n420), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n405), .A2(new_n406), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n461), .B(KEYINPUT39), .C1(new_n403), .C2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n464), .B(new_n403), .C1(new_n420), .C2(new_n460), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n465), .A2(new_n466), .A3(new_n429), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n466), .B1(new_n465), .B2(new_n429), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n469), .A2(KEYINPUT87), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n438), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n431), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT88), .B1(new_n469), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n465), .A2(new_n429), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT86), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n465), .A2(new_n466), .A3(new_n429), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT40), .A4(new_n463), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT87), .B1(new_n469), .B2(new_n470), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n473), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n397), .B1(new_n390), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n484), .B2(new_n390), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n486), .A2(KEYINPUT38), .B1(new_n390), .B2(new_n397), .ZN(new_n487));
  OR3_X1    g286(.A1(new_n379), .A2(new_n382), .A3(new_n385), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n388), .A2(new_n381), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n383), .B2(new_n245), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n488), .B(KEYINPUT37), .C1(new_n490), .C2(new_n325), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n487), .A2(new_n493), .A3(new_n435), .A4(new_n434), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n372), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n456), .B1(new_n483), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n449), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n498));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n499), .A2(G1gat), .ZN(new_n500));
  INV_X1    g299(.A(G8gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT16), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n502), .B2(G1gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n500), .B2(new_n503), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n498), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(KEYINPUT92), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  OR3_X1    g311(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n513), .A2(KEYINPUT91), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  NOR3_X1   g314(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT91), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n512), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  OAI22_X1  g320(.A1(new_n511), .A2(KEYINPUT15), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n513), .A2(new_n515), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  OAI22_X1  g322(.A1(new_n519), .A2(new_n522), .B1(new_n512), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n510), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT93), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n527), .A3(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n524), .B(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n508), .A3(new_n504), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n530), .B(KEYINPUT13), .Z(new_n536));
  AND2_X1   g335(.A1(new_n526), .A2(new_n528), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n510), .A2(new_n524), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n529), .A2(new_n532), .A3(KEYINPUT18), .A4(new_n530), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT11), .B(G169gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G197gat), .ZN(new_n543));
  XOR2_X1   g342(.A(G113gat), .B(G141gat), .Z(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT12), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n535), .A2(new_n539), .A3(new_n546), .A4(new_n540), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n497), .A2(KEYINPUT94), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT94), .B1(new_n497), .B2(new_n550), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT100), .ZN(new_n554));
  INV_X1    g353(.A(G99gat), .ZN(new_n555));
  INV_X1    g354(.A(G106gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(KEYINPUT8), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT99), .B(G92gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(G85gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n554), .B(new_n559), .C1(new_n562), .C2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n558), .A2(KEYINPUT8), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n395), .A2(KEYINPUT99), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G85gat), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n559), .A2(new_n554), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n557), .A2(KEYINPUT100), .A3(new_n558), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n563), .B(KEYINPUT7), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .A4(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n531), .A2(new_n566), .A3(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n566), .A2(new_n577), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n580), .B2(new_n524), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(G190gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n582), .A2(G190gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n306), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(G218gat), .A3(new_n583), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT98), .ZN(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n589), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(new_n305), .ZN(new_n595));
  INV_X1    g394(.A(new_n510), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(G64gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n393), .A2(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT96), .ZN(new_n601));
  NAND2_X1  g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT9), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n602), .A2(KEYINPUT95), .ZN(new_n608));
  OR2_X1    g407(.A1(G71gat), .A2(G78gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n602), .A2(KEYINPUT95), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n602), .B1(new_n609), .B2(new_n603), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n393), .A2(KEYINPUT97), .A3(G57gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n598), .A3(new_n616), .ZN(new_n617));
  AOI22_X1  g416(.A1(new_n607), .A2(new_n612), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(G183gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n596), .A2(new_n229), .A3(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n621), .B2(new_n622), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n595), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  INV_X1    g428(.A(new_n595), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n628), .A2(new_n631), .A3(new_n635), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n593), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G230gat), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(new_n204), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n605), .B1(new_n598), .B2(new_n599), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n611), .B1(new_n646), .B2(new_n604), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n617), .A2(new_n613), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n566), .B(new_n577), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n580), .A2(new_n618), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT101), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n580), .A2(new_n652), .A3(new_n618), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT10), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n643), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n653), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n657), .B1(new_n643), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT102), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G120gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n328), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n659), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n640), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n553), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n434), .A2(new_n435), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  OAI211_X1 g469(.A(new_n472), .B(new_n665), .C1(new_n551), .C2(new_n552), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n673), .B(new_n674), .C1(new_n675), .C2(G8gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n671), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n675), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n676), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT104), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n676), .A2(new_n678), .A3(new_n682), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1325gat));
  AND2_X1   g483(.A1(new_n304), .A2(new_n378), .ZN(new_n685));
  AOI21_X1  g484(.A(G15gat), .B1(new_n666), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n666), .A2(G15gat), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n451), .A2(new_n453), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n686), .B1(new_n688), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n666), .A2(new_n455), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(new_n639), .ZN(new_n695));
  INV_X1    g494(.A(new_n592), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n589), .B(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n664), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT105), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n553), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n520), .A3(new_n668), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n497), .A2(new_n697), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n695), .A2(KEYINPUT106), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n639), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n664), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(KEYINPUT107), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n497), .A2(new_n697), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n706), .A2(new_n550), .A3(new_n710), .A4(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G29gat), .B1(new_n714), .B2(new_n667), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n703), .A2(new_n715), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n521), .A3(new_n472), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n717), .A2(KEYINPUT46), .ZN(new_n718));
  OAI21_X1  g517(.A(G36gat), .B1(new_n714), .B2(new_n438), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(KEYINPUT46), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(G1329gat));
  INV_X1    g520(.A(G43gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n701), .A2(new_n722), .A3(new_n685), .ZN(new_n723));
  OAI21_X1  g522(.A(G43gat), .B1(new_n714), .B2(new_n689), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1330gat));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  INV_X1    g527(.A(G50gat), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n729), .B(new_n700), .C1(new_n551), .C2(new_n552), .ZN(new_n730));
  INV_X1    g529(.A(new_n455), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  OAI21_X1  g533(.A(G50gat), .B1(new_n714), .B2(new_n731), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n593), .B1(new_n449), .B2(new_n496), .ZN(new_n737));
  INV_X1    g536(.A(new_n705), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n713), .B(new_n550), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n710), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n739), .A2(new_n372), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n729), .B1(new_n741), .B2(KEYINPUT108), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n714), .B2(new_n372), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n732), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n728), .B(new_n736), .C1(new_n745), .C2(new_n734), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n738), .B1(new_n497), .B2(new_n697), .ZN(new_n747));
  INV_X1    g546(.A(new_n712), .ZN(new_n748));
  AOI211_X1 g547(.A(new_n593), .B(new_n748), .C1(new_n449), .C2(new_n496), .ZN(new_n749));
  INV_X1    g548(.A(new_n550), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n372), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n751), .A2(KEYINPUT108), .A3(new_n752), .A4(new_n710), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n744), .A2(new_n753), .A3(G50gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n734), .B1(new_n754), .B2(new_n733), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT109), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n746), .A2(new_n757), .ZN(G1331gat));
  AOI211_X1 g557(.A(new_n550), .B(new_n640), .C1(new_n449), .C2(new_n496), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n664), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n760), .A2(new_n667), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(new_n597), .ZN(G1332gat));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n438), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  INV_X1    g566(.A(new_n760), .ZN(new_n768));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n769), .A3(new_n685), .ZN(new_n770));
  OAI21_X1  g569(.A(G71gat), .B1(new_n760), .B2(new_n689), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g572(.A1(new_n768), .A2(new_n455), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n639), .A2(new_n550), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n706), .A2(new_n664), .A3(new_n713), .A4(new_n776), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n777), .A2(new_n572), .A3(new_n667), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  AND4_X1   g582(.A1(new_n737), .A2(new_n782), .A3(new_n776), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n782), .B1(new_n737), .B2(new_n776), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n784), .A2(new_n698), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n668), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n778), .B1(new_n572), .B2(new_n787), .ZN(G1336gat));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n395), .A3(new_n472), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n561), .B1(new_n777), .B2(new_n438), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT52), .ZN(G1337gat));
  OR3_X1    g591(.A1(new_n777), .A2(KEYINPUT111), .A3(new_n689), .ZN(new_n793));
  OAI21_X1  g592(.A(KEYINPUT111), .B1(new_n777), .B2(new_n689), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(G99gat), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n786), .A2(new_n555), .A3(new_n685), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1338gat));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n786), .A2(new_n556), .A3(new_n752), .ZN(new_n799));
  OAI21_X1  g598(.A(G106gat), .B1(new_n777), .B2(new_n731), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n803));
  OAI21_X1  g602(.A(G106gat), .B1(new_n777), .B2(new_n372), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(KEYINPUT113), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n803), .A2(new_n798), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(new_n806), .A3(new_n807), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n707), .A2(new_n709), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n658), .A2(new_n655), .ZN(new_n810));
  INV_X1    g609(.A(new_n656), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n642), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n812), .A2(KEYINPUT54), .A3(new_n657), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT114), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n812), .A2(new_n657), .A3(new_n815), .A4(KEYINPUT54), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n657), .A2(KEYINPUT54), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n663), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n659), .A2(new_n663), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n663), .A4(new_n818), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n821), .A2(new_n550), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n537), .A2(new_n538), .A3(new_n536), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n530), .B1(new_n529), .B2(new_n532), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n545), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n549), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n664), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n697), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n828), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n593), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n809), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n665), .A2(new_n750), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n731), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n667), .A2(new_n472), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(KEYINPUT115), .A3(new_n731), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n838), .A2(new_n685), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n750), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n835), .A2(new_n668), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n843), .A2(new_n472), .A3(new_n444), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n550), .C1(new_n259), .C2(new_n258), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n841), .B2(new_n698), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n247), .A3(new_n664), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1341gat));
  NOR3_X1   g648(.A1(new_n841), .A2(new_n266), .A3(new_n809), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n844), .A2(new_n639), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n266), .B2(new_n851), .ZN(G1342gat));
  NOR2_X1   g651(.A1(new_n843), .A2(new_n444), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n593), .A2(new_n472), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT116), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n265), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT56), .Z(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n841), .B2(new_n593), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1343gat));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n829), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n828), .A2(KEYINPUT117), .A3(new_n664), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n824), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n593), .ZN(new_n864));
  INV_X1    g663(.A(new_n832), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n639), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n834), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n455), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT57), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n689), .A2(new_n839), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n372), .B1(new_n833), .B2(new_n834), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n869), .A2(new_n873), .A3(new_n550), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT118), .B1(new_n874), .B2(G141gat), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(KEYINPUT58), .ZN(new_n876));
  INV_X1    g675(.A(new_n871), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n870), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n750), .A2(G141gat), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n874), .A2(G141gat), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n876), .B(new_n880), .ZN(G1344gat));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n328), .A3(new_n664), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n869), .A2(new_n873), .A3(new_n664), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(G148gat), .ZN(new_n885));
  INV_X1    g684(.A(new_n870), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n832), .B1(new_n593), .B2(new_n863), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n834), .B1(new_n887), .B2(new_n639), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n888), .B2(new_n455), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n872), .B(new_n372), .C1(new_n833), .C2(new_n834), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n664), .B(new_n886), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n884), .B1(new_n891), .B2(G148gat), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n882), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT119), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n895), .B(new_n882), .C1(new_n885), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(G1345gat));
  NAND2_X1  g696(.A1(new_n869), .A2(new_n873), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n339), .A3(new_n809), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n639), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT120), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n901), .B2(new_n339), .ZN(G1346gat));
  NAND3_X1  g701(.A1(new_n855), .A2(new_n340), .A3(new_n752), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n843), .A2(new_n903), .A3(new_n690), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n869), .A2(new_n697), .A3(new_n873), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G162gat), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT121), .ZN(G1347gat));
  NAND3_X1  g706(.A1(new_n452), .A2(new_n472), .A3(new_n372), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n668), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n835), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT123), .ZN(new_n913));
  INV_X1    g712(.A(G169gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n550), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT124), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n668), .A2(new_n438), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n838), .A2(new_n685), .A3(new_n840), .A4(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(G169gat), .B1(new_n918), .B2(new_n750), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1348gat));
  INV_X1    g719(.A(G176gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n918), .A2(new_n921), .A3(new_n698), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(KEYINPUT125), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(KEYINPUT125), .ZN(new_n924));
  AOI21_X1  g723(.A(G176gat), .B1(new_n913), .B2(new_n664), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n918), .B2(new_n809), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n639), .A2(new_n220), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n912), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n918), .B2(new_n593), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT126), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n933), .B(G190gat), .C1(new_n918), .C2(new_n593), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(KEYINPUT61), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n913), .A2(new_n219), .A3(new_n697), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(KEYINPUT126), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(G1351gat));
  NAND2_X1  g738(.A1(new_n689), .A2(new_n917), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n877), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(G197gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(new_n550), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n889), .A2(new_n890), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n944), .A2(new_n940), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n550), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n947), .B2(new_n942), .ZN(G1352gat));
  INV_X1    g747(.A(G204gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n949), .A3(new_n664), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(KEYINPUT62), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n944), .A2(new_n698), .A3(new_n940), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G204gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(G1353gat));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n305), .A3(new_n639), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n945), .A2(new_n639), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G1354gat));
  NAND3_X1  g761(.A1(new_n941), .A2(new_n306), .A3(new_n697), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n697), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n965), .B2(new_n306), .ZN(G1355gat));
endmodule


