//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986;
  AND2_X1   g000(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n203));
  OAI21_X1  g002(.A(G162gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT76), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT2), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G141gat), .B(G148gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n206), .A2(new_n208), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n209), .B1(new_n211), .B2(KEYINPUT74), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  OAI221_X1 g017(.A(new_n216), .B1(KEYINPUT74), .B2(new_n209), .C1(new_n218), .C2(new_n213), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221));
  INV_X1    g020(.A(G113gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G120gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(G120gat), .ZN(new_n224));
  INV_X1    g023(.A(G120gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G127gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G134gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G134gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(G127gat), .B2(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT67), .A2(G134gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(G127gat), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n231), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n222), .A2(G120gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n225), .A2(G113gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n232), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n229), .A2(new_n235), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n220), .A2(KEYINPUT4), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT68), .B1(new_n225), .B2(G113gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(new_n241), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT69), .B1(new_n247), .B2(new_n226), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n227), .A2(new_n228), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n235), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n239), .A2(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n215), .A2(new_n219), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n245), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(G225gat), .A2(G233gat), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n244), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n208), .A2(new_n214), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n207), .B1(new_n204), .B2(KEYINPUT2), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n257), .B(new_n219), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n215), .A2(KEYINPUT77), .A3(new_n257), .A4(new_n219), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n253), .A2(KEYINPUT3), .B1(new_n251), .B2(new_n250), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n264), .B2(new_n265), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n256), .B(KEYINPUT5), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G1gat), .B(G29gat), .Z(new_n270));
  XNOR2_X1  g069(.A(G57gat), .B(G85gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n244), .A2(new_n254), .A3(new_n255), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n264), .A2(new_n265), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT78), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n252), .B(new_n253), .ZN(new_n282));
  INV_X1    g081(.A(new_n255), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n269), .B(new_n275), .C1(new_n280), .C2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n269), .B1(new_n280), .B2(new_n284), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n274), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(new_n286), .A3(new_n285), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n289), .B1(new_n288), .B2(new_n274), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G204gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G197gat), .ZN(new_n295));
  INV_X1    g094(.A(G197gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G204gat), .ZN(new_n297));
  INV_X1    g096(.A(G211gat), .ZN(new_n298));
  INV_X1    g097(.A(G218gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n295), .B(new_n297), .C1(new_n300), .C2(KEYINPUT22), .ZN(new_n301));
  XNOR2_X1  g100(.A(G211gat), .B(G218gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n303), .A2(KEYINPUT81), .A3(KEYINPUT29), .ZN(new_n304));
  INV_X1    g103(.A(new_n302), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n301), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT81), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n304), .A2(new_n309), .A3(new_n257), .ZN(new_n310));
  AOI22_X1  g109(.A1(new_n310), .A2(new_n253), .B1(G228gat), .B2(G233gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n306), .B1(new_n264), .B2(new_n307), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n220), .B1(new_n257), .B2(new_n308), .ZN(new_n315));
  OAI211_X1 g114(.A(G228gat), .B(G233gat), .C1(new_n312), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT31), .B(G50gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(G22gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n317), .B(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n323));
  INV_X1    g122(.A(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT66), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G183gat), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT24), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NOR2_X1   g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT65), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(G169gat), .B2(G176gat), .ZN(new_n343));
  NAND3_X1  g142(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n335), .A2(new_n338), .A3(new_n345), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n331), .A2(new_n333), .B1(new_n324), .B2(new_n328), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(KEYINPUT23), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n339), .A3(new_n343), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n336), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT27), .B(G183gat), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n352), .A2(KEYINPUT28), .A3(new_n328), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT27), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n325), .B2(new_n327), .ZN(new_n355));
  NOR2_X1   g154(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n328), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT28), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n353), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n337), .B(KEYINPUT26), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n339), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n330), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n351), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n323), .B1(new_n363), .B2(new_n252), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n252), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n323), .A3(new_n252), .ZN(new_n367));
  INV_X1    g166(.A(G227gat), .ZN(new_n368));
  INV_X1    g167(.A(G233gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n363), .A2(new_n323), .A3(new_n252), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n371), .B1(new_n365), .B2(new_n364), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n368), .A2(new_n369), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n373), .B(KEYINPUT64), .Z(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT34), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n370), .A2(KEYINPUT34), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G15gat), .B(G43gat), .Z(new_n378));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n374), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n366), .B2(new_n367), .ZN(new_n382));
  XOR2_X1   g181(.A(KEYINPUT71), .B(KEYINPUT33), .Z(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n380), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT32), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n366), .A2(new_n367), .ZN(new_n389));
  AOI221_X4 g188(.A(new_n386), .B1(new_n384), .B2(new_n380), .C1(new_n389), .C2(new_n374), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n377), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT32), .B1(new_n372), .B2(new_n381), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n383), .B1(new_n372), .B2(new_n381), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n380), .ZN(new_n394));
  INV_X1    g193(.A(new_n380), .ZN(new_n395));
  OAI221_X1 g194(.A(KEYINPUT32), .B1(new_n383), .B2(new_n395), .C1(new_n372), .C2(new_n381), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n376), .A3(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n322), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  AND2_X1   g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n363), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n363), .B2(new_n307), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n401), .A2(new_n402), .A3(new_n303), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT72), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n303), .B1(new_n401), .B2(new_n402), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  OAI211_X1 g206(.A(KEYINPUT72), .B(new_n303), .C1(new_n401), .C2(new_n402), .ZN(new_n408));
  XOR2_X1   g207(.A(G8gat), .B(G36gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT73), .ZN(new_n410));
  XOR2_X1   g209(.A(G64gat), .B(G92gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n413), .B1(new_n406), .B2(new_n408), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n405), .A2(new_n404), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n363), .A2(new_n307), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n400), .B(new_n306), .C1(new_n417), .C2(new_n399), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n416), .A2(new_n408), .A3(new_n418), .A4(new_n413), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT30), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n414), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n293), .A2(new_n398), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT35), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n421), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n288), .A2(new_n274), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT80), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n285), .A2(new_n286), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n290), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n425), .B1(new_n429), .B2(new_n287), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(KEYINPUT35), .A3(new_n398), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n322), .ZN(new_n433));
  INV_X1    g232(.A(new_n293), .ZN(new_n434));
  INV_X1    g233(.A(new_n419), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT38), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n412), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n418), .A2(new_n405), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(KEYINPUT37), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n416), .A2(new_n408), .A3(new_n418), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(KEYINPUT37), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n435), .B1(new_n441), .B2(KEYINPUT83), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n440), .A2(KEYINPUT37), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(new_n439), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n413), .B1(new_n440), .B2(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n436), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n433), .B1(new_n434), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n244), .A2(new_n254), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n267), .B2(new_n268), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n283), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n278), .A2(new_n279), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n255), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  OR2_X1    g256(.A1(new_n282), .A2(new_n283), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT39), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n455), .B(new_n274), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT40), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n453), .A2(new_n283), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(KEYINPUT39), .A3(new_n458), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(KEYINPUT40), .A3(new_n274), .A4(new_n455), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n285), .B(new_n414), .C1(new_n415), .C2(new_n420), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n451), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n467), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(KEYINPUT82), .A3(new_n465), .A4(new_n462), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n450), .A2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n394), .A2(new_n376), .A3(new_n396), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n376), .B1(new_n394), .B2(new_n396), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT36), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n391), .A2(new_n476), .A3(new_n397), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n293), .A2(new_n421), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(new_n433), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n432), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G50gat), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT15), .B1(new_n482), .B2(G43gat), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(G43gat), .B2(new_n482), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(G29gat), .B2(G36gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT86), .B(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(G43gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(G43gat), .B2(new_n482), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n487), .A2(new_n488), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n486), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OR3_X1    g291(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n485), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G29gat), .A2(G36gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(KEYINPUT85), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n493), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n494), .A2(KEYINPUT85), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n484), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(KEYINPUT16), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n508), .B2(new_n507), .ZN(new_n510));
  INV_X1    g309(.A(G8gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n503), .A2(new_n512), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT18), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(new_n517), .A3(new_n515), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT18), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n503), .A2(new_n512), .ZN(new_n524));
  MUX2_X1   g323(.A(new_n523), .B(new_n522), .S(new_n524), .Z(new_n525));
  XOR2_X1   g324(.A(new_n517), .B(KEYINPUT13), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n518), .A2(new_n521), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(G169gat), .B(G197gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT84), .B(KEYINPUT11), .Z(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT12), .Z(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n534), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n518), .A2(new_n521), .A3(new_n527), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n481), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n541));
  XNOR2_X1  g340(.A(G134gat), .B(G162gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT92), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT7), .ZN(new_n545));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(KEYINPUT8), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n548), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT91), .B(G92gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(G85gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(G99gat), .B(G106gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n554), .B1(new_n504), .B2(new_n505), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n503), .ZN(new_n557));
  AND2_X1   g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT41), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G190gat), .B(G218gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n558), .A2(KEYINPUT41), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n562), .B1(new_n555), .B2(new_n560), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n566), .B1(new_n564), .B2(new_n567), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n544), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n564), .A2(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n565), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n573), .A2(new_n568), .A3(new_n543), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT89), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  OR2_X1    g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n580), .B(new_n581), .C1(new_n577), .C2(new_n582), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n512), .B1(new_n586), .B2(KEYINPUT21), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT90), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI211_X1 g390(.A(G231gat), .B(G233gat), .C1(new_n586), .C2(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n585), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT21), .ZN(new_n594));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n597), .B1(new_n592), .B2(new_n596), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n591), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n590), .A3(new_n598), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n588), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n603), .A3(new_n588), .ZN(new_n606));
  XOR2_X1   g405(.A(G183gat), .B(G211gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n610), .B2(new_n604), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n541), .B1(new_n576), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n609), .A2(new_n611), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(KEYINPUT93), .A3(new_n575), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT94), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n554), .B2(new_n586), .ZN(new_n617));
  INV_X1    g416(.A(new_n553), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n552), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(KEYINPUT94), .A3(new_n593), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n618), .B1(new_n552), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(KEYINPUT95), .B(new_n553), .C1(new_n549), .C2(new_n551), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n586), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n617), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n586), .A2(KEYINPUT10), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(new_n619), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n554), .A2(KEYINPUT96), .A3(KEYINPUT10), .A4(new_n586), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n617), .A2(new_n620), .A3(new_n636), .A4(new_n624), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n627), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G120gat), .B(G148gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT98), .ZN(new_n640));
  XOR2_X1   g439(.A(G176gat), .B(G204gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n630), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n635), .A2(new_n637), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n626), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n628), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n642), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n644), .A2(new_n645), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n645), .B1(new_n644), .B2(new_n649), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n540), .A2(new_n613), .A3(new_n615), .A4(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(new_n293), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n508), .ZN(G1324gat));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n421), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT42), .B1(new_n656), .B2(new_n511), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  MUX2_X1   g458(.A(KEYINPUT42), .B(new_n657), .S(new_n659), .Z(G1325gat));
  NOR3_X1   g459(.A1(new_n473), .A2(new_n474), .A3(KEYINPUT36), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n476), .B1(new_n391), .B2(new_n397), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G15gat), .B1(new_n653), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n473), .A2(new_n474), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(G15gat), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n664), .B1(new_n653), .B2(new_n667), .ZN(G1326gat));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n322), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NAND3_X1  g470(.A1(new_n652), .A2(new_n576), .A3(new_n612), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT100), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n540), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n674), .A2(G29gat), .A3(new_n293), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n675), .B(KEYINPUT45), .Z(new_n676));
  OAI21_X1  g475(.A(new_n663), .B1(new_n430), .B2(new_n322), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n677), .B1(new_n471), .B2(new_n450), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT44), .B(new_n576), .C1(new_n678), .C2(new_n432), .ZN(new_n679));
  INV_X1    g478(.A(new_n652), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(new_n539), .A3(new_n614), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n575), .A2(KEYINPUT101), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n571), .A2(new_n574), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n468), .A2(new_n470), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n443), .A2(new_n447), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n445), .B(new_n442), .C1(new_n688), .C2(new_n436), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n322), .B1(new_n689), .B2(new_n293), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n480), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n422), .A2(new_n423), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT35), .B1(new_n430), .B2(new_n398), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n686), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n679), .B(new_n681), .C1(KEYINPUT44), .C2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT102), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n481), .B2(new_n686), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n699), .A2(new_n700), .A3(new_n679), .A4(new_n681), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n434), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G29gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n676), .A2(new_n704), .ZN(G1328gat));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n425), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n702), .A2(KEYINPUT103), .A3(new_n425), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n708), .A2(G36gat), .A3(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n674), .A2(G36gat), .A3(new_n421), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT46), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1329gat));
  OAI21_X1  g512(.A(G43gat), .B1(new_n696), .B2(new_n663), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n666), .A2(G43gat), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n714), .B(KEYINPUT47), .C1(new_n674), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n674), .A2(new_n715), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n478), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(G43gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(KEYINPUT47), .ZN(G1330gat));
  XNOR2_X1  g519(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n697), .A2(new_n433), .A3(new_n701), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n540), .A2(new_n482), .A3(new_n433), .A4(new_n673), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT105), .B1(new_n722), .B2(G50gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G50gat), .B1(new_n696), .B2(new_n322), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1331gat));
  NAND3_X1  g529(.A1(new_n613), .A2(new_n615), .A3(new_n539), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n481), .A2(new_n652), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n434), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  INV_X1    g533(.A(KEYINPUT49), .ZN(new_n735));
  INV_X1    g534(.A(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n425), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT106), .Z(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n736), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1333gat));
  NAND2_X1  g540(.A1(new_n732), .A2(new_n478), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n666), .A2(G71gat), .ZN(new_n743));
  AOI22_X1  g542(.A1(new_n742), .A2(G71gat), .B1(new_n732), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n732), .A2(new_n433), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g546(.A1(new_n652), .A2(new_n614), .A3(new_n538), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n699), .A2(new_n679), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n749), .A2(new_n293), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G85gat), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n750), .A2(KEYINPUT107), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n614), .A2(new_n538), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n576), .B(new_n754), .C1(new_n678), .C2(new_n432), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT108), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n575), .B1(new_n691), .B2(new_n694), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT51), .A4(new_n754), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n755), .A2(new_n756), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n652), .A2(G85gat), .A3(new_n293), .ZN(new_n765));
  OAI22_X1  g564(.A1(new_n752), .A2(new_n753), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  NOR3_X1   g565(.A1(new_n652), .A2(G92gat), .A3(new_n421), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n699), .A2(new_n425), .A3(new_n679), .A4(new_n748), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n550), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n768), .A2(new_n774), .A3(new_n769), .A4(new_n771), .ZN(new_n775));
  INV_X1    g574(.A(new_n767), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n755), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT109), .B1(new_n758), .B2(new_n754), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n756), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n776), .B1(new_n780), .B2(new_n761), .ZN(new_n781));
  INV_X1    g580(.A(new_n771), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT110), .B(KEYINPUT52), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n755), .A2(new_n777), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n758), .A2(KEYINPUT109), .A3(new_n754), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n787), .A2(new_n756), .B1(new_n757), .B2(new_n760), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n771), .B1(new_n788), .B2(new_n776), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT110), .B1(new_n789), .B2(KEYINPUT52), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n773), .B(new_n775), .C1(new_n784), .C2(new_n790), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n749), .B2(new_n663), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n652), .A2(new_n666), .A3(G99gat), .ZN(new_n793));
  XOR2_X1   g592(.A(new_n793), .B(KEYINPUT112), .Z(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n764), .B2(new_n794), .ZN(G1338gat));
  OAI21_X1  g594(.A(G106gat), .B1(new_n749), .B2(new_n322), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n652), .A2(G106gat), .A3(new_n322), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT114), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n788), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT53), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n763), .A2(KEYINPUT115), .A3(new_n799), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT115), .B1(new_n763), .B2(new_n799), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n803), .B(new_n796), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n806), .ZN(G1339gat));
  NAND4_X1  g606(.A1(new_n613), .A2(new_n615), .A3(new_n539), .A4(new_n652), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n635), .A2(new_n637), .A3(new_n627), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n642), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(new_n638), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT116), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n811), .A2(new_n814), .A3(new_n818), .A4(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n815), .A2(new_n816), .B1(new_n630), .B2(new_n643), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n516), .A2(new_n517), .B1(new_n525), .B2(new_n526), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n533), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n537), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n685), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(new_n821), .A3(new_n538), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n650), .B2(new_n651), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n830), .B2(new_n685), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n809), .B1(new_n831), .B2(new_n612), .ZN(new_n832));
  INV_X1    g631(.A(new_n398), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n832), .A2(new_n293), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n421), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836), .B2(new_n538), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT117), .B1(new_n832), .B2(new_n433), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n685), .B1(new_n828), .B2(new_n829), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n571), .A2(new_n574), .A3(new_n683), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n683), .B1(new_n571), .B2(new_n574), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n826), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n822), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n612), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n808), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n322), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n434), .A2(new_n421), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n666), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n539), .A2(new_n222), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n837), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  AOI21_X1  g653(.A(G120gat), .B1(new_n836), .B2(new_n680), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n652), .A2(new_n225), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n852), .B2(new_n856), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n851), .B2(new_n612), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n230), .A3(new_n614), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  NOR2_X1   g659(.A1(new_n575), .A2(new_n425), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n834), .A2(new_n236), .A3(new_n237), .A4(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n862), .B2(KEYINPUT56), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n864), .A2(new_n865), .B1(KEYINPUT56), .B2(new_n862), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n851), .B2(new_n575), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n849), .A2(new_n478), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n845), .A2(new_n433), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n829), .A2(KEYINPUT119), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n826), .B(new_n874), .C1(new_n650), .C2(new_n651), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n828), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n843), .B1(new_n876), .B2(new_n575), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n808), .B1(new_n877), .B2(new_n614), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n872), .B1(new_n878), .B2(new_n433), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(G141gat), .A3(new_n538), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n663), .A2(new_n433), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT120), .Z(new_n883));
  NAND3_X1  g682(.A1(new_n845), .A2(new_n434), .A3(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n539), .A3(new_n425), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(G141gat), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n887), .B(new_n888), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n884), .A2(new_n425), .ZN(new_n890));
  INV_X1    g689(.A(G148gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n680), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n891), .C1(new_n880), .C2(new_n680), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n870), .A2(KEYINPUT57), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n823), .A2(KEYINPUT121), .A3(new_n576), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n822), .B2(new_n575), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n826), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n876), .A2(new_n575), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n614), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n872), .B(new_n433), .C1(new_n901), .C2(new_n809), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n895), .A2(new_n902), .A3(new_n680), .A4(new_n869), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n894), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n892), .B1(new_n893), .B2(new_n904), .ZN(G1345gat));
  NOR2_X1   g704(.A1(new_n202), .A2(new_n203), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n906), .A3(new_n614), .ZN(new_n907));
  INV_X1    g706(.A(new_n880), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n612), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n909), .B2(new_n906), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n908), .B2(new_n686), .ZN(new_n911));
  OR3_X1    g710(.A1(new_n575), .A2(G162gat), .A3(new_n425), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n884), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n832), .A2(new_n434), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n833), .A2(new_n421), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n538), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n434), .A2(new_n421), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n666), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n922), .B1(new_n838), .B2(new_n847), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n538), .A2(G169gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(G1348gat));
  INV_X1    g724(.A(G176gat), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n923), .B2(new_n680), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n916), .A2(G176gat), .A3(new_n652), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  AND4_X1   g728(.A1(new_n352), .A2(new_n914), .A3(new_n614), .A4(new_n915), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n923), .A2(new_n614), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT66), .B(G183gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n934), .A2(KEYINPUT122), .A3(KEYINPUT60), .ZN(new_n935));
  NOR2_X1   g734(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n936));
  AND2_X1   g735(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n935), .A2(new_n938), .ZN(G1350gat));
  AOI21_X1  g738(.A(new_n328), .B1(new_n923), .B2(new_n576), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT123), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT124), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n943), .A3(new_n941), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n846), .B1(new_n845), .B2(new_n322), .ZN(new_n945));
  AOI211_X1 g744(.A(KEYINPUT117), .B(new_n433), .C1(new_n844), .C2(new_n808), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n576), .B(new_n921), .C1(new_n945), .C2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G190gat), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT61), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n947), .A2(new_n941), .A3(G190gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT124), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n942), .A2(new_n944), .A3(new_n950), .A4(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n917), .A2(new_n328), .A3(new_n685), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1351gat));
  NOR2_X1   g754(.A1(new_n882), .A2(new_n421), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n914), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n538), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n895), .A2(new_n902), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n920), .A2(new_n478), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n539), .A2(new_n296), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(G1352gat));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n680), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT125), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n963), .A2(new_n968), .A3(new_n680), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n967), .A2(G204gat), .A3(new_n969), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n957), .A2(G204gat), .A3(new_n652), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1353gat));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n298), .A3(new_n614), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n895), .A2(new_n902), .A3(new_n614), .A4(new_n961), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n979), .B1(new_n976), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n974), .B1(new_n978), .B2(new_n980), .ZN(G1354gat));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n576), .B1(new_n963), .B2(new_n982), .ZN(new_n983));
  NOR3_X1   g782(.A1(new_n960), .A2(KEYINPUT127), .A3(new_n962), .ZN(new_n984));
  OAI21_X1  g783(.A(G218gat), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n958), .A2(new_n299), .A3(new_n685), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


