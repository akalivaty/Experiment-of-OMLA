

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U556 ( .A1(n541), .A2(G2104), .ZN(n888) );
  NOR2_X2 U557 ( .A1(G2104), .A2(n541), .ZN(n894) );
  NAND2_X1 U558 ( .A1(n750), .A2(n749), .ZN(n756) );
  INV_X1 U559 ( .A(KEYINPUT33), .ZN(n749) );
  XOR2_X1 U560 ( .A(KEYINPUT82), .B(n538), .Z(n521) );
  XOR2_X1 U561 ( .A(n747), .B(KEYINPUT96), .Z(n522) );
  NOR2_X1 U562 ( .A1(n693), .A2(n692), .ZN(n697) );
  INV_X1 U563 ( .A(KEYINPUT31), .ZN(n724) );
  XNOR2_X1 U564 ( .A(n725), .B(n724), .ZN(n726) );
  NAND2_X1 U565 ( .A1(n683), .A2(n798), .ZN(n728) );
  INV_X1 U566 ( .A(n764), .ZN(n748) );
  INV_X1 U567 ( .A(n976), .ZN(n753) );
  XNOR2_X1 U568 ( .A(KEYINPUT68), .B(KEYINPUT13), .ZN(n579) );
  NOR2_X1 U569 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U570 ( .A(n580), .B(n579), .ZN(n581) );
  NAND2_X1 U571 ( .A1(n756), .A2(n755), .ZN(n758) );
  NOR2_X1 U572 ( .A1(n630), .A2(n528), .ZN(n637) );
  XNOR2_X1 U573 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n555) );
  NOR2_X1 U574 ( .A1(G651), .A2(n630), .ZN(n647) );
  AND2_X1 U575 ( .A1(n585), .A2(n584), .ZN(n691) );
  XNOR2_X1 U576 ( .A(n556), .B(n555), .ZN(n557) );
  NOR2_X1 U577 ( .A1(n544), .A2(n543), .ZN(G164) );
  NOR2_X1 U578 ( .A1(G543), .A2(G651), .ZN(n523) );
  XNOR2_X1 U579 ( .A(n523), .B(KEYINPUT64), .ZN(n588) );
  NAND2_X1 U580 ( .A1(G89), .A2(n588), .ZN(n524) );
  XNOR2_X1 U581 ( .A(n524), .B(KEYINPUT4), .ZN(n526) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n630) );
  INV_X1 U583 ( .A(G651), .ZN(n528) );
  NAND2_X1 U584 ( .A1(G76), .A2(n637), .ZN(n525) );
  NAND2_X1 U585 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U586 ( .A(n527), .B(KEYINPUT5), .ZN(n534) );
  NOR2_X1 U587 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n529), .Z(n640) );
  NAND2_X1 U589 ( .A1(G63), .A2(n640), .ZN(n531) );
  NAND2_X1 U590 ( .A1(G51), .A2(n647), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U592 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U594 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U595 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U597 ( .A1(G114), .A2(n893), .ZN(n537) );
  INV_X1 U598 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U599 ( .A1(G126), .A2(n894), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U601 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT17), .B(n539), .Z(n553) );
  BUF_X1 U603 ( .A(n553), .Z(n889) );
  NAND2_X1 U604 ( .A1(n889), .A2(G138), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n521), .A2(n540), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G102), .A2(n888), .ZN(n542) );
  XNOR2_X1 U607 ( .A(KEYINPUT83), .B(n542), .ZN(n543) );
  NAND2_X1 U608 ( .A1(G72), .A2(n637), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G85), .A2(n588), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U611 ( .A1(G60), .A2(n640), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G47), .A2(n647), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U614 ( .A1(n550), .A2(n549), .ZN(G290) );
  NAND2_X1 U615 ( .A1(G113), .A2(n893), .ZN(n552) );
  NAND2_X1 U616 ( .A1(G125), .A2(n894), .ZN(n551) );
  AND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n679) );
  NAND2_X1 U618 ( .A1(G137), .A2(n553), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT66), .ZN(n558) );
  NAND2_X1 U620 ( .A1(G101), .A2(n888), .ZN(n556) );
  AND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n681) );
  AND2_X1 U622 ( .A1(n679), .A2(n681), .ZN(G160) );
  NAND2_X1 U623 ( .A1(G64), .A2(n640), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G52), .A2(n647), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U626 ( .A1(G77), .A2(n637), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G90), .A2(n588), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n563), .Z(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(G171) );
  AND2_X1 U631 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U632 ( .A(G132), .ZN(G219) );
  INV_X1 U633 ( .A(G82), .ZN(G220) );
  INV_X1 U634 ( .A(G108), .ZN(G238) );
  INV_X1 U635 ( .A(G120), .ZN(G236) );
  INV_X1 U636 ( .A(G57), .ZN(G237) );
  NAND2_X1 U637 ( .A1(G65), .A2(n640), .ZN(n567) );
  NAND2_X1 U638 ( .A1(G53), .A2(n647), .ZN(n566) );
  NAND2_X1 U639 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G78), .A2(n637), .ZN(n569) );
  NAND2_X1 U641 ( .A1(G91), .A2(n588), .ZN(n568) );
  NAND2_X1 U642 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U643 ( .A1(n571), .A2(n570), .ZN(n708) );
  INV_X1 U644 ( .A(n708), .ZN(G299) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U646 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U647 ( .A(G567), .ZN(n668) );
  NOR2_X1 U648 ( .A1(n668), .A2(G223), .ZN(n573) );
  XNOR2_X1 U649 ( .A(n573), .B(KEYINPUT11), .ZN(G234) );
  NAND2_X1 U650 ( .A1(n640), .A2(G56), .ZN(n574) );
  XNOR2_X1 U651 ( .A(n574), .B(KEYINPUT14), .ZN(n582) );
  NAND2_X1 U652 ( .A1(G68), .A2(n637), .ZN(n578) );
  XOR2_X1 U653 ( .A(KEYINPUT67), .B(KEYINPUT12), .Z(n576) );
  NAND2_X1 U654 ( .A1(G81), .A2(n588), .ZN(n575) );
  XNOR2_X1 U655 ( .A(n576), .B(n575), .ZN(n577) );
  NAND2_X1 U656 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U658 ( .A(n583), .B(KEYINPUT69), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G43), .A2(n647), .ZN(n584) );
  INV_X1 U660 ( .A(n691), .ZN(n996) );
  INV_X1 U661 ( .A(G860), .ZN(n621) );
  OR2_X1 U662 ( .A1(n996), .A2(n621), .ZN(G153) );
  XOR2_X1 U663 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U664 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U665 ( .A1(G66), .A2(n640), .ZN(n587) );
  NAND2_X1 U666 ( .A1(G79), .A2(n637), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n592) );
  NAND2_X1 U668 ( .A1(n647), .A2(G54), .ZN(n590) );
  NAND2_X1 U669 ( .A1(G92), .A2(n588), .ZN(n589) );
  NAND2_X1 U670 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U671 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U672 ( .A(KEYINPUT15), .B(n593), .Z(n980) );
  OR2_X1 U673 ( .A1(n980), .A2(G868), .ZN(n594) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(G284) );
  INV_X1 U675 ( .A(G868), .ZN(n658) );
  NOR2_X1 U676 ( .A1(G286), .A2(n658), .ZN(n597) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U678 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U679 ( .A1(G559), .A2(n621), .ZN(n598) );
  XOR2_X1 U680 ( .A(KEYINPUT71), .B(n598), .Z(n599) );
  NAND2_X1 U681 ( .A1(n599), .A2(n980), .ZN(n600) );
  XNOR2_X1 U682 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n996), .ZN(n603) );
  NAND2_X1 U684 ( .A1(G868), .A2(n980), .ZN(n601) );
  NOR2_X1 U685 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G111), .A2(n893), .ZN(n605) );
  NAND2_X1 U688 ( .A1(G99), .A2(n888), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G135), .A2(n889), .ZN(n606) );
  XNOR2_X1 U691 ( .A(n606), .B(KEYINPUT72), .ZN(n609) );
  NAND2_X1 U692 ( .A1(G123), .A2(n894), .ZN(n607) );
  XNOR2_X1 U693 ( .A(n607), .B(KEYINPUT18), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U695 ( .A1(n611), .A2(n610), .ZN(n931) );
  XNOR2_X1 U696 ( .A(n931), .B(G2096), .ZN(n613) );
  INV_X1 U697 ( .A(G2100), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G67), .A2(n640), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G80), .A2(n637), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n647), .A2(G55), .ZN(n617) );
  NAND2_X1 U703 ( .A1(G93), .A2(n588), .ZN(n616) );
  NAND2_X1 U704 ( .A1(n617), .A2(n616), .ZN(n618) );
  OR2_X1 U705 ( .A1(n619), .A2(n618), .ZN(n659) );
  NAND2_X1 U706 ( .A1(G559), .A2(n980), .ZN(n620) );
  XOR2_X1 U707 ( .A(n996), .B(n620), .Z(n656) );
  NAND2_X1 U708 ( .A1(n621), .A2(n656), .ZN(n622) );
  XNOR2_X1 U709 ( .A(n622), .B(KEYINPUT73), .ZN(n623) );
  XOR2_X1 U710 ( .A(n659), .B(n623), .Z(G145) );
  NAND2_X1 U711 ( .A1(G75), .A2(n637), .ZN(n625) );
  NAND2_X1 U712 ( .A1(G88), .A2(n588), .ZN(n624) );
  NAND2_X1 U713 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U714 ( .A1(G62), .A2(n640), .ZN(n627) );
  NAND2_X1 U715 ( .A1(G50), .A2(n647), .ZN(n626) );
  NAND2_X1 U716 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U717 ( .A1(n629), .A2(n628), .ZN(G166) );
  NAND2_X1 U718 ( .A1(G87), .A2(n630), .ZN(n631) );
  XNOR2_X1 U719 ( .A(n631), .B(KEYINPUT74), .ZN(n636) );
  NAND2_X1 U720 ( .A1(G49), .A2(n647), .ZN(n633) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U723 ( .A1(n640), .A2(n634), .ZN(n635) );
  NAND2_X1 U724 ( .A1(n636), .A2(n635), .ZN(G288) );
  XOR2_X1 U725 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n639) );
  NAND2_X1 U726 ( .A1(G73), .A2(n637), .ZN(n638) );
  XNOR2_X1 U727 ( .A(n639), .B(n638), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n640), .A2(G61), .ZN(n641) );
  XNOR2_X1 U729 ( .A(KEYINPUT75), .B(n641), .ZN(n642) );
  NOR2_X1 U730 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U731 ( .A1(G86), .A2(n588), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U733 ( .A(n646), .B(KEYINPUT77), .ZN(n649) );
  NAND2_X1 U734 ( .A1(G48), .A2(n647), .ZN(n648) );
  NAND2_X1 U735 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U736 ( .A(G166), .B(G288), .ZN(n655) );
  XNOR2_X1 U737 ( .A(KEYINPUT78), .B(KEYINPUT19), .ZN(n651) );
  XNOR2_X1 U738 ( .A(G305), .B(n708), .ZN(n650) );
  XNOR2_X1 U739 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U740 ( .A(n659), .B(n652), .Z(n653) );
  XNOR2_X1 U741 ( .A(n653), .B(G290), .ZN(n654) );
  XNOR2_X1 U742 ( .A(n655), .B(n654), .ZN(n909) );
  XOR2_X1 U743 ( .A(n909), .B(n656), .Z(n657) );
  NOR2_X1 U744 ( .A1(n658), .A2(n657), .ZN(n661) );
  NOR2_X1 U745 ( .A1(G868), .A2(n659), .ZN(n660) );
  NOR2_X1 U746 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G236), .A2(G238), .ZN(n666) );
  NAND2_X1 U754 ( .A1(G69), .A2(n666), .ZN(n667) );
  NOR2_X1 U755 ( .A1(G237), .A2(n667), .ZN(n834) );
  NOR2_X1 U756 ( .A1(n834), .A2(n668), .ZN(n675) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U759 ( .A1(G218), .A2(n670), .ZN(n671) );
  XOR2_X1 U760 ( .A(KEYINPUT79), .B(n671), .Z(n672) );
  NAND2_X1 U761 ( .A1(G96), .A2(n672), .ZN(n832) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n832), .ZN(n673) );
  XOR2_X1 U763 ( .A(KEYINPUT80), .B(n673), .Z(n674) );
  NOR2_X1 U764 ( .A1(n675), .A2(n674), .ZN(G319) );
  INV_X1 U765 ( .A(G319), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U767 ( .A1(n677), .A2(n676), .ZN(n831) );
  NAND2_X1 U768 ( .A1(n831), .A2(G36), .ZN(n678) );
  XOR2_X1 U769 ( .A(KEYINPUT81), .B(n678), .Z(G176) );
  XOR2_X1 U770 ( .A(KEYINPUT84), .B(G166), .Z(G303) );
  AND2_X1 U771 ( .A1(n679), .A2(G40), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U773 ( .A(KEYINPUT85), .B(n682), .Z(n797) );
  INV_X1 U774 ( .A(n797), .ZN(n683) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n798) );
  INV_X1 U776 ( .A(n728), .ZN(n702) );
  OR2_X1 U777 ( .A1(n702), .A2(G1961), .ZN(n685) );
  XNOR2_X1 U778 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NAND2_X1 U779 ( .A1(n702), .A2(n955), .ZN(n684) );
  NAND2_X1 U780 ( .A1(n685), .A2(n684), .ZN(n721) );
  NAND2_X1 U781 ( .A1(n721), .A2(G171), .ZN(n714) );
  NAND2_X1 U782 ( .A1(G2067), .A2(n702), .ZN(n687) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n728), .ZN(n686) );
  NAND2_X1 U784 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U785 ( .A(KEYINPUT91), .B(n688), .Z(n695) );
  INV_X1 U786 ( .A(G1996), .ZN(n949) );
  NOR2_X1 U787 ( .A1(n728), .A2(n949), .ZN(n689) );
  XNOR2_X1 U788 ( .A(n689), .B(KEYINPUT26), .ZN(n693) );
  NAND2_X1 U789 ( .A1(n728), .A2(G1341), .ZN(n690) );
  NAND2_X1 U790 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U791 ( .A1(n697), .A2(n980), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U793 ( .A(n696), .B(KEYINPUT92), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n980), .A2(n697), .ZN(n698) );
  XNOR2_X1 U795 ( .A(KEYINPUT93), .B(n698), .ZN(n699) );
  NAND2_X1 U796 ( .A1(n700), .A2(n699), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n702), .A2(G2072), .ZN(n701) );
  XNOR2_X1 U798 ( .A(n701), .B(KEYINPUT27), .ZN(n704) );
  INV_X1 U799 ( .A(G1956), .ZN(n1013) );
  NOR2_X1 U800 ( .A1(n1013), .A2(n702), .ZN(n703) );
  NOR2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n711) );
  NOR2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U805 ( .A(n709), .B(KEYINPUT28), .Z(n710) );
  NAND2_X1 U806 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U807 ( .A(KEYINPUT29), .B(n712), .Z(n713) );
  NAND2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n727) );
  INV_X1 U809 ( .A(KEYINPUT30), .ZN(n718) );
  NAND2_X1 U810 ( .A1(G8), .A2(n728), .ZN(n764) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n764), .ZN(n740) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n728), .ZN(n737) );
  INV_X1 U813 ( .A(n737), .ZN(n715) );
  NAND2_X1 U814 ( .A1(G8), .A2(n715), .ZN(n716) );
  NOR2_X1 U815 ( .A1(n740), .A2(n716), .ZN(n717) );
  XNOR2_X1 U816 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U817 ( .A1(n719), .A2(G168), .ZN(n720) );
  XNOR2_X1 U818 ( .A(n720), .B(KEYINPUT94), .ZN(n723) );
  NOR2_X1 U819 ( .A1(n721), .A2(G171), .ZN(n722) );
  NOR2_X1 U820 ( .A1(n723), .A2(n722), .ZN(n725) );
  NAND2_X1 U821 ( .A1(n727), .A2(n726), .ZN(n738) );
  NAND2_X1 U822 ( .A1(n738), .A2(G286), .ZN(n733) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n764), .ZN(n730) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n728), .ZN(n729) );
  NOR2_X1 U825 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U826 ( .A1(n731), .A2(G303), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n734), .A2(G8), .ZN(n736) );
  XOR2_X1 U829 ( .A(KEYINPUT95), .B(KEYINPUT32), .Z(n735) );
  XNOR2_X1 U830 ( .A(n736), .B(n735), .ZN(n744) );
  NAND2_X1 U831 ( .A1(G8), .A2(n737), .ZN(n742) );
  INV_X1 U832 ( .A(n738), .ZN(n739) );
  NOR2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n744), .A2(n743), .ZN(n763) );
  NOR2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U837 ( .A1(G303), .A2(G1971), .ZN(n745) );
  NOR2_X1 U838 ( .A1(n751), .A2(n745), .ZN(n990) );
  NAND2_X1 U839 ( .A1(n763), .A2(n990), .ZN(n746) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n989) );
  NAND2_X1 U841 ( .A1(n746), .A2(n989), .ZN(n747) );
  NAND2_X1 U842 ( .A1(n522), .A2(n748), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n752), .A2(n764), .ZN(n754) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n976) );
  INV_X1 U846 ( .A(KEYINPUT97), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n758), .B(n757), .ZN(n813) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U849 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  NOR2_X1 U850 ( .A1(n764), .A2(n760), .ZN(n768) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n761) );
  NAND2_X1 U852 ( .A1(G8), .A2(n761), .ZN(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U855 ( .A(n766), .B(KEYINPUT98), .Z(n767) );
  NOR2_X1 U856 ( .A1(n768), .A2(n767), .ZN(n811) );
  NAND2_X1 U857 ( .A1(G104), .A2(n888), .ZN(n770) );
  NAND2_X1 U858 ( .A1(G140), .A2(n889), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n771), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G116), .A2(n893), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G128), .A2(n894), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U864 ( .A(n774), .B(KEYINPUT35), .Z(n775) );
  NOR2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT36), .B(n777), .Z(n778) );
  XNOR2_X1 U867 ( .A(KEYINPUT86), .B(n778), .ZN(n906) );
  XOR2_X1 U868 ( .A(KEYINPUT37), .B(G2067), .Z(n805) );
  OR2_X1 U869 ( .A1(n906), .A2(n805), .ZN(n779) );
  XNOR2_X1 U870 ( .A(n779), .B(KEYINPUT100), .ZN(n940) );
  NAND2_X1 U871 ( .A1(n894), .A2(G129), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G117), .A2(n893), .ZN(n781) );
  NAND2_X1 U873 ( .A1(G141), .A2(n889), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n888), .A2(G105), .ZN(n782) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n782), .Z(n783) );
  NOR2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U879 ( .A(KEYINPUT89), .B(n787), .ZN(n903) );
  AND2_X1 U880 ( .A1(n949), .A2(n903), .ZN(n926) );
  NAND2_X1 U881 ( .A1(G95), .A2(n888), .ZN(n789) );
  NAND2_X1 U882 ( .A1(G131), .A2(n889), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U884 ( .A(KEYINPUT88), .B(n790), .Z(n794) );
  NAND2_X1 U885 ( .A1(G107), .A2(n893), .ZN(n792) );
  NAND2_X1 U886 ( .A1(G119), .A2(n894), .ZN(n791) );
  AND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n900) );
  AND2_X1 U889 ( .A1(n900), .A2(G1991), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n949), .A2(n903), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n928) );
  INV_X1 U892 ( .A(n928), .ZN(n799) );
  NOR2_X1 U893 ( .A1(n798), .A2(n797), .ZN(n818) );
  NAND2_X1 U894 ( .A1(n799), .A2(n818), .ZN(n815) );
  INV_X1 U895 ( .A(n815), .ZN(n802) );
  NOR2_X1 U896 ( .A1(G1991), .A2(n900), .ZN(n930) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U898 ( .A1(n930), .A2(n800), .ZN(n801) );
  NOR2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n926), .A2(n803), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n804), .B(KEYINPUT39), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n906), .A2(n805), .ZN(n806) );
  XNOR2_X1 U903 ( .A(n806), .B(KEYINPUT87), .ZN(n938) );
  NAND2_X1 U904 ( .A1(n818), .A2(n938), .ZN(n816) );
  NAND2_X1 U905 ( .A1(n807), .A2(n816), .ZN(n808) );
  XOR2_X1 U906 ( .A(KEYINPUT99), .B(n808), .Z(n809) );
  NAND2_X1 U907 ( .A1(n940), .A2(n809), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n810), .A2(n818), .ZN(n814) );
  AND2_X1 U909 ( .A1(n811), .A2(n814), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n824) );
  INV_X1 U911 ( .A(n814), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U913 ( .A(n817), .B(KEYINPUT90), .ZN(n820) );
  XNOR2_X1 U914 ( .A(G1986), .B(G290), .ZN(n986) );
  AND2_X1 U915 ( .A1(n986), .A2(n818), .ZN(n819) );
  NOR2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n821) );
  OR2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U919 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U920 ( .A(G223), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(G2106), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(KEYINPUT104), .ZN(G217) );
  NAND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n828) );
  XNOR2_X1 U924 ( .A(KEYINPUT105), .B(n828), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n829), .A2(G661), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U927 ( .A1(n831), .A2(n830), .ZN(G188) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  INV_X1 U930 ( .A(n832), .ZN(n833) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G261) );
  INV_X1 U932 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U933 ( .A(G2427), .B(G2443), .ZN(n844) );
  XOR2_X1 U934 ( .A(G2430), .B(KEYINPUT102), .Z(n836) );
  XNOR2_X1 U935 ( .A(G2454), .B(G2435), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U937 ( .A(G2438), .B(KEYINPUT101), .Z(n838) );
  XNOR2_X1 U938 ( .A(G1341), .B(G1348), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U940 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U941 ( .A(G2446), .B(G2451), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n845), .A2(G14), .ZN(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT103), .B(n846), .ZN(G401) );
  XOR2_X1 U946 ( .A(G2100), .B(G2096), .Z(n848) );
  XNOR2_X1 U947 ( .A(KEYINPUT42), .B(G2678), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(KEYINPUT43), .B(G2090), .Z(n850) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U955 ( .A(G2474), .B(G1976), .Z(n856) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1961), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U958 ( .A(n857), .B(KEYINPUT106), .Z(n859) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(G1971), .B(G1956), .Z(n861) );
  XNOR2_X1 U962 ( .A(G1981), .B(G1966), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(KEYINPUT41), .B(KEYINPUT107), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G112), .A2(n893), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G100), .A2(n888), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(KEYINPUT108), .B(n868), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n894), .A2(G124), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G136), .A2(n889), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(G162) );
  XOR2_X1 U976 ( .A(G162), .B(n931), .Z(n875) );
  XNOR2_X1 U977 ( .A(G164), .B(G160), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n875), .B(n874), .ZN(n887) );
  XOR2_X1 U979 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n885) );
  NAND2_X1 U980 ( .A1(G103), .A2(n888), .ZN(n877) );
  NAND2_X1 U981 ( .A1(G139), .A2(n889), .ZN(n876) );
  NAND2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G115), .A2(n893), .ZN(n879) );
  NAND2_X1 U984 ( .A1(G127), .A2(n894), .ZN(n878) );
  NAND2_X1 U985 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U986 ( .A(KEYINPUT111), .B(n880), .ZN(n881) );
  XNOR2_X1 U987 ( .A(KEYINPUT47), .B(n881), .ZN(n882) );
  NOR2_X1 U988 ( .A1(n883), .A2(n882), .ZN(n920) );
  XNOR2_X1 U989 ( .A(n920), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U990 ( .A(n885), .B(n884), .ZN(n886) );
  XOR2_X1 U991 ( .A(n887), .B(n886), .Z(n905) );
  NAND2_X1 U992 ( .A1(G106), .A2(n888), .ZN(n891) );
  NAND2_X1 U993 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n892), .B(KEYINPUT45), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G118), .A2(n893), .ZN(n896) );
  NAND2_X1 U997 ( .A1(G130), .A2(n894), .ZN(n895) );
  NAND2_X1 U998 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(KEYINPUT109), .B(n897), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n901) );
  XOR2_X1 U1001 ( .A(n901), .B(n900), .Z(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n908) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n908), .ZN(G395) );
  XOR2_X1 U1006 ( .A(n909), .B(G286), .Z(n911) );
  XNOR2_X1 U1007 ( .A(G171), .B(n980), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n912), .B(n996), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n913), .ZN(G397) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(KEYINPUT112), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n916), .ZN(n917) );
  AND2_X1 U1015 ( .A1(G319), .A2(n917), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1020 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(G2072), .B(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G164), .B(G2078), .ZN(n921) );
  NAND2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n924), .B(n923), .ZN(n944) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1027 ( .A(KEYINPUT51), .B(n927), .Z(n936) );
  XNOR2_X1 U1028 ( .A(G160), .B(G2084), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(KEYINPUT113), .B(n932), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(KEYINPUT114), .B(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1037 ( .A(KEYINPUT115), .B(n942), .Z(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1039 ( .A(KEYINPUT52), .B(n945), .Z(n946) );
  NOR2_X1 U1040 ( .A1(KEYINPUT55), .A2(n946), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT117), .B(n947), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(G29), .ZN(n975) );
  INV_X1 U1043 ( .A(G29), .ZN(n971) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n951) );
  XNOR2_X1 U1045 ( .A(n949), .B(G32), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G25), .B(G1991), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n960) );
  XOR2_X1 U1049 ( .A(G2072), .B(G33), .Z(n954) );
  NAND2_X1 U1050 ( .A1(n954), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G27), .B(n955), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT119), .B(n956), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT53), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G2084), .B(KEYINPUT54), .Z(n962) );
  XNOR2_X1 U1057 ( .A(G34), .B(n962), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT118), .B(G2090), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(G35), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT55), .B(n968), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(KEYINPUT120), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(G11), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n973), .B(KEYINPUT121), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n1031) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n978), .B(KEYINPUT122), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(KEYINPUT57), .B(n979), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(n980), .B(G1348), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G171), .B(G1961), .Z(n982) );
  XNOR2_X1 U1075 ( .A(G299), .B(G1956), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n995) );
  AND2_X1 U1080 ( .A1(G303), .A2(G1971), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(n993), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1085 ( .A(G1341), .B(n996), .Z(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1029) );
  INV_X1 U1088 ( .A(G16), .ZN(n1027) );
  XNOR2_X1 U1089 ( .A(G1986), .B(G24), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(G1976), .B(G23), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT127), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT58), .B(n1006), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G1966), .B(G21), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(G5), .B(G1961), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1024) );
  XOR2_X1 U1100 ( .A(G1348), .B(KEYINPUT59), .Z(n1011) );
  XNOR2_X1 U1101 ( .A(G4), .B(n1011), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(G1341), .B(G19), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(n1012), .B(KEYINPUT124), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(G1981), .B(G6), .Z(n1015) );
  XNOR2_X1 U1105 ( .A(n1013), .B(G20), .ZN(n1014) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(n1018), .B(KEYINPUT125), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1110 ( .A(KEYINPUT126), .B(n1021), .Z(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT60), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1117 ( .A(n1032), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

