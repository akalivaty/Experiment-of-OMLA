//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G58), .ZN(new_n207));
  INV_X1    g0007(.A(G232), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G77), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT65), .B(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n212), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  OAI21_X1  g0024(.A(G50), .B1(G58), .B2(G68), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n226), .A2(G20), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(G13), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n230), .B(G250), .C1(G257), .C2(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT0), .ZN(new_n232));
  NAND3_X1  g0032(.A1(new_n224), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(new_n203), .A2(G20), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  INV_X1    g0051(.A(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n253), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n250), .B1(new_n251), .B2(new_n254), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n227), .B1(new_n206), .B2(new_n253), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n267), .A2(new_n264), .A3(G13), .A4(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n202), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n259), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n264), .A2(G20), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n273), .B(KEYINPUT69), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(G50), .A3(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n263), .A2(KEYINPUT9), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n271), .B(new_n275), .C1(new_n261), .C2(new_n262), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G223), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G222), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n227), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n284), .B(new_n286), .C1(new_n214), .C2(new_n280), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G226), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n228), .B1(new_n253), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n288), .A2(KEYINPUT66), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT66), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n296), .B(new_n264), .C1(G41), .C2(G45), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n287), .B(new_n291), .C1(new_n292), .C2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g0101(.A(KEYINPUT75), .B(G200), .Z(new_n302));
  INV_X1    g0102(.A(KEYINPUT77), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n299), .A2(new_n302), .B1(new_n303), .B2(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n276), .A2(new_n279), .A3(new_n301), .A4(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n299), .A2(G179), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n277), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n291), .B1(new_n298), .B2(new_n208), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n292), .A2(G1698), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n280), .B(new_n314), .C1(G223), .C2(G1698), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G33), .A2(G87), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT84), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n294), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G179), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n308), .B2(new_n319), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n280), .B2(G20), .ZN(new_n323));
  AND2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n252), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n220), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n207), .A2(new_n220), .ZN(new_n329));
  OAI21_X1  g0129(.A(G20), .B1(new_n329), .B2(new_n201), .ZN(new_n330));
  INV_X1    g0130(.A(G159), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n254), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n328), .B1(KEYINPUT82), .B2(new_n332), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n332), .A2(KEYINPUT82), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(KEYINPUT16), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n328), .B2(new_n332), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n259), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT83), .ZN(new_n339));
  INV_X1    g0139(.A(new_n255), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n274), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n272), .A2(new_n341), .B1(new_n270), .B2(new_n255), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n339), .B1(new_n338), .B2(new_n342), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n321), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(KEYINPUT85), .A3(KEYINPUT18), .ZN(new_n346));
  OAI21_X1  g0146(.A(G200), .B1(new_n313), .B2(new_n318), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n338), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT87), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n319), .A2(G190), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT86), .B(KEYINPUT17), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n338), .A2(new_n350), .A3(new_n342), .A4(new_n347), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT17), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT87), .B1(new_n354), .B2(new_n351), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n338), .A2(new_n342), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT83), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g0161(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n362));
  NAND2_X1  g0162(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n361), .A2(new_n321), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n346), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n266), .A2(KEYINPUT74), .A3(new_n268), .ZN(new_n366));
  AOI21_X1  g0166(.A(KEYINPUT74), .B1(new_n266), .B2(new_n268), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n259), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n368), .A2(new_n274), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G77), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n213), .B1(new_n366), .B2(new_n367), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n255), .A2(new_n254), .B1(new_n213), .B2(new_n252), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n374), .B(KEYINPUT73), .ZN(new_n375));
  XOR2_X1   g0175(.A(KEYINPUT15), .B(G87), .Z(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n377), .A2(new_n257), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n259), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n372), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n294), .A2(new_n295), .A3(new_n215), .A4(new_n297), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n291), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT70), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n280), .A2(G232), .A3(new_n282), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT71), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n326), .A2(G107), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n280), .A2(KEYINPUT71), .A3(G232), .A4(new_n282), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n280), .A2(G238), .A3(G1698), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n387), .A2(new_n388), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n286), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT72), .B1(new_n384), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT70), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n383), .B(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT72), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(new_n392), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(new_n398), .A3(new_n302), .ZN(new_n399));
  INV_X1    g0199(.A(new_n398), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n396), .B2(new_n392), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n381), .B(new_n399), .C1(new_n402), .C2(new_n300), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n312), .A2(new_n365), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT12), .B(new_n220), .C1(new_n366), .C2(new_n367), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n256), .A2(G77), .B1(G20), .B2(new_n220), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT80), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n202), .B2(new_n254), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(new_n259), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n410), .A2(KEYINPUT11), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(KEYINPUT11), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n406), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n270), .A2(KEYINPUT12), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n220), .B1(new_n370), .B2(KEYINPUT12), .ZN(new_n415));
  NOR3_X1   g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n298), .A2(new_n221), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n290), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n292), .A2(G1698), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n324), .B2(new_n325), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT78), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT78), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n419), .B(new_n424), .C1(new_n325), .C2(new_n324), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n421), .A2(new_n422), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n426), .A2(new_n427), .A3(new_n286), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n426), .B2(new_n286), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n418), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT13), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT13), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n418), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G200), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n426), .A2(new_n286), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT79), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n426), .A2(new_n427), .A3(new_n286), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n432), .B1(new_n439), .B2(new_n418), .ZN(new_n440));
  INV_X1    g0240(.A(new_n433), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G190), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n416), .A2(new_n435), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n440), .B2(new_n441), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT14), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(G179), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT14), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n434), .A2(new_n449), .A3(G169), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT81), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT81), .A4(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n416), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n445), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n402), .A2(new_n308), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT76), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n394), .A2(new_n398), .ZN(new_n460));
  INV_X1    g0260(.A(G179), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI211_X1 g0262(.A(KEYINPUT76), .B(G179), .C1(new_n394), .C2(new_n398), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n458), .B(new_n380), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n405), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(G264), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT90), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT90), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n280), .A2(new_n468), .A3(G264), .A4(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n326), .A2(G303), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n280), .A2(G257), .A3(new_n282), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT88), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT5), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G41), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n293), .A2(KEYINPUT88), .A3(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n264), .A2(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n286), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n472), .A2(new_n286), .B1(G270), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n475), .A2(new_n476), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(KEYINPUT5), .B2(new_n293), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n483), .A2(new_n486), .A3(new_n289), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n482), .A2(G190), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT74), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n269), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n266), .A2(KEYINPUT74), .A3(new_n268), .ZN(new_n492));
  INV_X1    g0292(.A(G116), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n264), .B2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n369), .A4(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n366), .B2(new_n367), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  INV_X1    g0297(.A(G97), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n252), .C1(G33), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n493), .A2(G20), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n259), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT20), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n499), .A2(new_n259), .A3(KEYINPUT20), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n495), .A2(new_n496), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AOI221_X4 g0307(.A(new_n487), .B1(G270), .B2(new_n481), .C1(new_n472), .C2(new_n286), .ZN(new_n508));
  INV_X1    g0308(.A(G200), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n489), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT91), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(KEYINPUT21), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n506), .A2(G169), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n508), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n472), .A2(new_n286), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n481), .A2(G270), .ZN(new_n516));
  AND4_X1   g0316(.A1(G179), .A2(new_n515), .A3(new_n488), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n506), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n482), .A2(new_n488), .ZN(new_n519));
  INV_X1    g0319(.A(new_n512), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n519), .A2(G169), .A3(new_n506), .A4(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n510), .A2(new_n514), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n252), .B(G87), .C1(new_n324), .C2(new_n325), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n280), .A2(new_n526), .A3(new_n252), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n256), .A2(G116), .ZN(new_n529));
  INV_X1    g0329(.A(G107), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n530), .A2(KEYINPUT23), .A3(G20), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT23), .B1(new_n530), .B2(G20), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AND4_X1   g0334(.A1(new_n523), .A2(new_n528), .A3(new_n529), .A4(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n525), .B2(new_n527), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n523), .B1(new_n536), .B2(new_n529), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n259), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G264), .B(new_n294), .C1(new_n483), .C2(new_n486), .ZN(new_n539));
  OAI211_X1 g0339(.A(G250), .B(new_n282), .C1(new_n324), .C2(new_n325), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n324), .C2(new_n325), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G33), .A2(G294), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n286), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n488), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT25), .B1(new_n269), .B2(G107), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n264), .A2(G33), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n269), .A2(new_n369), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G107), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT25), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n270), .A2(new_n551), .A3(new_n530), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n538), .A2(new_n546), .A3(new_n547), .A4(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n545), .A2(new_n300), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n522), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n538), .A2(new_n547), .A3(new_n554), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n545), .A2(new_n308), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n545), .A2(G179), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n530), .B1(new_n323), .B2(new_n327), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n254), .A2(new_n371), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT6), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n498), .A2(new_n530), .ZN(new_n567));
  NOR2_X1   g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n530), .A2(KEYINPUT6), .A3(G97), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n252), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OR3_X1    g0371(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n259), .B1(new_n498), .B2(new_n270), .ZN(new_n573));
  OR2_X1    g0373(.A1(KEYINPUT3), .A2(G33), .ZN(new_n574));
  NAND2_X1  g0374(.A1(KEYINPUT3), .A2(G33), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n210), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  OAI21_X1  g0377(.A(G1698), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(G244), .B1(new_n324), .B2(new_n325), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(new_n577), .B1(G33), .B2(G283), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n577), .A2(G1698), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(G244), .C1(new_n325), .C2(new_n324), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n286), .B1(G257), .B2(new_n481), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(G190), .A3(new_n488), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n549), .A2(G97), .ZN(new_n586));
  INV_X1    g0386(.A(G244), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n574), .B2(new_n575), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n582), .B(new_n497), .C1(new_n588), .C2(KEYINPUT4), .ZN(new_n589));
  OAI21_X1  g0389(.A(G250), .B1(new_n324), .B2(new_n325), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n282), .B1(new_n590), .B2(KEYINPUT4), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n286), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n481), .A2(G257), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n488), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(G200), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n573), .A2(new_n585), .A3(new_n586), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n270), .A2(new_n498), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n597), .B(new_n586), .C1(new_n598), .C2(new_n369), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n584), .A2(new_n461), .A3(new_n488), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n594), .A2(new_n308), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n221), .A2(new_n282), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n587), .A2(G1698), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(new_n605), .C1(new_n324), .C2(new_n325), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G33), .A2(G116), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n294), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n479), .A2(new_n289), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n479), .B(G250), .C1(new_n285), .C2(new_n227), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G190), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT89), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(G20), .B1(new_n574), .B2(new_n575), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G68), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT19), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n257), .B2(new_n498), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n209), .A2(new_n498), .A3(new_n530), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n423), .A2(new_n252), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT19), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n259), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n269), .A2(new_n369), .A3(G87), .A4(new_n548), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n377), .B1(new_n366), .B2(new_n367), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n609), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n606), .A2(new_n607), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n610), .C1(new_n630), .C2(new_n294), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n302), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n612), .A2(KEYINPUT89), .A3(G190), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n615), .A2(new_n628), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n549), .A2(new_n376), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n624), .A3(new_n626), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n631), .A2(new_n308), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(G179), .C2(new_n631), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g0439(.A1(new_n563), .A2(new_n603), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n465), .A2(new_n558), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT92), .ZN(G372));
  AND3_X1   g0442(.A1(new_n514), .A2(new_n518), .A3(new_n521), .ZN(new_n643));
  INV_X1    g0443(.A(new_n302), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n612), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n627), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n643), .A2(new_n562), .B1(new_n646), .B2(new_n613), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n603), .A2(new_n557), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n639), .B2(new_n602), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT93), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n631), .A2(new_n651), .A3(new_n308), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n652), .A2(new_n636), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n637), .A2(KEYINPUT93), .B1(new_n461), .B2(new_n612), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n653), .A2(new_n654), .B1(new_n646), .B2(new_n613), .ZN(new_n655));
  INV_X1    g0455(.A(new_n602), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n654), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n650), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n649), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n465), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n311), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n416), .B1(new_n453), .B2(new_n454), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n445), .A2(new_n464), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n357), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n358), .A2(new_n321), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n670), .B2(new_n307), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n662), .A2(new_n671), .ZN(G369));
  INV_X1    g0472(.A(G13), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(G20), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n264), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n562), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n559), .A2(new_n680), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n556), .B2(new_n555), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n562), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n643), .A2(new_n680), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n681), .ZN(new_n687));
  INV_X1    g0487(.A(new_n643), .ZN(new_n688));
  INV_X1    g0488(.A(new_n680), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n507), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n522), .B2(new_n690), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(G330), .A3(new_n684), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(G399));
  NAND2_X1  g0494(.A1(new_n230), .A2(new_n293), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G1), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n620), .A2(G116), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n696), .A2(new_n697), .B1(new_n225), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n680), .B1(new_n649), .B2(new_n660), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n656), .A2(new_n657), .A3(new_n634), .A4(new_n638), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n655), .A2(new_n656), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n649), .A2(new_n659), .A3(new_n703), .A4(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n706), .A2(new_n689), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n702), .B1(new_n707), .B2(new_n701), .ZN(new_n708));
  INV_X1    g0508(.A(new_n560), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n526), .B1(new_n616), .B2(G87), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n529), .B(new_n534), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT24), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n536), .A2(new_n523), .A3(new_n529), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n553), .B1(new_n715), .B2(new_n259), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n709), .B1(new_n716), .B2(new_n547), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n639), .B1(new_n717), .B2(new_n561), .ZN(new_n718));
  INV_X1    g0518(.A(new_n603), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n558), .A2(new_n718), .A3(new_n719), .A4(new_n689), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT96), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n640), .A2(KEYINPUT96), .A3(new_n558), .A4(new_n689), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n488), .B1(new_n584), .B2(new_n482), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n461), .A3(new_n545), .A4(new_n631), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT95), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n726), .A2(new_n727), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n544), .A2(new_n539), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n482), .A3(G179), .A4(new_n488), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n592), .A2(new_n612), .A3(new_n488), .A4(new_n593), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND4_X1   g0534(.A1(new_n488), .A2(new_n592), .A3(new_n612), .A4(new_n593), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n517), .A2(new_n735), .A3(new_n728), .A4(new_n731), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n725), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  INV_X1    g0539(.A(new_n737), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(new_n689), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n722), .A2(new_n723), .A3(new_n738), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n708), .B1(G330), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n699), .B1(new_n743), .B2(G1), .ZN(G364));
  OR2_X1    g0544(.A1(new_n692), .A2(G330), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT97), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n692), .A2(G330), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n696), .B1(G45), .B2(new_n674), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n252), .A2(new_n300), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n461), .A2(new_n509), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n252), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G50), .A2(new_n754), .B1(new_n757), .B2(G68), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n461), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n751), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n755), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n758), .B1(new_n207), .B2(new_n760), .C1(new_n213), .C2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G179), .A2(G200), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n252), .B1(new_n763), .B2(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n498), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n762), .A2(new_n326), .A3(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n755), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n644), .A2(G179), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n755), .A2(new_n763), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(KEYINPUT32), .A3(G159), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT32), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n769), .B2(new_n331), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n768), .A2(G107), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n302), .A2(new_n461), .A3(new_n751), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n766), .B(new_n774), .C1(new_n209), .C2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT98), .ZN(new_n777));
  INV_X1    g0577(.A(G294), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n326), .B1(new_n764), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n757), .A2(new_n780), .B1(new_n770), .B2(G329), .ZN(new_n781));
  INV_X1    g0581(.A(new_n761), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G311), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n754), .A2(G326), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n779), .B(new_n785), .C1(G283), .C2(new_n768), .ZN(new_n786));
  INV_X1    g0586(.A(G303), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n775), .A2(KEYINPUT99), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n775), .A2(KEYINPUT99), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G322), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n786), .B1(new_n787), .B2(new_n790), .C1(new_n791), .C2(new_n760), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n777), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n227), .B1(G20), .B2(new_n308), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n749), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n326), .A2(new_n230), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n226), .A2(new_n484), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n797), .B(new_n798), .C1(new_n245), .C2(new_n484), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n280), .A2(G355), .A3(new_n230), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G116), .C2(new_n230), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n794), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n804), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n795), .B(new_n806), .C1(new_n692), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n750), .A2(new_n808), .ZN(G396));
  OAI21_X1  g0609(.A(KEYINPUT76), .B1(new_n402), .B2(G179), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n460), .A2(new_n459), .A3(new_n461), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n812), .A2(new_n458), .A3(new_n380), .A4(new_n689), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n380), .A2(new_n680), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n403), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n464), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(new_n700), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n700), .A2(new_n813), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n742), .A2(G330), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n821), .B(new_n822), .Z(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n749), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n817), .A2(new_n802), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G283), .A2(new_n757), .B1(new_n782), .B2(G116), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n778), .B2(new_n760), .C1(new_n787), .C2(new_n753), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G87), .B2(new_n768), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n280), .B(new_n765), .C1(G311), .C2(new_n770), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n530), .C2(new_n790), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n768), .A2(G68), .ZN(new_n831));
  INV_X1    g0631(.A(new_n760), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n832), .B1(new_n757), .B2(G150), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n834), .B2(new_n753), .C1(new_n331), .C2(new_n761), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT34), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n831), .B1(new_n207), .B2(new_n764), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n280), .B1(new_n769), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n835), .B2(new_n836), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n202), .B2(new_n790), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n830), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n794), .A2(new_n802), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n842), .A2(new_n794), .B1(new_n371), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n825), .A2(new_n748), .A3(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT100), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n824), .A2(new_n846), .ZN(G384));
  INV_X1    g0647(.A(KEYINPUT40), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n449), .B1(new_n434), .B2(G169), .ZN(new_n849));
  AOI211_X1 g0649(.A(KEYINPUT14), .B(new_n308), .C1(new_n431), .C2(new_n433), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(KEYINPUT81), .B1(new_n851), .B2(new_n448), .ZN(new_n852));
  INV_X1    g0652(.A(new_n454), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n456), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n689), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT102), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n416), .A2(new_n689), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n857), .B1(new_n457), .B2(new_n859), .ZN(new_n860));
  NOR4_X1   g0660(.A1(new_n664), .A2(KEYINPUT102), .A3(new_n445), .A4(new_n858), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n856), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n738), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n737), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n680), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n866), .A2(new_n722), .A3(new_n741), .A4(new_n723), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT106), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n862), .A2(new_n818), .A3(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n678), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n335), .A2(new_n259), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT16), .B1(new_n333), .B2(new_n334), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n342), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n365), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n345), .A2(new_n354), .ZN(new_n875));
  XOR2_X1   g0675(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n361), .B2(new_n870), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n873), .A2(new_n321), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n870), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n354), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n874), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n848), .B1(new_n869), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n854), .A2(new_n444), .A3(new_n859), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT102), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n457), .A2(new_n857), .A3(new_n859), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n855), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n817), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n870), .B1(new_n343), .B2(new_n344), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n354), .A3(new_n667), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n875), .A2(new_n877), .B1(new_n896), .B2(new_n876), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n895), .B1(new_n669), .B2(new_n357), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n892), .A2(KEYINPUT40), .A3(new_n900), .A4(new_n868), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n887), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n868), .A2(new_n465), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n902), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(G330), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n465), .A2(new_n708), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n671), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT104), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n906), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT39), .B1(new_n893), .B2(new_n899), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n886), .B2(KEYINPUT39), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n854), .A2(new_n680), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n669), .A2(new_n870), .ZN(new_n915));
  INV_X1    g0715(.A(new_n885), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n893), .ZN(new_n917));
  AND4_X1   g0717(.A1(new_n661), .A2(new_n689), .A3(new_n813), .A4(new_n816), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n464), .A2(new_n680), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT101), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT101), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n820), .A2(new_n921), .A3(new_n813), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n862), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n914), .A2(new_n915), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n910), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n264), .B2(new_n674), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n569), .A2(new_n570), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT35), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n252), .B(new_n227), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n930), .B(G116), .C1(new_n929), .C2(new_n928), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n213), .A2(new_n329), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n933), .A2(new_n225), .B1(G50), .B2(new_n220), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G1), .A3(new_n673), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n927), .A2(new_n932), .A3(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n599), .A2(new_n680), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n719), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n602), .B2(new_n689), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n686), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT42), .Z(new_n941));
  OAI21_X1  g0741(.A(new_n602), .B1(new_n938), .B2(new_n562), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n689), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n655), .B1(new_n628), .B2(new_n689), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n653), .A2(new_n654), .A3(new_n627), .A4(new_n680), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n941), .A2(new_n943), .B1(KEYINPUT43), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n947), .B(new_n948), .Z(new_n949));
  INV_X1    g0749(.A(KEYINPUT107), .ZN(new_n950));
  INV_X1    g0750(.A(new_n693), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n939), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n950), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n695), .B(KEYINPUT41), .Z(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n687), .A2(new_n939), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT44), .Z(new_n960));
  NAND2_X1  g0760(.A1(new_n687), .A2(new_n939), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT45), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n960), .A2(new_n951), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n951), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n684), .A2(new_n685), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n686), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT109), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n747), .B2(KEYINPUT108), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT109), .B1(new_n692), .B2(G330), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n967), .B2(new_n969), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n743), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n965), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n958), .B1(new_n975), .B2(new_n743), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n264), .B1(new_n674), .B2(G45), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n955), .B(new_n956), .C1(new_n976), .C2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n326), .B1(new_n764), .B2(new_n530), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n754), .A2(G311), .B1(new_n770), .B2(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n778), .B2(new_n756), .C1(new_n787), .C2(new_n760), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(G97), .C2(new_n768), .ZN(new_n983));
  INV_X1    g0783(.A(G283), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  INV_X1    g0785(.A(new_n790), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n985), .B1(new_n986), .B2(G116), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n775), .A2(KEYINPUT46), .A3(new_n493), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n983), .B1(new_n984), .B2(new_n761), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G150), .A2(new_n832), .B1(new_n782), .B2(G50), .ZN(new_n990));
  INV_X1    g0790(.A(G143), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n834), .B2(new_n769), .C1(new_n991), .C2(new_n753), .ZN(new_n992));
  AOI211_X1 g0792(.A(new_n326), .B(new_n992), .C1(G159), .C2(new_n757), .ZN(new_n993));
  INV_X1    g0793(.A(new_n764), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(G68), .ZN(new_n995));
  INV_X1    g0795(.A(new_n775), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(G58), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n768), .A2(new_n214), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n993), .A2(new_n995), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n989), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n749), .B1(new_n1001), .B2(new_n794), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n805), .B1(new_n230), .B2(new_n377), .C1(new_n241), .C2(new_n796), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n807), .C2(new_n946), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n979), .A2(new_n1004), .ZN(G387));
  NAND2_X1  g0805(.A1(new_n973), .A2(new_n978), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT110), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G311), .A2(new_n757), .B1(new_n832), .B2(G317), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n787), .B2(new_n761), .C1(new_n791), .C2(new_n753), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT48), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n984), .B2(new_n764), .C1(new_n778), .C2(new_n775), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT49), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n770), .A2(G326), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n280), .B1(new_n768), .B2(G116), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n775), .A2(new_n213), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n377), .A2(new_n764), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n280), .B1(new_n760), .B2(new_n202), .C1(new_n331), .C2(new_n753), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(G150), .C2(new_n770), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT112), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n756), .A2(new_n255), .B1(new_n761), .B2(new_n220), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n768), .A2(G97), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n1023), .A2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1017), .B1(new_n1018), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n794), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n340), .A2(new_n202), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n697), .B1(new_n1029), .B2(KEYINPUT50), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(G68), .A2(G77), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n484), .A4(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n797), .B(new_n1033), .C1(new_n238), .C2(new_n484), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n697), .A2(new_n230), .A3(new_n280), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(G107), .C2(new_n230), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT111), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n749), .B1(new_n1037), .B2(new_n805), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1028), .B(new_n1038), .C1(new_n684), .C2(new_n807), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n695), .B(KEYINPUT113), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n973), .B(new_n743), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1007), .B(new_n1039), .C1(new_n1040), .C2(new_n1041), .ZN(G393));
  XNOR2_X1  g0842(.A(new_n965), .B(KEYINPUT114), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n978), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n753), .A2(new_n251), .B1(new_n760), .B2(new_n331), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT115), .Z(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT51), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n768), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1048), .A2(new_n209), .B1(new_n220), .B2(new_n775), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n756), .A2(new_n202), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n326), .B1(new_n782), .B2(new_n340), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n994), .A2(G77), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n991), .C2(new_n769), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT116), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n756), .A2(new_n787), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G317), .A2(new_n754), .B1(new_n832), .B2(G311), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n326), .B1(new_n769), .B2(new_n791), .C1(new_n778), .C2(new_n761), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G116), .B2(new_n994), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n768), .A2(G107), .B1(new_n996), .B2(G283), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1055), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n749), .B1(new_n1063), .B2(new_n794), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n805), .B1(new_n498), .B2(new_n230), .C1(new_n248), .C2(new_n796), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n939), .A2(new_n807), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1044), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1040), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n965), .A2(new_n974), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n975), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1071), .ZN(G390));
  AOI21_X1  g0872(.A(new_n913), .B1(new_n893), .B2(new_n899), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n919), .B1(new_n707), .B2(new_n816), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1073), .B1(new_n891), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(G330), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n817), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n742), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n862), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n913), .B1(new_n862), .B2(new_n923), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1075), .B(new_n1080), .C1(new_n1081), .C2(new_n912), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(KEYINPUT117), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n913), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n921), .B1(new_n820), .B2(new_n813), .ZN(new_n1085));
  AOI211_X1 g0885(.A(KEYINPUT101), .B(new_n919), .C1(new_n700), .C2(new_n816), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n891), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT39), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n900), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n917), .B2(new_n1089), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT117), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1092), .A2(new_n1093), .A3(new_n1075), .A4(new_n1080), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1075), .B1(new_n1081), .B2(new_n912), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n867), .A2(KEYINPUT106), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n867), .A2(KEYINPUT106), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1077), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n891), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1096), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n671), .B(new_n907), .C1(new_n903), .C2(new_n1076), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n856), .B(new_n1078), .C1(new_n860), .C2(new_n861), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n891), .B2(new_n1099), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n923), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n891), .A2(new_n1099), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n1080), .A3(new_n1074), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1103), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1040), .B1(new_n1102), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1095), .A2(KEYINPUT118), .A3(new_n1101), .A4(new_n1109), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1083), .A2(new_n1109), .A3(new_n1094), .A4(new_n1101), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT118), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1095), .A2(new_n978), .A3(new_n1101), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n326), .B1(new_n769), .B2(new_n778), .C1(new_n493), .C2(new_n760), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n756), .A2(new_n530), .B1(new_n761), .B2(new_n498), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT119), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(G283), .C2(new_n754), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n986), .A2(G87), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1122), .A2(new_n831), .A3(new_n1052), .A4(new_n1123), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT54), .B(G143), .Z(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1126), .A2(new_n761), .B1(new_n1127), .B2(new_n769), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G128), .B2(new_n754), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n838), .B2(new_n760), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n326), .B(new_n1130), .C1(G159), .C2(new_n994), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n775), .A2(new_n251), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n202), .C2(new_n1048), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n756), .A2(new_n834), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1124), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1136), .A2(new_n794), .B1(new_n255), .B2(new_n843), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n748), .B(new_n1137), .C1(new_n912), .C2(new_n803), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1117), .A2(new_n1118), .A3(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1103), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n914), .A2(new_n915), .A3(new_n924), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n902), .B2(new_n1076), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n312), .B(KEYINPUT55), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n277), .A2(new_n870), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT56), .Z(new_n1146));
  XNOR2_X1  g0946(.A(new_n1144), .B(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n925), .A2(G330), .A3(new_n887), .A4(new_n901), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1143), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1140), .B1(new_n1141), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1147), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1143), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1113), .B(KEYINPUT118), .ZN(new_n1158));
  OAI211_X1 g0958(.A(KEYINPUT57), .B(new_n1157), .C1(new_n1158), .C2(new_n1103), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1152), .A2(new_n1159), .A3(new_n1069), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n753), .A2(new_n1127), .B1(new_n764), .B2(new_n251), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT120), .Z(new_n1162));
  NAND2_X1  g0962(.A1(new_n832), .A2(G128), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n756), .A2(new_n838), .B1(new_n761), .B2(new_n834), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n996), .B2(new_n1125), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1162), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT59), .Z(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n768), .B2(G159), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G33), .B1(new_n770), .B2(G124), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n202), .B1(new_n324), .B2(G41), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G116), .A2(new_n754), .B1(new_n832), .B2(G107), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n984), .B2(new_n769), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G97), .B2(new_n757), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n768), .A2(G58), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n326), .B1(new_n377), .B2(new_n761), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1018), .A2(new_n1176), .A3(G41), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n995), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT58), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1170), .A2(new_n1171), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n749), .B1(new_n1180), .B2(new_n794), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1154), .B2(new_n803), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n202), .B2(new_n843), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1157), .B2(new_n978), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1160), .A2(new_n1184), .ZN(G375));
  OAI21_X1  g0985(.A(new_n280), .B1(new_n764), .B2(new_n202), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G150), .A2(new_n782), .B1(new_n770), .B2(G128), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n838), .B2(new_n753), .C1(new_n834), .C2(new_n760), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G58), .C2(new_n768), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n331), .B2(new_n790), .C1(new_n756), .C2(new_n1126), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n790), .A2(new_n498), .B1(new_n787), .B2(new_n769), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1191), .B(KEYINPUT122), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G294), .A2(new_n754), .B1(new_n832), .B2(G283), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n530), .B2(new_n761), .ZN(new_n1194));
  OR3_X1    g0994(.A1(new_n1192), .A2(new_n1019), .A3(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n326), .B1(new_n493), .B2(new_n756), .C1(new_n1048), .C2(new_n371), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1190), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT123), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n749), .B1(new_n1198), .B2(new_n794), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n862), .B2(new_n803), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n220), .B2(new_n843), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n977), .B(KEYINPUT121), .Z(new_n1203));
  AOI21_X1  g1003(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1106), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n957), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1206), .B2(new_n1109), .ZN(G381));
  NOR2_X1   g1007(.A1(G375), .A2(G378), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1068), .A2(new_n979), .A3(new_n1004), .A4(new_n1071), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(G381), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1208), .A2(new_n1210), .A3(new_n1211), .ZN(G407));
  INV_X1    g1012(.A(G213), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1208), .B2(new_n679), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(G407), .ZN(G409));
  INV_X1    g1015(.A(G378), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n957), .B1(new_n1158), .B2(new_n1103), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1203), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1151), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1216), .B1(new_n1219), .B2(new_n1183), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1160), .A2(G378), .A3(new_n1184), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1213), .A2(G343), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT60), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1109), .B1(new_n1226), .B2(new_n1205), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1227), .B(new_n1069), .C1(new_n1226), .C2(new_n1205), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n1228), .A2(G384), .A3(new_n1204), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G384), .B1(new_n1228), .B2(new_n1204), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1223), .A2(G2897), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT125), .Z(new_n1233));
  XNOR2_X1  g1033(.A(new_n1231), .B(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT61), .B1(new_n1225), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1222), .A2(new_n1224), .A3(new_n1231), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT62), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1223), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1231), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1236), .A2(new_n1238), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G390), .A2(G387), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G393), .B(G396), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1243), .A2(new_n1209), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1243), .B2(new_n1209), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1247), .B(new_n1250), .C1(new_n1239), .C2(new_n1234), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1231), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1223), .B(new_n1254), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1253), .B1(new_n1255), .B2(KEYINPUT63), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1237), .A2(KEYINPUT124), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(KEYINPUT63), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1252), .A2(new_n1256), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1249), .A2(new_n1260), .ZN(G405));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1221), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(G378), .B1(new_n1160), .B2(new_n1184), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1254), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1265), .A2(new_n1254), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1264), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G375), .A2(new_n1216), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1231), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1247), .B(KEYINPUT127), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1248), .A2(KEYINPUT127), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n1273), .ZN(G402));
endmodule


