

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761;

  NOR2_X1 U371 ( .A1(n398), .A2(n397), .ZN(n427) );
  NOR2_X1 U372 ( .A1(n655), .A2(n654), .ZN(n580) );
  INV_X1 U373 ( .A(n605), .ZN(n650) );
  AND2_X2 U374 ( .A1(n597), .A2(n598), .ZN(n610) );
  NAND2_X2 U375 ( .A1(n605), .A2(n604), .ZN(n617) );
  XNOR2_X2 U376 ( .A(n387), .B(n359), .ZN(n757) );
  XNOR2_X2 U377 ( .A(n453), .B(G122), .ZN(n518) );
  XNOR2_X2 U378 ( .A(G107), .B(G116), .ZN(n453) );
  XNOR2_X2 U379 ( .A(n536), .B(n535), .ZN(n577) );
  XNOR2_X2 U380 ( .A(n505), .B(n542), .ZN(n731) );
  XNOR2_X2 U381 ( .A(n464), .B(n350), .ZN(n605) );
  NAND2_X1 U382 ( .A1(n610), .A2(n642), .ZN(n599) );
  AND2_X1 U383 ( .A1(n470), .A2(n472), .ZN(n463) );
  XNOR2_X1 U384 ( .A(n426), .B(n480), .ZN(n475) );
  XOR2_X2 U385 ( .A(KEYINPUT6), .B(n658), .Z(n616) );
  INV_X2 U386 ( .A(n606), .ZN(n658) );
  XNOR2_X1 U387 ( .A(n386), .B(n461), .ZN(n756) );
  OR2_X1 U388 ( .A1(n644), .A2(n414), .ZN(n413) );
  XNOR2_X1 U389 ( .A(n500), .B(n499), .ZN(n609) );
  XNOR2_X1 U390 ( .A(G119), .B(KEYINPUT67), .ZN(n431) );
  XNOR2_X1 U391 ( .A(n436), .B(n503), .ZN(n711) );
  XNOR2_X2 U392 ( .A(n440), .B(n504), .ZN(n542) );
  XNOR2_X2 U393 ( .A(n631), .B(KEYINPUT38), .ZN(n642) );
  NAND2_X1 U394 ( .A1(G237), .A2(G234), .ZN(n512) );
  XNOR2_X1 U395 ( .A(n459), .B(n519), .ZN(n559) );
  XOR2_X1 U396 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n519) );
  XNOR2_X1 U397 ( .A(G902), .B(KEYINPUT15), .ZN(n679) );
  XNOR2_X1 U398 ( .A(n479), .B(G125), .ZN(n373) );
  XNOR2_X1 U399 ( .A(n534), .B(n533), .ZN(n535) );
  NOR2_X1 U400 ( .A1(n721), .A2(G902), .ZN(n536) );
  INV_X1 U401 ( .A(KEYINPUT13), .ZN(n533) );
  XNOR2_X1 U402 ( .A(n603), .B(n388), .ZN(n563) );
  INV_X1 U403 ( .A(KEYINPUT94), .ZN(n388) );
  NAND2_X1 U404 ( .A1(n723), .A2(G478), .ZN(n407) );
  INV_X1 U405 ( .A(KEYINPUT47), .ZN(n384) );
  XOR2_X1 U406 ( .A(G140), .B(G131), .Z(n523) );
  XNOR2_X1 U407 ( .A(G122), .B(G113), .ZN(n522) );
  XNOR2_X1 U408 ( .A(n451), .B(n450), .ZN(n585) );
  INV_X1 U409 ( .A(KEYINPUT101), .ZN(n450) );
  NOR2_X1 U410 ( .A1(n584), .A2(n646), .ZN(n451) );
  XNOR2_X1 U411 ( .A(n431), .B(KEYINPUT3), .ZN(n440) );
  XOR2_X1 U412 ( .A(KEYINPUT88), .B(KEYINPUT76), .Z(n506) );
  XOR2_X1 U413 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n501) );
  XNOR2_X1 U414 ( .A(n543), .B(n494), .ZN(n503) );
  XNOR2_X1 U415 ( .A(n729), .B(KEYINPUT69), .ZN(n494) );
  XNOR2_X1 U416 ( .A(n564), .B(n361), .ZN(n433) );
  XNOR2_X1 U417 ( .A(n518), .B(KEYINPUT16), .ZN(n505) );
  XNOR2_X1 U418 ( .A(n429), .B(n520), .ZN(n724) );
  XNOR2_X1 U419 ( .A(n517), .B(n430), .ZN(n429) );
  XNOR2_X1 U420 ( .A(n485), .B(n484), .ZN(n721) );
  NOR2_X1 U421 ( .A1(n609), .A2(n608), .ZN(n614) );
  NAND2_X1 U422 ( .A1(n411), .A2(n408), .ZN(n640) );
  AND2_X1 U423 ( .A1(n415), .A2(n412), .ZN(n411) );
  NOR2_X1 U424 ( .A1(n421), .A2(n609), .ZN(n597) );
  XNOR2_X1 U425 ( .A(n589), .B(n588), .ZN(n598) );
  NAND2_X1 U426 ( .A1(n650), .A2(n422), .ZN(n421) );
  NAND2_X1 U427 ( .A1(n650), .A2(n563), .ZN(n654) );
  INV_X1 U428 ( .A(KEYINPUT0), .ZN(n435) );
  XNOR2_X1 U429 ( .A(n482), .B(n481), .ZN(n586) );
  INV_X1 U430 ( .A(KEYINPUT100), .ZN(n481) );
  INV_X1 U431 ( .A(n724), .ZN(n406) );
  INV_X1 U432 ( .A(n684), .ZN(n491) );
  AND2_X1 U433 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U434 ( .A1(n376), .A2(n375), .ZN(n374) );
  AND2_X1 U435 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U436 ( .A(n688), .ZN(n492) );
  XNOR2_X1 U437 ( .A(G116), .B(G137), .ZN(n544) );
  NAND2_X1 U438 ( .A1(n710), .A2(n709), .ZN(n473) );
  NOR2_X1 U439 ( .A1(n633), .A2(n474), .ZN(n471) );
  INV_X1 U440 ( .A(G953), .ZN(n510) );
  XNOR2_X1 U441 ( .A(n418), .B(G140), .ZN(n555) );
  INV_X1 U442 ( .A(G137), .ZN(n418) );
  XNOR2_X1 U443 ( .A(G134), .B(KEYINPUT7), .ZN(n516) );
  INV_X1 U444 ( .A(G104), .ZN(n524) );
  XNOR2_X1 U445 ( .A(n373), .B(KEYINPUT10), .ZN(n554) );
  XNOR2_X1 U446 ( .A(n555), .B(n417), .ZN(n496) );
  INV_X1 U447 ( .A(G107), .ZN(n417) );
  NAND2_X1 U448 ( .A1(n641), .A2(n601), .ZN(n410) );
  NAND2_X1 U449 ( .A1(n413), .A2(KEYINPUT41), .ZN(n412) );
  INV_X1 U450 ( .A(n641), .ZN(n414) );
  NAND2_X1 U451 ( .A1(n416), .A2(KEYINPUT41), .ZN(n415) );
  NAND2_X1 U452 ( .A1(G214), .A2(n508), .ZN(n641) );
  OR2_X1 U453 ( .A1(G902), .A2(G237), .ZN(n508) );
  AND2_X1 U454 ( .A1(n563), .A2(n595), .ZN(n422) );
  XNOR2_X1 U455 ( .A(n587), .B(KEYINPUT106), .ZN(n588) );
  NOR2_X1 U456 ( .A1(n734), .A2(G953), .ZN(n735) );
  XNOR2_X1 U457 ( .A(n425), .B(KEYINPUT92), .ZN(n424) );
  XNOR2_X1 U458 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n425) );
  XNOR2_X1 U459 ( .A(G128), .B(G119), .ZN(n423) );
  XNOR2_X1 U460 ( .A(n554), .B(n555), .ZN(n746) );
  XNOR2_X1 U461 ( .A(G110), .B(KEYINPUT68), .ZN(n556) );
  INV_X1 U462 ( .A(n679), .ZN(n683) );
  AND2_X1 U463 ( .A1(n681), .A2(KEYINPUT81), .ZN(n490) );
  AND2_X1 U464 ( .A1(n681), .A2(n468), .ZN(n684) );
  NOR2_X1 U465 ( .A1(n637), .A2(n349), .ZN(n468) );
  XNOR2_X1 U466 ( .A(n731), .B(n487), .ZN(n436) );
  NAND2_X1 U467 ( .A1(n684), .A2(n443), .ZN(n371) );
  INV_X1 U468 ( .A(n611), .ZN(n631) );
  XNOR2_X1 U469 ( .A(n540), .B(KEYINPUT22), .ZN(n572) );
  XNOR2_X1 U470 ( .A(n609), .B(KEYINPUT1), .ZN(n655) );
  NOR2_X1 U471 ( .A1(n724), .A2(G902), .ZN(n521) );
  NOR2_X1 U472 ( .A1(n726), .A2(G902), .ZN(n464) );
  INV_X1 U473 ( .A(KEYINPUT64), .ZN(n460) );
  XNOR2_X1 U474 ( .A(n561), .B(n465), .ZN(n726) );
  XNOR2_X1 U475 ( .A(n452), .B(n560), .ZN(n465) );
  XNOR2_X1 U476 ( .A(n746), .B(n558), .ZN(n561) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n560) );
  XNOR2_X1 U478 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n461) );
  NAND2_X1 U479 ( .A1(n640), .A2(n614), .ZN(n386) );
  NAND2_X1 U480 ( .A1(n632), .A2(n689), .ZN(n387) );
  XNOR2_X1 U481 ( .A(n568), .B(KEYINPUT35), .ZN(n759) );
  XNOR2_X1 U482 ( .A(n402), .B(n360), .ZN(n567) );
  INV_X1 U483 ( .A(n661), .ZN(n434) );
  NOR2_X1 U484 ( .A1(n583), .A2(n658), .ZN(n467) );
  NOR2_X1 U485 ( .A1(n654), .A2(n609), .ZN(n596) );
  XNOR2_X1 U486 ( .A(n743), .B(n456), .ZN(G69) );
  XNOR2_X1 U487 ( .A(n744), .B(n457), .ZN(n456) );
  INV_X1 U488 ( .A(KEYINPUT122), .ZN(n457) );
  INV_X1 U489 ( .A(KEYINPUT118), .ZN(n403) );
  INV_X1 U490 ( .A(KEYINPUT60), .ZN(n446) );
  INV_X1 U491 ( .A(KEYINPUT56), .ZN(n438) );
  INV_X1 U492 ( .A(G110), .ZN(n432) );
  AND2_X1 U493 ( .A1(n368), .A2(n358), .ZN(n347) );
  AND2_X1 U494 ( .A1(n374), .A2(KEYINPUT72), .ZN(n348) );
  INV_X1 U495 ( .A(G146), .ZN(n479) );
  XNOR2_X1 U496 ( .A(KEYINPUT78), .B(n638), .ZN(n349) );
  XOR2_X1 U497 ( .A(n553), .B(n552), .Z(n350) );
  XOR2_X1 U498 ( .A(n550), .B(G472), .Z(n351) );
  OR2_X1 U499 ( .A1(n648), .A2(n647), .ZN(n352) );
  AND2_X2 U500 ( .A1(n390), .A2(n491), .ZN(n723) );
  AND2_X1 U501 ( .A1(n710), .A2(n471), .ZN(n353) );
  NOR2_X1 U502 ( .A1(n684), .A2(n443), .ZN(n354) );
  OR2_X1 U503 ( .A1(n478), .A2(n477), .ZN(n355) );
  AND2_X1 U504 ( .A1(G210), .A2(n508), .ZN(n356) );
  AND2_X1 U505 ( .A1(n675), .A2(n674), .ZN(n357) );
  AND2_X1 U506 ( .A1(n357), .A2(n371), .ZN(n358) );
  XOR2_X1 U507 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n359) );
  XOR2_X1 U508 ( .A(KEYINPUT70), .B(KEYINPUT34), .Z(n360) );
  XNOR2_X1 U509 ( .A(KEYINPUT102), .B(KEYINPUT33), .ZN(n361) );
  INV_X1 U510 ( .A(KEYINPUT72), .ZN(n477) );
  XOR2_X1 U511 ( .A(n685), .B(KEYINPUT62), .Z(n362) );
  XOR2_X1 U512 ( .A(n713), .B(n712), .Z(n363) );
  XOR2_X1 U513 ( .A(n721), .B(n720), .Z(n364) );
  XNOR2_X1 U514 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n365) );
  NAND2_X1 U515 ( .A1(n683), .A2(KEYINPUT2), .ZN(n366) );
  INV_X1 U516 ( .A(KEYINPUT83), .ZN(n474) );
  INV_X1 U517 ( .A(KEYINPUT44), .ZN(n576) );
  NOR2_X1 U518 ( .A1(n752), .A2(G952), .ZN(n728) );
  INV_X1 U519 ( .A(n728), .ZN(n441) );
  XOR2_X1 U520 ( .A(KEYINPUT63), .B(KEYINPUT85), .Z(n367) );
  NOR2_X1 U521 ( .A1(n572), .A2(n621), .ZN(n570) );
  NAND2_X1 U522 ( .A1(n347), .A2(n370), .ZN(n372) );
  NAND2_X1 U523 ( .A1(n369), .A2(n354), .ZN(n368) );
  INV_X1 U524 ( .A(n639), .ZN(n369) );
  NAND2_X1 U525 ( .A1(n639), .A2(n443), .ZN(n370) );
  XNOR2_X1 U526 ( .A(n372), .B(n678), .ZN(G75) );
  XNOR2_X1 U527 ( .A(n373), .B(n506), .ZN(n507) );
  NAND2_X1 U528 ( .A1(n377), .A2(n374), .ZN(n383) );
  NAND2_X1 U529 ( .A1(n348), .A2(n377), .ZN(n380) );
  NOR2_X1 U530 ( .A1(n646), .A2(n384), .ZN(n375) );
  INV_X1 U531 ( .A(n695), .ZN(n376) );
  NAND2_X1 U532 ( .A1(n646), .A2(n384), .ZN(n378) );
  NAND2_X1 U533 ( .A1(n695), .A2(n384), .ZN(n379) );
  NAND2_X1 U534 ( .A1(n381), .A2(n380), .ZN(n398) );
  NAND2_X1 U535 ( .A1(n383), .A2(n382), .ZN(n381) );
  NOR2_X1 U536 ( .A1(n699), .A2(KEYINPUT72), .ZN(n382) );
  XNOR2_X2 U537 ( .A(n385), .B(G146), .ZN(n545) );
  XNOR2_X1 U538 ( .A(n747), .B(n385), .ZN(n751) );
  XNOR2_X2 U539 ( .A(G134), .B(G131), .ZN(n385) );
  NAND2_X1 U540 ( .A1(n757), .A2(n756), .ZN(n419) );
  XNOR2_X2 U541 ( .A(n599), .B(KEYINPUT39), .ZN(n632) );
  INV_X1 U542 ( .A(n603), .ZN(n651) );
  XNOR2_X2 U543 ( .A(n389), .B(n351), .ZN(n606) );
  OR2_X2 U544 ( .A1(n685), .A2(G902), .ZN(n389) );
  XNOR2_X1 U545 ( .A(n454), .B(n548), .ZN(n685) );
  NAND2_X1 U546 ( .A1(n391), .A2(n366), .ZN(n390) );
  NAND2_X1 U547 ( .A1(n393), .A2(n392), .ZN(n391) );
  NAND2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n392) );
  NAND2_X1 U549 ( .A1(n490), .A2(n682), .ZN(n393) );
  XNOR2_X2 U550 ( .A(n394), .B(KEYINPUT45), .ZN(n681) );
  NAND2_X1 U551 ( .A1(n395), .A2(n400), .ZN(n394) );
  XNOR2_X1 U552 ( .A(n396), .B(n576), .ZN(n395) );
  NAND2_X1 U553 ( .A1(n401), .A2(n760), .ZN(n396) );
  NAND2_X1 U554 ( .A1(n708), .A2(n355), .ZN(n397) );
  NAND2_X1 U555 ( .A1(n433), .A2(n399), .ZN(n402) );
  NAND2_X1 U556 ( .A1(n399), .A2(n539), .ZN(n540) );
  AND2_X1 U557 ( .A1(n434), .A2(n399), .ZN(n582) );
  NAND2_X1 U558 ( .A1(n399), .A2(n596), .ZN(n583) );
  XNOR2_X2 U559 ( .A(n466), .B(n435), .ZN(n399) );
  NOR2_X1 U560 ( .A1(n585), .A2(n492), .ZN(n400) );
  NOR2_X1 U561 ( .A1(n571), .A2(n759), .ZN(n401) );
  XNOR2_X1 U562 ( .A(n404), .B(n403), .ZN(G63) );
  NAND2_X1 U563 ( .A1(n405), .A2(n441), .ZN(n404) );
  XNOR2_X1 U564 ( .A(n407), .B(n406), .ZN(n405) );
  NAND2_X1 U565 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U566 ( .A1(n642), .A2(n409), .ZN(n408) );
  NOR2_X1 U567 ( .A1(n644), .A2(n410), .ZN(n409) );
  INV_X1 U568 ( .A(n642), .ZN(n416) );
  AND2_X1 U569 ( .A1(n352), .A2(n433), .ZN(n649) );
  NAND2_X1 U570 ( .A1(n664), .A2(n433), .ZN(n675) );
  XNOR2_X1 U571 ( .A(n419), .B(n365), .ZN(n428) );
  XNOR2_X1 U572 ( .A(n420), .B(KEYINPUT74), .ZN(n680) );
  XNOR2_X1 U573 ( .A(n420), .B(n751), .ZN(n753) );
  NOR2_X1 U574 ( .A1(n734), .A2(n420), .ZN(n634) );
  NAND2_X2 U575 ( .A1(n463), .A2(n462), .ZN(n420) );
  NAND2_X1 U576 ( .A1(n428), .A2(n427), .ZN(n426) );
  XNOR2_X1 U577 ( .A(n518), .B(n516), .ZN(n430) );
  XNOR2_X1 U578 ( .A(n571), .B(n432), .ZN(G12) );
  XNOR2_X1 U579 ( .A(n718), .B(n719), .ZN(n445) );
  INV_X2 U580 ( .A(n437), .ZN(n515) );
  XNOR2_X2 U581 ( .A(G143), .B(G128), .ZN(n437) );
  XNOR2_X1 U582 ( .A(n439), .B(n438), .ZN(G51) );
  NAND2_X1 U583 ( .A1(n442), .A2(n441), .ZN(n439) );
  XNOR2_X1 U584 ( .A(n547), .B(n549), .ZN(n454) );
  XNOR2_X1 U585 ( .A(n714), .B(n363), .ZN(n442) );
  XNOR2_X2 U586 ( .A(n575), .B(KEYINPUT32), .ZN(n760) );
  XNOR2_X1 U587 ( .A(n469), .B(KEYINPUT19), .ZN(n615) );
  INV_X1 U588 ( .A(KEYINPUT82), .ZN(n443) );
  XNOR2_X1 U589 ( .A(n444), .B(n367), .ZN(G57) );
  NAND2_X1 U590 ( .A1(n448), .A2(n441), .ZN(n444) );
  AND2_X1 U591 ( .A1(n445), .A2(n441), .ZN(G54) );
  XNOR2_X1 U592 ( .A(n447), .B(n446), .ZN(G60) );
  NAND2_X1 U593 ( .A1(n449), .A2(n441), .ZN(n447) );
  XNOR2_X1 U594 ( .A(n686), .B(n362), .ZN(n448) );
  XNOR2_X1 U595 ( .A(n722), .B(n364), .ZN(n449) );
  OR2_X2 U596 ( .A1(n711), .A2(n683), .ZN(n476) );
  NAND2_X1 U597 ( .A1(n559), .A2(G221), .ZN(n452) );
  NAND2_X1 U598 ( .A1(n752), .A2(G234), .ZN(n459) );
  NAND2_X1 U599 ( .A1(n611), .A2(n641), .ZN(n509) );
  XNOR2_X2 U600 ( .A(n476), .B(n356), .ZN(n611) );
  NOR2_X1 U601 ( .A1(n606), .A2(n617), .ZN(n607) );
  NAND2_X1 U602 ( .A1(n455), .A2(n741), .ZN(n742) );
  XNOR2_X1 U603 ( .A(n735), .B(KEYINPUT121), .ZN(n455) );
  XNOR2_X1 U604 ( .A(n458), .B(n501), .ZN(n502) );
  NAND2_X1 U605 ( .A1(n752), .A2(G224), .ZN(n458) );
  XNOR2_X2 U606 ( .A(n460), .B(G953), .ZN(n752) );
  OR2_X1 U607 ( .A1(n475), .A2(KEYINPUT83), .ZN(n462) );
  NAND2_X1 U608 ( .A1(n615), .A2(n514), .ZN(n466) );
  XNOR2_X2 U609 ( .A(n509), .B(KEYINPUT84), .ZN(n469) );
  NAND2_X1 U610 ( .A1(n467), .A2(n704), .ZN(n691) );
  NAND2_X1 U611 ( .A1(n467), .A2(n689), .ZN(n690) );
  NOR2_X1 U612 ( .A1(n705), .A2(n467), .ZN(n584) );
  NOR2_X1 U613 ( .A1(n623), .A2(n469), .ZN(n620) );
  NAND2_X1 U614 ( .A1(n475), .A2(n710), .ZN(n637) );
  NAND2_X1 U615 ( .A1(n475), .A2(n353), .ZN(n470) );
  NAND2_X1 U616 ( .A1(n473), .A2(n474), .ZN(n472) );
  INV_X1 U617 ( .A(n699), .ZN(n478) );
  NOR2_X2 U618 ( .A1(n680), .A2(n679), .ZN(n682) );
  XNOR2_X1 U619 ( .A(n502), .B(n507), .ZN(n487) );
  INV_X1 U620 ( .A(KEYINPUT48), .ZN(n480) );
  NAND2_X1 U621 ( .A1(n579), .A2(n578), .ZN(n482) );
  XNOR2_X1 U622 ( .A(n577), .B(n483), .ZN(n579) );
  INV_X1 U623 ( .A(KEYINPUT99), .ZN(n483) );
  XNOR2_X1 U624 ( .A(n554), .B(n530), .ZN(n484) );
  XNOR2_X1 U625 ( .A(n531), .B(n486), .ZN(n485) );
  XNOR2_X1 U626 ( .A(n532), .B(n525), .ZN(n486) );
  XNOR2_X2 U627 ( .A(n745), .B(G101), .ZN(n543) );
  INV_X1 U628 ( .A(KEYINPUT81), .ZN(n488) );
  NAND2_X1 U629 ( .A1(n682), .A2(n681), .ZN(n489) );
  NOR2_X1 U630 ( .A1(n586), .A2(n704), .ZN(n646) );
  XNOR2_X1 U631 ( .A(n524), .B(KEYINPUT98), .ZN(n525) );
  INV_X1 U632 ( .A(KEYINPUT79), .ZN(n635) );
  INV_X1 U633 ( .A(n602), .ZN(n595) );
  INV_X1 U634 ( .A(KEYINPUT59), .ZN(n720) );
  INV_X1 U635 ( .A(n655), .ZN(n621) );
  XNOR2_X1 U636 ( .A(KEYINPUT66), .B(G469), .ZN(n500) );
  XNOR2_X2 U637 ( .A(n515), .B(KEYINPUT4), .ZN(n745) );
  XNOR2_X1 U638 ( .A(G104), .B(KEYINPUT73), .ZN(n493) );
  XNOR2_X1 U639 ( .A(n493), .B(G110), .ZN(n729) );
  NAND2_X1 U640 ( .A1(G227), .A2(n752), .ZN(n495) );
  XNOR2_X1 U641 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U642 ( .A(n497), .B(n545), .ZN(n498) );
  XNOR2_X1 U643 ( .A(n503), .B(n498), .ZN(n715) );
  NOR2_X1 U644 ( .A1(G902), .A2(n715), .ZN(n499) );
  XNOR2_X1 U645 ( .A(KEYINPUT87), .B(G113), .ZN(n504) );
  XOR2_X1 U646 ( .A(KEYINPUT89), .B(G898), .Z(n739) );
  NOR2_X1 U647 ( .A1(n739), .A2(n510), .ZN(n732) );
  NAND2_X1 U648 ( .A1(G902), .A2(n732), .ZN(n511) );
  NAND2_X1 U649 ( .A1(G952), .A2(n510), .ZN(n592) );
  AND2_X1 U650 ( .A1(n511), .A2(n592), .ZN(n513) );
  XNOR2_X1 U651 ( .A(n512), .B(KEYINPUT14), .ZN(n594) );
  INV_X1 U652 ( .A(n594), .ZN(n672) );
  NOR2_X1 U653 ( .A1(n513), .A2(n672), .ZN(n514) );
  XOR2_X1 U654 ( .A(KEYINPUT9), .B(n515), .Z(n517) );
  NAND2_X1 U655 ( .A1(G217), .A2(n559), .ZN(n520) );
  XNOR2_X1 U656 ( .A(G478), .B(n521), .ZN(n578) );
  INV_X1 U657 ( .A(n578), .ZN(n565) );
  XNOR2_X1 U658 ( .A(n523), .B(n522), .ZN(n532) );
  XOR2_X1 U659 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n527) );
  XNOR2_X1 U660 ( .A(KEYINPUT96), .B(KEYINPUT12), .ZN(n526) );
  XNOR2_X1 U661 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U662 ( .A(G143), .B(n528), .ZN(n531) );
  NOR2_X1 U663 ( .A1(G953), .A2(G237), .ZN(n529) );
  XOR2_X1 U664 ( .A(KEYINPUT75), .B(n529), .Z(n541) );
  NAND2_X1 U665 ( .A1(n541), .A2(G214), .ZN(n530) );
  INV_X1 U666 ( .A(G475), .ZN(n534) );
  NOR2_X1 U667 ( .A1(n565), .A2(n577), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n679), .A2(G234), .ZN(n537) );
  XNOR2_X1 U669 ( .A(n537), .B(KEYINPUT20), .ZN(n551) );
  NAND2_X1 U670 ( .A1(G221), .A2(n551), .ZN(n538) );
  XNOR2_X1 U671 ( .A(KEYINPUT21), .B(n538), .ZN(n603) );
  AND2_X1 U672 ( .A1(n600), .A2(n563), .ZN(n539) );
  NAND2_X1 U673 ( .A1(n541), .A2(G210), .ZN(n549) );
  XNOR2_X1 U674 ( .A(n542), .B(n543), .ZN(n548) );
  XNOR2_X1 U675 ( .A(n544), .B(KEYINPUT5), .ZN(n546) );
  XOR2_X1 U676 ( .A(n546), .B(n545), .Z(n547) );
  INV_X1 U677 ( .A(KEYINPUT71), .ZN(n550) );
  XOR2_X1 U678 ( .A(KEYINPUT25), .B(KEYINPUT93), .Z(n553) );
  NAND2_X1 U679 ( .A1(n551), .A2(G217), .ZN(n552) );
  XOR2_X1 U680 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n557) );
  XNOR2_X1 U681 ( .A(n557), .B(n556), .ZN(n558) );
  NOR2_X1 U682 ( .A1(n616), .A2(n605), .ZN(n562) );
  NAND2_X1 U683 ( .A1(n570), .A2(n562), .ZN(n688) );
  NAND2_X1 U684 ( .A1(n580), .A2(n616), .ZN(n564) );
  NAND2_X1 U685 ( .A1(n565), .A2(n577), .ZN(n613) );
  XNOR2_X1 U686 ( .A(KEYINPUT77), .B(n613), .ZN(n566) );
  NAND2_X1 U687 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U688 ( .A1(n658), .A2(n650), .ZN(n569) );
  NOR2_X1 U689 ( .A1(n572), .A2(n650), .ZN(n574) );
  NOR2_X1 U690 ( .A1(n655), .A2(n616), .ZN(n573) );
  NAND2_X1 U691 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U692 ( .A1(n579), .A2(n578), .ZN(n704) );
  NAND2_X1 U693 ( .A1(n658), .A2(n580), .ZN(n661) );
  XNOR2_X1 U694 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n581) );
  XNOR2_X1 U695 ( .A(n582), .B(n581), .ZN(n705) );
  INV_X1 U696 ( .A(n681), .ZN(n734) );
  BUF_X1 U697 ( .A(n586), .Z(n689) );
  NAND2_X1 U698 ( .A1(n641), .A2(n658), .ZN(n589) );
  INV_X1 U699 ( .A(KEYINPUT30), .ZN(n587) );
  NOR2_X1 U700 ( .A1(n752), .A2(G900), .ZN(n590) );
  NAND2_X1 U701 ( .A1(G902), .A2(n590), .ZN(n591) );
  NAND2_X1 U702 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U703 ( .A1(n594), .A2(n593), .ZN(n602) );
  INV_X1 U704 ( .A(n600), .ZN(n644) );
  INV_X1 U705 ( .A(KEYINPUT41), .ZN(n601) );
  NOR2_X1 U706 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U707 ( .A(KEYINPUT28), .B(n607), .Z(n608) );
  NAND2_X1 U708 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U709 ( .A1(n613), .A2(n612), .ZN(n699) );
  NAND2_X1 U710 ( .A1(n615), .A2(n614), .ZN(n695) );
  INV_X1 U711 ( .A(n616), .ZN(n618) );
  NOR2_X1 U712 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U713 ( .A1(n619), .A2(n689), .ZN(n623) );
  XNOR2_X1 U714 ( .A(KEYINPUT36), .B(n620), .ZN(n622) );
  NAND2_X1 U715 ( .A1(n622), .A2(n621), .ZN(n708) );
  INV_X1 U716 ( .A(n623), .ZN(n624) );
  NAND2_X1 U717 ( .A1(n624), .A2(n641), .ZN(n625) );
  XNOR2_X1 U718 ( .A(n625), .B(KEYINPUT103), .ZN(n626) );
  NAND2_X1 U719 ( .A1(n626), .A2(n655), .ZN(n629) );
  XOR2_X1 U720 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n627) );
  XNOR2_X1 U721 ( .A(KEYINPUT43), .B(n627), .ZN(n628) );
  XNOR2_X1 U722 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U723 ( .A1(n631), .A2(n630), .ZN(n710) );
  NAND2_X1 U724 ( .A1(n632), .A2(n704), .ZN(n709) );
  INV_X1 U725 ( .A(n709), .ZN(n633) );
  NOR2_X1 U726 ( .A1(n634), .A2(KEYINPUT2), .ZN(n636) );
  XNOR2_X1 U727 ( .A(n636), .B(n635), .ZN(n639) );
  NAND2_X1 U728 ( .A1(KEYINPUT2), .A2(n709), .ZN(n638) );
  BUF_X1 U729 ( .A(n640), .Z(n664) );
  NOR2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U733 ( .A(n649), .B(KEYINPUT113), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n652), .B(KEYINPUT112), .ZN(n653) );
  XNOR2_X1 U736 ( .A(n653), .B(KEYINPUT49), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U738 ( .A(KEYINPUT50), .B(n656), .Z(n657) );
  NOR2_X1 U739 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U742 ( .A(KEYINPUT51), .B(n663), .Z(n665) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(KEYINPUT114), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n669), .B(KEYINPUT52), .ZN(n670) );
  NAND2_X1 U747 ( .A1(n670), .A2(G952), .ZN(n671) );
  NOR2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U749 ( .A1(G953), .A2(n673), .ZN(n674) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(KEYINPUT116), .Z(n677) );
  INV_X1 U751 ( .A(KEYINPUT115), .ZN(n676) );
  XNOR2_X1 U752 ( .A(n677), .B(n676), .ZN(n678) );
  NAND2_X1 U753 ( .A1(n723), .A2(G472), .ZN(n686) );
  XOR2_X1 U754 ( .A(G101), .B(KEYINPUT109), .Z(n687) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(G3) );
  INV_X1 U756 ( .A(n689), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n690), .B(G104), .ZN(G6) );
  XNOR2_X1 U758 ( .A(G107), .B(KEYINPUT27), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT26), .B(KEYINPUT110), .Z(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U761 ( .A(n694), .B(n693), .ZN(G9) );
  INV_X1 U762 ( .A(n704), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U764 ( .A(G128), .B(KEYINPUT29), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n698), .B(n697), .ZN(G30) );
  XOR2_X1 U766 ( .A(G143), .B(n699), .Z(G45) );
  NOR2_X1 U767 ( .A1(n700), .A2(n695), .ZN(n701) );
  XOR2_X1 U768 ( .A(G146), .B(n701), .Z(G48) );
  XOR2_X1 U769 ( .A(G113), .B(KEYINPUT111), .Z(n703) );
  NAND2_X1 U770 ( .A1(n705), .A2(n689), .ZN(n702) );
  XNOR2_X1 U771 ( .A(n703), .B(n702), .ZN(G15) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U773 ( .A(n706), .B(G116), .ZN(G18) );
  XOR2_X1 U774 ( .A(G125), .B(KEYINPUT37), .Z(n707) );
  XNOR2_X1 U775 ( .A(n708), .B(n707), .ZN(G27) );
  XNOR2_X1 U776 ( .A(G134), .B(n709), .ZN(G36) );
  XNOR2_X1 U777 ( .A(G140), .B(n710), .ZN(G42) );
  XOR2_X1 U778 ( .A(KEYINPUT86), .B(KEYINPUT55), .Z(n713) );
  XNOR2_X1 U779 ( .A(n711), .B(KEYINPUT54), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n723), .A2(G210), .ZN(n714) );
  XOR2_X1 U781 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  XNOR2_X1 U782 ( .A(n715), .B(KEYINPUT117), .ZN(n716) );
  XNOR2_X1 U783 ( .A(n717), .B(n716), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n723), .A2(G469), .ZN(n718) );
  NAND2_X1 U785 ( .A1(n723), .A2(G475), .ZN(n722) );
  NAND2_X1 U786 ( .A1(G217), .A2(n723), .ZN(n725) );
  XNOR2_X1 U787 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n728), .A2(n727), .ZN(G66) );
  XOR2_X1 U789 ( .A(G101), .B(n729), .Z(n730) );
  XNOR2_X1 U790 ( .A(n731), .B(n730), .ZN(n733) );
  NOR2_X1 U791 ( .A1(n733), .A2(n732), .ZN(n744) );
  XOR2_X1 U792 ( .A(KEYINPUT61), .B(KEYINPUT119), .Z(n737) );
  NAND2_X1 U793 ( .A1(G224), .A2(G953), .ZN(n736) );
  XNOR2_X1 U794 ( .A(n737), .B(n736), .ZN(n738) );
  NAND2_X1 U795 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U796 ( .A(KEYINPUT120), .B(n740), .ZN(n741) );
  XNOR2_X1 U797 ( .A(n742), .B(KEYINPUT123), .ZN(n743) );
  XNOR2_X1 U798 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U799 ( .A(G227), .B(n751), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(G900), .ZN(n749) );
  XNOR2_X1 U801 ( .A(KEYINPUT124), .B(n749), .ZN(n750) );
  NAND2_X1 U802 ( .A1(n750), .A2(G953), .ZN(n755) );
  NAND2_X1 U803 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n755), .A2(n754), .ZN(G72) );
  XNOR2_X1 U805 ( .A(n756), .B(G137), .ZN(G39) );
  XNOR2_X1 U806 ( .A(n757), .B(G131), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n758), .B(KEYINPUT126), .ZN(G33) );
  XOR2_X1 U808 ( .A(n759), .B(G122), .Z(G24) );
  XOR2_X1 U809 ( .A(n760), .B(G119), .Z(n761) );
  XNOR2_X1 U810 ( .A(KEYINPUT125), .B(n761), .ZN(G21) );
endmodule

