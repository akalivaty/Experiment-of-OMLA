//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G77), .A2(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(G97), .A2(G257), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n206), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(new_n201), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n219), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n210), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  NAND2_X1  g0040(.A1(G68), .A2(G77), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n203), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(new_n209), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(G20), .B1(new_n221), .B2(G50), .ZN(new_n250));
  INV_X1    g0050(.A(G150), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n225), .A2(G33), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n250), .B1(new_n251), .B2(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n224), .ZN(new_n258));
  INV_X1    g0058(.A(G50), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n256), .A2(new_n258), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n258), .B1(new_n260), .B2(G20), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n259), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT66), .A2(G223), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT66), .A2(G223), .ZN(new_n268));
  OAI21_X1  g0068(.A(G1698), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G222), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n273), .B(new_n277), .C1(G77), .C2(new_n270), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n276), .A2(new_n279), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G226), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n278), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n266), .B1(new_n285), .B2(G179), .ZN(new_n286));
  INV_X1    g0086(.A(G169), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT9), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n266), .A2(new_n290), .B1(G200), .B2(new_n285), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n291), .B(new_n293), .C1(new_n290), .C2(new_n266), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(KEYINPUT10), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n289), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT13), .ZN(new_n298));
  AND2_X1   g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  NOR2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  OAI211_X1 g0100(.A(G232), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT67), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n270), .A2(KEYINPUT67), .A3(G232), .A4(G1698), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G97), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n270), .A2(G226), .A3(new_n271), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n277), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n283), .A2(G238), .ZN(new_n309));
  AND4_X1   g0109(.A1(new_n298), .A2(new_n308), .A3(new_n282), .A4(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n281), .B1(new_n307), .B2(new_n277), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n298), .B1(new_n311), .B2(new_n309), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n313), .A2(new_n287), .B1(KEYINPUT70), .B2(KEYINPUT14), .ZN(new_n314));
  NAND2_X1  g0114(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n309), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n311), .A2(new_n298), .A3(new_n309), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(G169), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n313), .A2(G179), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n314), .A2(new_n315), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n201), .A2(G20), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n324), .B1(new_n254), .B2(new_n202), .C1(new_n253), .C2(new_n259), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n258), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n262), .A2(new_n201), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT12), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n325), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n264), .A2(G68), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n328), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT69), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n323), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n317), .A2(G190), .A3(new_n318), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT68), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n317), .A2(new_n338), .A3(G190), .A4(new_n318), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n334), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n341), .B1(new_n317), .B2(new_n318), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n299), .A2(new_n300), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G232), .B2(new_n271), .ZN(new_n346));
  INV_X1    g0146(.A(G238), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(new_n271), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n277), .C1(G107), .C2(new_n270), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n283), .A2(G244), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n282), .A3(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(G179), .ZN(new_n352));
  INV_X1    g0152(.A(new_n255), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n354));
  XOR2_X1   g0154(.A(KEYINPUT15), .B(G87), .Z(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n356), .B2(new_n254), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n258), .B1(new_n202), .B2(new_n262), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(new_n202), .B2(new_n265), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n351), .A2(new_n287), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n352), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n297), .A2(new_n335), .A3(new_n344), .A4(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n220), .A2(new_n201), .ZN(new_n363));
  NOR2_X1   g0163(.A1(G58), .A2(G68), .ZN(new_n364));
  OAI21_X1  g0164(.A(G20), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(KEYINPUT72), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n252), .A2(G159), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT72), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n368), .B(G20), .C1(new_n363), .C2(new_n364), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  NOR4_X1   g0171(.A1(new_n299), .A2(new_n300), .A3(new_n371), .A4(G20), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n299), .A2(new_n300), .A3(G20), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT71), .B1(new_n373), .B2(KEYINPUT7), .ZN(new_n374));
  OR2_X1    g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  NAND2_X1  g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n225), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT71), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n371), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n372), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT16), .B(new_n370), .C1(new_n380), .C2(new_n201), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  INV_X1    g0182(.A(new_n372), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n377), .A2(new_n371), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n201), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n381), .A2(new_n258), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n255), .A2(new_n261), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n264), .B2(new_n255), .ZN(new_n390));
  OAI211_X1 g0190(.A(G226), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n391));
  OAI211_X1 g0191(.A(G223), .B(new_n271), .C1(new_n299), .C2(new_n300), .ZN(new_n392));
  INV_X1    g0192(.A(G87), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n391), .B(new_n392), .C1(new_n274), .C2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n281), .B1(new_n394), .B2(new_n277), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n276), .A2(G232), .A3(new_n279), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n292), .A3(new_n397), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n281), .B(new_n396), .C1(new_n394), .C2(new_n277), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(G200), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n388), .A2(new_n390), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT17), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT17), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n388), .A2(new_n400), .A3(new_n403), .A4(new_n390), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n402), .A2(KEYINPUT73), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT73), .B1(new_n402), .B2(new_n404), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n388), .A2(new_n390), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n395), .A2(G179), .A3(new_n397), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n287), .B1(new_n395), .B2(new_n397), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n408), .A2(new_n412), .A3(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n359), .B1(G200), .B2(new_n351), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n292), .B2(new_n351), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n407), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n362), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT77), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n260), .A2(G45), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n426));
  INV_X1    g0226(.A(G45), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(G1), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT5), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G41), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(KEYINPUT77), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n425), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G270), .A3(new_n276), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT80), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT80), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n432), .A2(new_n435), .A3(G270), .A4(new_n276), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(G257), .B(new_n271), .C1(new_n299), .C2(new_n300), .ZN(new_n438));
  OAI211_X1 g0238(.A(G264), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n375), .A2(G303), .A3(new_n376), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n277), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n425), .A2(new_n431), .A3(G274), .A4(new_n426), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n277), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n437), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G200), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n434), .B2(new_n436), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G190), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n260), .A2(G33), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n261), .A2(new_n450), .A3(new_n224), .A4(new_n257), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G116), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n262), .A2(new_n209), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n257), .A2(new_n224), .B1(G20), .B2(new_n209), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n456), .B(new_n225), .C1(G33), .C2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n455), .A2(KEYINPUT20), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT20), .B1(new_n455), .B2(new_n458), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n453), .B(new_n454), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n447), .A2(new_n449), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(G169), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n437), .B2(new_n445), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT21), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT21), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n448), .B2(new_n465), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n448), .A2(G179), .A3(new_n461), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT81), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n437), .A2(new_n445), .A3(G179), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(new_n461), .B1(new_n466), .B2(KEYINPUT21), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(new_n463), .A3(new_n475), .A4(new_n469), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G107), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n451), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(KEYINPUT22), .B(G87), .C1(new_n299), .C2(new_n300), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n225), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n270), .A2(new_n225), .A3(G87), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT22), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT23), .ZN(new_n487));
  OAI211_X1 g0287(.A(G20), .B(new_n478), .C1(new_n487), .C2(KEYINPUT83), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n489));
  XNOR2_X1  g0289(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n483), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(KEYINPUT82), .B(KEYINPUT24), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n491), .B(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n479), .B1(new_n494), .B2(new_n258), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n270), .A2(G257), .A3(G1698), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n270), .A2(G250), .A3(new_n271), .ZN(new_n497));
  INV_X1    g0297(.A(G294), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n496), .B(new_n497), .C1(new_n274), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n277), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n432), .A2(G264), .A3(new_n276), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n443), .A2(new_n277), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n500), .A2(new_n504), .A3(new_n501), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G190), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n262), .B(new_n478), .C1(KEYINPUT84), .C2(KEYINPUT25), .ZN(new_n509));
  NAND2_X1  g0309(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n495), .A2(new_n506), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n491), .A2(new_n493), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n482), .A2(new_n225), .B1(new_n484), .B2(new_n485), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n492), .B1(new_n514), .B2(new_n490), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n258), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n479), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(new_n517), .A3(new_n511), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n505), .A2(new_n287), .ZN(new_n519));
  INV_X1    g0319(.A(G179), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n507), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n261), .A2(KEYINPUT75), .A3(G97), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n261), .A2(G97), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT75), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n451), .A2(new_n457), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT7), .B1(new_n345), .B2(new_n225), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n528), .B2(new_n372), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT74), .B1(new_n252), .B2(G77), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  AND2_X1   g0331(.A1(G97), .A2(G107), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n478), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n530), .B1(new_n536), .B2(G20), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n252), .A2(KEYINPUT74), .A3(G77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n529), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n524), .B(new_n527), .C1(new_n539), .C2(new_n258), .ZN(new_n540));
  OAI211_X1 g0340(.A(G244), .B(new_n271), .C1(new_n299), .C2(new_n300), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n270), .A2(KEYINPUT4), .A3(G244), .A4(new_n271), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(new_n456), .ZN(new_n545));
  OAI211_X1 g0345(.A(G250), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT76), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT76), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n270), .A2(new_n548), .A3(G250), .A4(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n277), .B1(new_n545), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n432), .A2(G257), .A3(new_n276), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n504), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n540), .B(new_n554), .C1(new_n292), .C2(new_n553), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n355), .A2(new_n261), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n225), .B1(new_n305), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n533), .A2(new_n393), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n225), .A2(G33), .A3(G97), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n558), .A2(new_n559), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n270), .A2(new_n225), .A3(G68), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n556), .B1(new_n563), .B2(new_n258), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n452), .A2(new_n355), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G238), .B(new_n271), .C1(new_n299), .C2(new_n300), .ZN(new_n567));
  OAI211_X1 g0367(.A(G244), .B(G1698), .C1(new_n299), .C2(new_n300), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(new_n568), .A3(new_n481), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n277), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n260), .A2(G45), .A3(G274), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT78), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT78), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n573), .A2(new_n260), .A3(G45), .A4(G274), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  AND2_X1   g0376(.A1(G33), .A2(G41), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n424), .B(G250), .C1(new_n577), .C2(new_n224), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n576), .B1(new_n575), .B2(new_n578), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n520), .B(new_n570), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n573), .B1(new_n428), .B2(G274), .ZN(new_n582));
  INV_X1    g0382(.A(new_n574), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(KEYINPUT79), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n586));
  AOI22_X1  g0386(.A1(new_n585), .A2(new_n586), .B1(new_n277), .B2(new_n569), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n566), .B(new_n581), .C1(new_n587), .C2(G169), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n451), .A2(new_n393), .ZN(new_n589));
  AOI211_X1 g0389(.A(new_n556), .B(new_n589), .C1(new_n563), .C2(new_n258), .ZN(new_n590));
  OAI211_X1 g0390(.A(G190), .B(new_n570), .C1(new_n579), .C2(new_n580), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n587), .C2(new_n341), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n553), .A2(new_n287), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n539), .A2(new_n258), .ZN(new_n595));
  INV_X1    g0395(.A(new_n524), .ZN(new_n596));
  INV_X1    g0396(.A(new_n527), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n551), .A2(new_n504), .A3(new_n520), .A4(new_n552), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n555), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n523), .A2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n421), .A2(new_n477), .A3(new_n602), .ZN(G372));
  AND2_X1   g0403(.A1(new_n323), .A2(new_n334), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n361), .B1(new_n340), .B2(new_n343), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT87), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT87), .ZN(new_n607));
  AOI211_X1 g0407(.A(new_n342), .B(new_n334), .C1(new_n337), .C2(new_n339), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n335), .B(new_n607), .C1(new_n608), .C2(new_n361), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n606), .A2(new_n407), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n417), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n295), .A2(new_n296), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n289), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n421), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n588), .A2(new_n592), .ZN(new_n615));
  XNOR2_X1  g0415(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n600), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n600), .A2(new_n615), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n588), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n471), .A2(KEYINPUT85), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT85), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n467), .A2(new_n469), .A3(new_n622), .A4(new_n470), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n522), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n508), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n507), .A2(new_n341), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n518), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n601), .ZN(new_n628));
  AOI211_X1 g0428(.A(new_n617), .B(new_n620), .C1(new_n624), .C2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n613), .B1(new_n614), .B2(new_n629), .ZN(G369));
  NAND2_X1  g0430(.A1(new_n621), .A2(new_n623), .ZN(new_n631));
  INV_X1    g0431(.A(G13), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(G20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n260), .ZN(new_n634));
  OR2_X1    g0434(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(KEYINPUT27), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(G213), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(G343), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n461), .ZN(new_n640));
  MUX2_X1   g0440(.A(new_n631), .B(new_n477), .S(new_n640), .Z(new_n641));
  XNOR2_X1  g0441(.A(KEYINPUT88), .B(G330), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n518), .A2(new_n639), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n512), .A2(new_n522), .A3(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(KEYINPUT89), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n522), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n639), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n639), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n471), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n646), .B2(new_n647), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n522), .A2(new_n639), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n657), .ZN(G399));
  INV_X1    g0458(.A(new_n228), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n559), .A2(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G1), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n222), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT28), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT91), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n620), .B1(new_n624), .B2(new_n628), .ZN(new_n667));
  INV_X1    g0467(.A(new_n617), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n639), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n666), .B1(new_n669), .B2(KEYINPUT29), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n551), .A2(new_n504), .A3(new_n552), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n527), .B1(new_n539), .B2(new_n258), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n671), .A2(new_n520), .B1(new_n672), .B2(new_n596), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n593), .A2(new_n619), .A3(new_n673), .A4(new_n594), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n616), .B1(new_n600), .B2(new_n615), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n588), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT92), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n522), .A2(new_n474), .A3(new_n469), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n555), .A2(new_n593), .A3(new_n600), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n512), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT92), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n674), .A2(new_n675), .A3(new_n681), .A4(new_n588), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n683), .A2(KEYINPUT29), .A3(new_n653), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT29), .ZN(new_n685));
  OAI211_X1 g0485(.A(KEYINPUT91), .B(new_n685), .C1(new_n629), .C2(new_n639), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n670), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n477), .A2(new_n602), .A3(new_n653), .ZN(new_n688));
  INV_X1    g0488(.A(new_n587), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n505), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n551), .A2(new_n552), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n473), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n507), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  AOI21_X1  g0497(.A(G179), .B1(new_n587), .B2(KEYINPUT90), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n697), .A2(new_n446), .A3(new_n553), .A4(new_n698), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n690), .A2(KEYINPUT30), .A3(new_n473), .A4(new_n692), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n695), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n639), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n688), .A2(KEYINPUT31), .A3(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(KEYINPUT31), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n642), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n687), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT93), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n687), .A2(new_n706), .A3(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n665), .B1(new_n711), .B2(G1), .ZN(G364));
  AOI21_X1  g0512(.A(new_n260), .B1(new_n633), .B2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n660), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n659), .A2(new_n270), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n223), .A2(new_n427), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n717), .B(new_n718), .C1(new_n245), .C2(new_n427), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n270), .A2(G355), .A3(new_n228), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n719), .B(new_n720), .C1(G116), .C2(new_n228), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n224), .B1(G20), .B2(new_n287), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n716), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n726), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n225), .A2(G190), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G179), .A2(G200), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G159), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT32), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n341), .A2(G179), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G107), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n225), .B1(new_n731), .B2(G190), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n457), .ZN(new_n744));
  NAND3_X1  g0544(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n292), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n744), .B1(new_n746), .B2(G50), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n225), .A2(new_n292), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n739), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n393), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n520), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n730), .A2(new_n751), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n752), .A2(new_n220), .B1(new_n753), .B2(new_n202), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n745), .A2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n270), .B1(new_n756), .B2(new_n201), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n750), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n738), .A2(new_n742), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT96), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G303), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n345), .B1(new_n743), .B2(new_n498), .C1(new_n763), .C2(new_n749), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT97), .B(G326), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n762), .B(new_n764), .C1(new_n746), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G322), .ZN(new_n767));
  INV_X1    g0567(.A(G311), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n752), .A2(new_n767), .B1(new_n753), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n735), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(G329), .ZN(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n766), .B(new_n771), .C1(new_n772), .C2(new_n740), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n760), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n725), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n728), .B1(new_n729), .B2(new_n774), .C1(new_n641), .C2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n643), .A2(new_n716), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n641), .A2(new_n642), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(G396));
  NAND2_X1  g0579(.A1(new_n770), .A2(G311), .ZN(new_n780));
  INV_X1    g0580(.A(new_n753), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G116), .ZN(new_n782));
  INV_X1    g0582(.A(new_n746), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n756), .A2(new_n772), .B1(new_n783), .B2(new_n763), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n345), .B1(new_n740), .B2(new_n393), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n784), .A2(new_n744), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n749), .ZN(new_n787));
  INV_X1    g0587(.A(new_n752), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G107), .A2(new_n787), .B1(new_n788), .B2(G294), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n780), .A2(new_n782), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n781), .A2(G159), .B1(G137), .B2(new_n746), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(new_n251), .B2(new_n756), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(G143), .B2(new_n788), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT34), .ZN(new_n794));
  INV_X1    g0594(.A(G132), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n270), .B1(new_n735), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT98), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT98), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n741), .A2(G68), .ZN(new_n799));
  INV_X1    g0599(.A(new_n743), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n787), .A2(G50), .B1(new_n800), .B2(G58), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n790), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n726), .A2(new_n723), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(new_n726), .B1(new_n202), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n359), .A2(new_n639), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n419), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n361), .ZN(new_n808));
  INV_X1    g0608(.A(new_n361), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n653), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n715), .B(new_n805), .C1(new_n811), .C2(new_n724), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n812), .B(KEYINPUT99), .Z(new_n813));
  XNOR2_X1  g0613(.A(new_n669), .B(new_n811), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n706), .B(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n813), .B1(new_n815), .B2(new_n715), .ZN(G384));
  INV_X1    g0616(.A(KEYINPUT40), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT38), .ZN(new_n818));
  INV_X1    g0618(.A(new_n258), .ZN(new_n819));
  INV_X1    g0619(.A(new_n379), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n378), .B1(new_n377), .B2(new_n371), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n383), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n386), .B1(new_n822), .B2(G68), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n819), .B1(new_n823), .B2(KEYINPUT16), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(KEYINPUT16), .B2(new_n823), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n825), .A2(new_n390), .B1(new_n411), .B2(new_n637), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n388), .A2(new_n390), .A3(new_n400), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT37), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n637), .B(KEYINPUT100), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n408), .B1(new_n412), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n401), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n402), .A2(new_n404), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT73), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n402), .A2(KEYINPUT73), .A3(new_n404), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(new_n417), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n637), .B1(new_n825), .B2(new_n390), .ZN(new_n840));
  AOI221_X4 g0640(.A(new_n818), .B1(new_n828), .B2(new_n834), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n828), .A2(new_n834), .ZN(new_n843));
  AOI21_X1  g0643(.A(KEYINPUT38), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n334), .B(new_n639), .C1(new_n608), .C2(new_n323), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n334), .A2(new_n639), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n335), .A2(new_n344), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n703), .A2(new_n849), .A3(new_n704), .A4(new_n811), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n817), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  AND4_X1   g0651(.A1(new_n703), .A2(new_n849), .A3(new_n704), .A4(new_n811), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n843), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n411), .A2(new_n829), .B1(new_n388), .B2(new_n390), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n832), .B1(new_n854), .B2(new_n827), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT102), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n834), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n854), .A2(new_n827), .A3(new_n832), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT102), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n415), .A2(new_n416), .B1(new_n402), .B2(new_n404), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n829), .B1(new_n388), .B2(new_n390), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n857), .B(new_n859), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n818), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n817), .B1(new_n853), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n852), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n851), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n705), .A2(new_n421), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n642), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n670), .A2(new_n421), .A3(new_n684), .A4(new_n686), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n613), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n870), .B(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n846), .A2(new_n848), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n624), .A2(new_n628), .ZN(new_n875));
  INV_X1    g0675(.A(new_n620), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n668), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n653), .A3(new_n811), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n874), .B1(new_n878), .B2(new_n810), .ZN(new_n879));
  INV_X1    g0679(.A(new_n840), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n407), .B2(new_n417), .ZN(new_n881));
  INV_X1    g0681(.A(new_n843), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n818), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n853), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n415), .A2(new_n416), .A3(new_n829), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n883), .B2(new_n853), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n853), .A2(new_n864), .A3(new_n887), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n335), .A2(new_n639), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n885), .B(new_n886), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n873), .B(new_n893), .Z(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n260), .B2(new_n633), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n209), .B1(new_n536), .B2(KEYINPUT35), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n896), .B(new_n226), .C1(KEYINPUT35), .C2(new_n536), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT36), .ZN(new_n898));
  OAI21_X1  g0698(.A(G77), .B1(new_n220), .B2(new_n201), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n222), .A2(new_n899), .B1(G50), .B2(new_n201), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(G1), .A3(new_n632), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(new_n898), .A3(new_n901), .ZN(G367));
  NOR2_X1   g0702(.A1(new_n600), .A2(new_n653), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT104), .Z(new_n904));
  OAI211_X1 g0704(.A(new_n555), .B(new_n600), .C1(new_n540), .C2(new_n653), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n652), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n653), .A2(new_n590), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT103), .ZN(new_n911));
  MUX2_X1   g0711(.A(new_n588), .B(new_n615), .S(new_n911), .Z(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n655), .A2(new_n906), .ZN(new_n915));
  OR3_X1    g0715(.A1(new_n915), .A2(KEYINPUT105), .A3(KEYINPUT42), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n600), .B1(new_n907), .B2(new_n522), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n653), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT105), .B1(new_n915), .B2(KEYINPUT42), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n916), .A2(new_n918), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n909), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n909), .B1(new_n921), .B2(new_n914), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OR3_X1    g0726(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n923), .B2(new_n924), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n660), .B(KEYINPUT41), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n657), .A2(new_n906), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT106), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT106), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n657), .A2(new_n933), .A3(new_n906), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT45), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n657), .A2(new_n906), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT44), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(KEYINPUT45), .A3(new_n934), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT107), .B1(new_n941), .B2(new_n651), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n651), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  MUX2_X1   g0744(.A(new_n648), .B(new_n650), .S(new_n654), .Z(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n643), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n709), .B2(new_n710), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n941), .A2(KEYINPUT107), .A3(new_n651), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n930), .B1(new_n949), .B2(new_n711), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n927), .B(new_n928), .C1(new_n950), .C2(new_n714), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n345), .B1(new_n740), .B2(new_n457), .C1(new_n772), .C2(new_n753), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n783), .A2(new_n768), .B1(new_n743), .B2(new_n478), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n954), .B1(new_n955), .B2(new_n735), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT108), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n787), .A2(KEYINPUT46), .A3(G116), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT46), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n749), .B2(new_n209), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n960), .C1(new_n498), .C2(new_n756), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n956), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n962), .B1(new_n957), .B2(new_n961), .C1(new_n763), .C2(new_n752), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n752), .A2(new_n251), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n743), .A2(new_n201), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n270), .B1(new_n740), .B2(new_n202), .C1(new_n220), .C2(new_n749), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(G143), .C2(new_n746), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n756), .A2(new_n736), .B1(new_n753), .B2(new_n259), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n770), .A2(G137), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n963), .B1(new_n964), .B2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT47), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n716), .B1(new_n973), .B2(new_n726), .ZN(new_n974));
  INV_X1    g0774(.A(new_n717), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n727), .B1(new_n228), .B2(new_n356), .C1(new_n239), .C2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(new_n775), .C2(new_n913), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n951), .A2(new_n977), .ZN(G387));
  AND2_X1   g0778(.A1(new_n770), .A2(new_n765), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n781), .A2(G303), .B1(G322), .B2(new_n746), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n768), .B2(new_n756), .C1(new_n955), .C2(new_n752), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT48), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n772), .B2(new_n743), .C1(new_n498), .C2(new_n749), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT49), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n270), .B(new_n979), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n984), .B2(new_n983), .C1(new_n209), .C2(new_n740), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n749), .A2(new_n202), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G50), .B2(new_n788), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n735), .B2(new_n251), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n356), .A2(new_n743), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n755), .B2(new_n353), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n345), .B1(new_n741), .B2(G97), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n736), .C2(new_n783), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n989), .B(new_n993), .C1(G68), .C2(new_n781), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT111), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n986), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n716), .B1(new_n996), .B2(new_n726), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(new_n353), .B2(new_n259), .ZN(new_n999));
  INV_X1    g0799(.A(new_n662), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n353), .A2(new_n998), .A3(new_n259), .ZN(new_n1002));
  AND4_X1   g0802(.A1(new_n427), .A2(new_n1001), .A3(new_n241), .A4(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n717), .B1(new_n236), .B2(new_n427), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n228), .A3(new_n270), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n228), .A2(G107), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n727), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n650), .A2(new_n725), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n997), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n946), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n660), .B1(new_n1011), .B2(new_n711), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1010), .B1(new_n713), .B2(new_n946), .C1(new_n1012), .C2(new_n947), .ZN(G393));
  OR2_X1    g0813(.A1(new_n941), .A2(new_n651), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT112), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n1015), .A3(new_n943), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n941), .A2(KEYINPUT112), .A3(new_n651), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n660), .B(new_n949), .C1(new_n1018), .C2(new_n947), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n907), .A2(new_n725), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n727), .B1(new_n457), .B2(new_n228), .C1(new_n248), .C2(new_n975), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n735), .A2(new_n767), .B1(new_n772), .B2(new_n749), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT113), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n788), .A2(G311), .B1(G317), .B2(new_n746), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n270), .B(new_n1025), .C1(G294), .C2(new_n781), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n742), .B1(new_n209), .B2(new_n743), .C1(new_n756), .C2(new_n763), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT52), .B2(new_n1024), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1023), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n749), .A2(new_n201), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n743), .A2(new_n202), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n270), .B1(new_n740), .B2(new_n393), .C1(new_n255), .C2(new_n753), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(G50), .C2(new_n755), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n783), .A2(new_n251), .B1(new_n752), .B2(new_n736), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT51), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n770), .A2(G143), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1029), .B1(new_n1030), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n716), .B1(new_n1038), .B2(new_n726), .ZN(new_n1039));
  AND3_X1   g0839(.A1(new_n1020), .A2(new_n1021), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n1018), .B2(new_n714), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1019), .A2(new_n1041), .ZN(G390));
  OAI21_X1  g0842(.A(KEYINPUT39), .B1(new_n841), .B2(new_n844), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n853), .A2(new_n864), .A3(new_n887), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(new_n879), .C2(new_n891), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n408), .A2(new_n412), .A3(KEYINPUT18), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT18), .B1(new_n408), .B2(new_n412), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n835), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1048), .A2(new_n861), .B1(KEYINPUT102), .B2(new_n858), .ZN(new_n1049));
  AOI21_X1  g0849(.A(KEYINPUT38), .B1(new_n1049), .B2(new_n857), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n892), .B1(new_n841), .B2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n683), .A2(new_n653), .A3(new_n808), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1052), .A2(new_n810), .B1(new_n848), .B2(new_n846), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n703), .A2(new_n642), .A3(new_n704), .A4(new_n811), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(new_n874), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1045), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n669), .A2(new_n808), .B1(new_n809), .B2(new_n653), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n892), .B1(new_n1059), .B2(new_n874), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1058), .B1(new_n890), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(G330), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n850), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1057), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n890), .A2(new_n723), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n755), .A2(G137), .B1(new_n746), .B2(G128), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n800), .A2(G159), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n270), .B1(new_n740), .B2(new_n259), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n749), .A2(new_n251), .ZN(new_n1070));
  XOR2_X1   g0870(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1071));
  XNOR2_X1  g0871(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  XOR2_X1   g0872(.A(KEYINPUT54), .B(G143), .Z(new_n1073));
  AOI211_X1 g0873(.A(new_n1069), .B(new_n1072), .C1(new_n781), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n770), .A2(G125), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1068), .B(new_n1076), .C1(G132), .C2(new_n788), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1031), .B1(new_n755), .B2(G107), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n772), .B2(new_n783), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n799), .B1(new_n457), .B2(new_n753), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n270), .B1(new_n787), .B2(G87), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(KEYINPUT117), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(KEYINPUT117), .B2(new_n1081), .C1(new_n498), .C2(new_n735), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1079), .B(new_n1083), .C1(G116), .C2(new_n788), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n726), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n804), .A2(new_n255), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n715), .A3(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT118), .Z(new_n1088));
  AOI22_X1  g0888(.A1(new_n1064), .A2(new_n714), .B1(new_n1065), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1064), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n705), .A2(new_n421), .A3(G330), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n613), .A2(new_n871), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1059), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1055), .A2(new_n874), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1093), .B1(new_n1094), .B2(new_n1063), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n703), .A2(G330), .A3(new_n704), .A4(new_n811), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n874), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1052), .A2(new_n810), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n874), .C2(new_n1055), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1092), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1090), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g0902(.A1(new_n1064), .A2(KEYINPUT114), .A3(new_n1100), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT114), .B1(new_n1064), .B2(new_n1100), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n660), .B(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT115), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1089), .B1(new_n1107), .B2(new_n1108), .ZN(G378));
  INV_X1    g0909(.A(new_n1092), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n851), .A2(new_n866), .A3(G330), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n893), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n851), .A2(new_n866), .A3(G330), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n891), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1114), .A2(new_n886), .A3(new_n1116), .A4(new_n885), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n637), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n266), .A2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n297), .B(new_n1120), .Z(new_n1121));
  INV_X1    g0921(.A(KEYINPUT55), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1123), .A2(KEYINPUT56), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT56), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1113), .A2(new_n1117), .A3(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1111), .A2(KEYINPUT57), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT57), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1104), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1064), .A2(new_n1100), .A3(KEYINPUT114), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1092), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1131), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT121), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1111), .A2(new_n1140), .A3(new_n1131), .A4(KEYINPUT57), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1133), .A2(new_n660), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n726), .A2(G50), .A3(new_n723), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n274), .A2(new_n275), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n770), .A2(G124), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G128), .A2(new_n788), .B1(new_n781), .B2(G137), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n800), .A2(G150), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n787), .A2(new_n1073), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n755), .A2(G132), .B1(new_n746), .B2(G125), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1145), .B(new_n1146), .C1(KEYINPUT59), .C2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(KEYINPUT59), .B2(new_n1151), .C1(new_n736), .C2(new_n740), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n345), .A2(new_n275), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1145), .A2(new_n259), .A3(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n752), .A2(new_n478), .B1(new_n740), .B2(new_n220), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n770), .B2(G283), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n756), .A2(new_n457), .B1(new_n783), .B2(new_n209), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1158), .A2(new_n965), .A3(new_n987), .A4(new_n1154), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(new_n356), .C2(new_n753), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT58), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1153), .A2(new_n1155), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n726), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n715), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1143), .B(new_n1164), .C1(new_n1127), .C2(new_n723), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1131), .B2(new_n714), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(new_n1166), .B(KEYINPUT120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1142), .A2(new_n1167), .ZN(G375));
  NAND3_X1  g0968(.A1(new_n874), .A2(KEYINPUT122), .A3(new_n723), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT122), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n849), .B2(new_n724), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n749), .A2(new_n736), .B1(new_n753), .B2(new_n251), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n770), .B2(G128), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n270), .B1(new_n740), .B2(new_n220), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT124), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n788), .A2(G137), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n783), .A2(new_n795), .B1(new_n743), .B2(new_n259), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n755), .B2(new_n1073), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1173), .A2(new_n1175), .A3(new_n1176), .A4(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n755), .A2(G116), .B1(new_n746), .B2(G294), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n478), .B2(new_n753), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n1181), .B(KEYINPUT123), .Z(new_n1182));
  OAI21_X1  g0982(.A(new_n345), .B1(new_n740), .B2(new_n202), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1183), .B(new_n990), .C1(G97), .C2(new_n787), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(new_n763), .C2(new_n735), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n752), .A2(new_n772), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1187), .A2(new_n726), .B1(new_n201), .B2(new_n804), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1169), .A2(new_n1171), .A3(new_n715), .A4(new_n1188), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n713), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1095), .A2(new_n1092), .A3(new_n1099), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n929), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1100), .B2(new_n1194), .ZN(G381));
  OR2_X1    g0995(.A1(G393), .A2(G396), .ZN(new_n1196));
  NOR4_X1   g0996(.A1(G387), .A2(G384), .A3(G390), .A4(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(G375), .ZN(new_n1198));
  INV_X1    g0998(.A(G381), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1105), .A2(new_n1089), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(G407));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n638), .A3(new_n1200), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(G407), .A2(G213), .A3(new_n1202), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT125), .Z(G409));
  AOI21_X1  g1004(.A(G390), .B1(new_n951), .B2(new_n977), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(G393), .A2(G396), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n951), .A2(new_n977), .A3(G390), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n1196), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1196), .A2(new_n1207), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1208), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1205), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT60), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n661), .B1(new_n1193), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n1101), .C1(new_n1214), .C2(new_n1193), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1192), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(G384), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n638), .A2(G213), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1142), .A2(G378), .A3(new_n1167), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1111), .A2(new_n929), .A3(new_n1131), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n1166), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1200), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT126), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT126), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n1225), .A3(new_n1200), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1218), .B(new_n1219), .C1(new_n1220), .C2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT127), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT62), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1222), .A2(new_n1225), .A3(new_n1200), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1225), .B1(new_n1222), .B2(new_n1200), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1142), .A2(new_n1167), .A3(G378), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT127), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1235), .A2(new_n1236), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1229), .A2(new_n1230), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1219), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n638), .A2(G213), .A3(G2897), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1218), .B(new_n1240), .Z(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT61), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1228), .A2(KEYINPUT62), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1213), .B1(new_n1238), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1237), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1233), .A2(new_n1234), .B1(G213), .B2(new_n638), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1236), .B1(new_n1248), .B2(new_n1218), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1228), .A2(new_n1246), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(new_n1213), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1242), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1245), .A2(new_n1253), .ZN(G405));
  NAND2_X1  g1054(.A1(G375), .A2(new_n1200), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1234), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(new_n1218), .ZN(new_n1257));
  XNOR2_X1  g1057(.A(new_n1257), .B(new_n1213), .ZN(G402));
endmodule


