//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  XOR2_X1   g000(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT67), .A3(G116), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(new_n199), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n202), .A2(new_n192), .A3(new_n191), .A4(new_n194), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT68), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n209), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT64), .B1(new_n211), .B2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n212), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT1), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(KEYINPUT64), .A3(G143), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n217), .A2(new_n218), .A3(G128), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(KEYINPUT66), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n220), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(G137), .ZN(new_n230));
  INV_X1    g044(.A(G137), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT11), .A3(G134), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(G137), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n230), .A2(new_n232), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n238), .B2(G131), .ZN(new_n239));
  AOI211_X1 g053(.A(KEYINPUT65), .B(new_n233), .C1(new_n234), .C2(new_n237), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n227), .A2(new_n235), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(new_n221), .B2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n221), .A2(G146), .ZN(new_n245));
  OAI211_X1 g059(.A(G128), .B(new_n219), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n225), .A2(new_n210), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT0), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT0), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(new_n214), .B2(new_n210), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n230), .A2(new_n234), .A3(new_n232), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n248), .A2(new_n250), .B1(new_n252), .B2(new_n235), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n208), .B1(new_n242), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n250), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n252), .A2(KEYINPUT69), .A3(new_n235), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT69), .B1(new_n252), .B2(new_n235), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n227), .A2(new_n235), .A3(new_n241), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n206), .A2(new_n207), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n188), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(G237), .A2(G953), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G210), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n266), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT70), .ZN(new_n270));
  OR3_X1    g084(.A1(new_n262), .A2(new_n264), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n273), .B1(new_n242), .B2(new_n253), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n258), .A2(KEYINPUT30), .A3(new_n259), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n208), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n261), .ZN(new_n277));
  INV_X1    g091(.A(new_n269), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n272), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n264), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n258), .A2(new_n259), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n208), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n261), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n287), .B2(new_n263), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n269), .A2(KEYINPUT29), .ZN(new_n289));
  OAI221_X1 g103(.A(new_n282), .B1(new_n281), .B2(new_n280), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n276), .A2(new_n261), .A3(new_n269), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT31), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n276), .A2(new_n294), .A3(new_n261), .A4(new_n269), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n270), .B1(new_n262), .B2(new_n264), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT72), .B(new_n270), .C1(new_n262), .C2(new_n264), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n296), .A2(KEYINPUT73), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n299), .A2(new_n295), .A3(new_n293), .A4(new_n300), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G472), .A2(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT32), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n301), .A2(new_n304), .A3(new_n308), .A4(new_n305), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n307), .A2(new_n309), .B1(KEYINPUT74), .B2(new_n306), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n291), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT92), .ZN(new_n314));
  INV_X1    g128(.A(G469), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  INV_X1    g130(.A(G107), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G104), .ZN(new_n318));
  INV_X1    g132(.A(G104), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G107), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G101), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT82), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n319), .A2(KEYINPUT3), .A3(G107), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g139(.A(G101), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .A4(new_n320), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT82), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n321), .A2(new_n328), .A3(G101), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n323), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(new_n227), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n217), .A2(new_n219), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n220), .B1(new_n332), .B2(new_n213), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n331), .A2(new_n334), .B1(new_n252), .B2(new_n235), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT12), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n256), .A2(new_n257), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n331), .B2(new_n334), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(KEYINPUT12), .B2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n324), .A2(new_n325), .A3(new_n320), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G101), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT4), .A3(new_n327), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n345), .A3(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n255), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n330), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n341), .A2(new_n337), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G140), .ZN(new_n350));
  INV_X1    g164(.A(G227), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G953), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n350), .B(new_n352), .Z(new_n353));
  AND2_X1   g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n339), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n341), .A2(new_n347), .A3(new_n348), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n256), .B2(new_n257), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n353), .B1(new_n357), .B2(new_n349), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n315), .B(new_n316), .C1(new_n355), .C2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n339), .A2(new_n349), .ZN(new_n360));
  INV_X1    g174(.A(new_n353), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n354), .A2(new_n357), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(G469), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n315), .A2(new_n316), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G221), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT9), .B(G234), .Z(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n316), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n369), .ZN(new_n373));
  INV_X1    g187(.A(G217), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n373), .A2(new_n374), .A3(G953), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n210), .A2(G143), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT88), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n221), .A2(G128), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(KEYINPUT89), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT89), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n229), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n378), .A2(new_n379), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(G134), .A3(new_n380), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G116), .B(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n317), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n190), .A2(KEYINPUT14), .A3(G122), .ZN(new_n391));
  INV_X1    g205(.A(new_n389), .ZN(new_n392));
  OAI211_X1 g206(.A(G107), .B(new_n391), .C1(new_n392), .C2(KEYINPUT14), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n388), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(G134), .B1(new_n386), .B2(new_n380), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n379), .B(KEYINPUT13), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n229), .B1(new_n378), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n389), .B(G107), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n376), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n388), .A2(new_n390), .A3(new_n393), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n375), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(KEYINPUT90), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT90), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n401), .A2(new_n402), .A3(new_n405), .A4(new_n375), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n316), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n407), .B(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n372), .A2(new_n411), .ZN(new_n412));
  OR2_X1    g226(.A1(KEYINPUT91), .A2(G952), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT91), .A2(G952), .ZN(new_n414));
  AOI21_X1  g228(.A(G953), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(G234), .A2(G237), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT21), .B(G898), .Z(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(G902), .A3(G953), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G214), .B1(G237), .B2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT83), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n227), .A2(G125), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n248), .A2(G125), .A3(new_n250), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n426), .A2(new_n424), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G953), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G224), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT84), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(KEYINPUT7), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n427), .B2(new_n428), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n193), .A3(G116), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n195), .B2(new_n436), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n203), .B1(new_n438), .B2(new_n196), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n323), .A2(new_n327), .A3(new_n329), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  XOR2_X1   g255(.A(G110), .B(G122), .Z(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT8), .Z(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n439), .A2(new_n440), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n206), .A2(new_n344), .A3(new_n207), .A4(new_n346), .ZN(new_n446));
  INV_X1    g260(.A(new_n442), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n433), .A2(new_n435), .A3(new_n444), .A4(new_n448), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n427), .A2(new_n432), .A3(new_n428), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n446), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n442), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT6), .A3(new_n448), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n432), .B1(new_n427), .B2(new_n428), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n455), .A3(new_n442), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n450), .A2(new_n453), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n457), .A3(new_n316), .ZN(new_n458));
  OAI21_X1  g272(.A(G210), .B1(G237), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n449), .A2(new_n457), .A3(new_n316), .A4(new_n459), .ZN(new_n462));
  AOI211_X1 g276(.A(new_n421), .B(new_n423), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n265), .A2(G214), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(G143), .ZN(new_n465));
  NAND2_X1  g279(.A1(KEYINPUT18), .A2(G131), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G125), .ZN(new_n469));
  INV_X1    g283(.A(G140), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G140), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(G140), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT79), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n472), .A2(G140), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n480));
  OAI21_X1  g294(.A(G125), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT79), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n477), .A2(new_n478), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n478), .B1(new_n477), .B2(new_n483), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n484), .A2(new_n485), .A3(new_n211), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n470), .A2(G125), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n487), .A2(new_n475), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n211), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT80), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT86), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n477), .A2(new_n483), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT85), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n477), .A2(new_n483), .A3(new_n478), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(G146), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT86), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n490), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n468), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT16), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n487), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n493), .B2(KEYINPUT16), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n503), .A2(new_n211), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n465), .A2(new_n505), .A3(new_n233), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n465), .B(G131), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n505), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n503), .A2(new_n211), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G113), .B(G122), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n319), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n499), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n496), .A2(new_n497), .A3(new_n490), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n497), .B1(new_n496), .B2(new_n490), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n467), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n513), .B1(new_n518), .B2(new_n510), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n316), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G475), .ZN(new_n521));
  INV_X1    g335(.A(G475), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n465), .B(new_n233), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n488), .A2(KEYINPUT19), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n494), .A2(new_n495), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n524), .B1(new_n525), .B2(KEYINPUT19), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n504), .B(new_n523), .C1(new_n526), .C2(G146), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n513), .B1(new_n518), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n522), .B(new_n316), .C1(new_n515), .C2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT87), .B1(new_n529), .B2(KEYINPUT20), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(KEYINPUT20), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n529), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n463), .B(new_n521), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n314), .B1(new_n412), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n504), .A2(new_n509), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n193), .A2(G128), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT77), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(KEYINPUT23), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT23), .B1(new_n210), .B2(G119), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n193), .B2(G128), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G110), .ZN(new_n543));
  XNOR2_X1  g357(.A(G119), .B(G128), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT76), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT24), .B(G110), .Z(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n536), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  OAI22_X1  g362(.A1(new_n545), .A2(new_n546), .B1(new_n542), .B2(G110), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n504), .A2(new_n549), .A3(new_n490), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT22), .B(G137), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n430), .A2(G221), .A3(G234), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n551), .B(new_n552), .Z(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n548), .B2(new_n550), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT81), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT25), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n559), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n557), .A2(new_n316), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n556), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n564), .A2(new_n316), .A3(new_n562), .A4(new_n554), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n560), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n374), .B1(G234), .B2(new_n316), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(G902), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n557), .A2(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n411), .A2(new_n367), .A3(new_n371), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n523), .B1(new_n503), .B2(new_n211), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT19), .B1(new_n484), .B2(new_n485), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n574), .B1(KEYINPUT19), .B2(new_n488), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n575), .B2(new_n211), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n514), .B1(new_n499), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n518), .A2(new_n513), .A3(new_n510), .ZN(new_n578));
  AOI21_X1  g392(.A(G475), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT20), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n316), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n579), .B2(new_n316), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n582), .B2(KEYINPUT87), .ZN(new_n583));
  OR3_X1    g397(.A1(new_n529), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n583), .A2(new_n584), .B1(G475), .B2(new_n520), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n572), .A2(new_n585), .A3(KEYINPUT92), .A4(new_n463), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n313), .A2(new_n535), .A3(new_n571), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  NAND2_X1  g402(.A1(new_n571), .A2(new_n372), .ZN(new_n589));
  INV_X1    g403(.A(new_n463), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n301), .A2(new_n304), .A3(new_n316), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n306), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n521), .B1(new_n532), .B2(new_n533), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n404), .A2(new_n596), .A3(new_n406), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n400), .A2(KEYINPUT33), .A3(new_n403), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n408), .A2(G902), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT93), .B(G478), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n599), .A2(new_n600), .B1(new_n407), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n594), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  NOR2_X1   g422(.A1(new_n531), .A2(new_n582), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n520), .A2(new_n610), .A3(G475), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n514), .B1(new_n499), .B2(new_n511), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n612), .B2(new_n578), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT94), .B1(new_n613), .B2(new_n522), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n609), .A2(new_n411), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n594), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT35), .B(G107), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  NAND2_X1  g433(.A1(new_n548), .A2(new_n550), .ZN(new_n620));
  INV_X1    g434(.A(new_n553), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n620), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n569), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n568), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n593), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n535), .A2(new_n586), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT37), .B(G110), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT95), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n628), .B(new_n630), .ZN(G12));
  NAND2_X1  g445(.A1(new_n461), .A2(new_n462), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n422), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n417), .B1(G900), .B2(new_n419), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n616), .A2(KEYINPUT96), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT96), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n611), .A2(new_n614), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n407), .B(new_n409), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n529), .A2(KEYINPUT20), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n581), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n638), .A2(new_n639), .A3(new_n641), .A4(new_n635), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n637), .B1(new_n642), .B2(new_n633), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n313), .A3(new_n372), .A4(new_n625), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  NAND2_X1  g460(.A1(new_n595), .A2(new_n639), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n632), .B(KEYINPUT38), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n635), .B(KEYINPUT39), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n372), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT40), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n422), .B(new_n648), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n647), .B(new_n653), .C1(new_n652), .C2(new_n651), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n307), .A2(new_n309), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n306), .A2(KEYINPUT74), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n311), .ZN(new_n658));
  INV_X1    g472(.A(G472), .ZN(new_n659));
  INV_X1    g473(.A(new_n270), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n292), .B1(new_n287), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n659), .B1(new_n661), .B2(new_n316), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n654), .A2(new_n626), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT97), .B(G143), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G45));
  AOI21_X1  g481(.A(new_n626), .B1(new_n658), .B2(new_n291), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n595), .A2(new_n634), .A3(new_n603), .A4(new_n635), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT98), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n668), .A2(new_n672), .A3(new_n372), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  AOI21_X1  g489(.A(new_n358), .B1(new_n339), .B2(new_n354), .ZN(new_n676));
  OAI21_X1  g490(.A(G469), .B1(new_n676), .B2(G902), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n677), .A2(new_n359), .A3(new_n371), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n463), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n313), .A2(new_n571), .A3(new_n605), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  AND2_X1   g497(.A1(new_n680), .A2(new_n616), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n313), .A2(new_n684), .A3(new_n571), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NOR3_X1   g500(.A1(new_n595), .A2(new_n679), .A3(new_n639), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n313), .A2(new_n625), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  AOI21_X1  g503(.A(new_n660), .B1(new_n288), .B2(KEYINPUT99), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(KEYINPUT99), .B2(new_n288), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n296), .ZN(new_n692));
  AOI22_X1  g506(.A1(new_n591), .A2(G472), .B1(new_n692), .B2(new_n305), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n571), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n639), .A3(new_n595), .A4(new_n680), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G122), .ZN(G24));
  INV_X1    g510(.A(new_n669), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n693), .A2(new_n625), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n678), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G125), .ZN(G27));
  INV_X1    g514(.A(new_n635), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n461), .A2(new_n422), .A3(new_n462), .ZN(new_n702));
  NOR4_X1   g516(.A1(new_n585), .A2(new_n602), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n364), .A2(KEYINPUT100), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n364), .A2(KEYINPUT100), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n359), .A3(new_n366), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n371), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n313), .A2(new_n571), .A3(new_n703), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT101), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n711));
  INV_X1    g525(.A(new_n702), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n595), .A2(new_n603), .A3(new_n635), .A4(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n707), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n313), .A4(new_n571), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n655), .A2(new_n291), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n718), .A2(new_n719), .A3(new_n571), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n719), .B1(new_n718), .B2(new_n571), .ZN(new_n721));
  OAI211_X1 g535(.A(KEYINPUT42), .B(new_n714), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G131), .ZN(G33));
  INV_X1    g538(.A(new_n642), .ZN(new_n725));
  AND4_X1   g539(.A1(new_n313), .A2(new_n571), .A3(new_n725), .A4(new_n712), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n708), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G134), .ZN(G36));
  AND2_X1   g542(.A1(new_n585), .A2(KEYINPUT105), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n585), .A2(KEYINPUT105), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n729), .A2(new_n730), .A3(new_n602), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT43), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT104), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n585), .B1(new_n603), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n733), .B2(new_n603), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n732), .B1(KEYINPUT43), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(new_n593), .A3(new_n625), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n702), .B(KEYINPUT106), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n362), .A2(new_n363), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(G469), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT46), .B1(new_n745), .B2(new_n366), .ZN(new_n746));
  INV_X1    g560(.A(new_n359), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(KEYINPUT46), .A3(new_n366), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n370), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n650), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT103), .Z(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n738), .B2(new_n737), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n741), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g568(.A(KEYINPUT107), .B(G137), .Z(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(G39));
  XNOR2_X1  g570(.A(new_n750), .B(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n703), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n313), .A3(new_n571), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n470), .ZN(G42));
  INV_X1    g574(.A(new_n664), .ZN(new_n761));
  INV_X1    g575(.A(new_n571), .ZN(new_n762));
  NOR4_X1   g576(.A1(new_n762), .A2(new_n648), .A3(new_n370), .A4(new_n423), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n677), .A2(new_n359), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n764), .B(KEYINPUT49), .Z(new_n765));
  NAND4_X1  g579(.A1(new_n761), .A2(new_n731), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT108), .Z(new_n767));
  AND3_X1   g581(.A1(new_n736), .A2(new_n416), .A3(new_n415), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n694), .A3(new_n740), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n764), .A2(new_n371), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n757), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n769), .A2(new_n770), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n768), .A2(new_n678), .A3(new_n694), .ZN(new_n776));
  INV_X1    g590(.A(new_n648), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n423), .A3(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n776), .A2(new_n423), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n702), .A2(new_n764), .A3(new_n370), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n761), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n762), .A2(new_n417), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n585), .A3(new_n602), .A4(new_n786), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n775), .A2(new_n780), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n768), .A2(new_n783), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n698), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n790), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n775), .A2(new_n780), .A3(new_n782), .A4(new_n787), .ZN(new_n796));
  INV_X1    g610(.A(new_n792), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g613(.A1(new_n784), .A2(new_n762), .A3(new_n417), .A4(new_n604), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n717), .A2(new_n722), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n681), .A2(new_n685), .A3(new_n688), .A4(new_n695), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n604), .B1(new_n411), .B2(new_n595), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n594), .A2(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n587), .A2(new_n628), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n609), .A2(new_n615), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n313), .A2(new_n572), .A3(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n605), .A2(new_n693), .A3(new_n708), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n626), .A2(new_n701), .A3(new_n702), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n803), .A2(new_n806), .A3(new_n812), .A4(new_n727), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n801), .B1(new_n802), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n673), .A2(new_n313), .A3(new_n372), .A4(new_n625), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n645), .B(new_n699), .C1(new_n816), .C2(new_n671), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n647), .A2(new_n707), .A3(new_n633), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n664), .A2(new_n626), .A3(new_n635), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n815), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n645), .A2(new_n699), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(KEYINPUT52), .A3(new_n674), .A4(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n810), .A2(new_n811), .B1(new_n726), .B2(new_n708), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n681), .A2(new_n685), .A3(new_n688), .A4(new_n695), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n587), .A2(new_n628), .A3(new_n805), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n723), .A2(KEYINPUT109), .A3(new_n825), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n814), .A2(new_n824), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  INV_X1    g647(.A(new_n813), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n824), .A2(new_n834), .A3(KEYINPUT53), .A4(new_n723), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n824), .A4(new_n829), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n833), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT110), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n832), .A2(new_n837), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT54), .ZN(new_n841));
  AND4_X1   g655(.A1(KEYINPUT53), .A2(new_n824), .A3(new_n834), .A4(new_n723), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n831), .B2(new_n830), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n833), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT110), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n839), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n791), .B1(new_n720), .B2(new_n721), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT48), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n776), .A2(new_n634), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n849), .A2(new_n415), .A3(new_n850), .ZN(new_n851));
  NOR4_X1   g665(.A1(new_n799), .A2(new_n800), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(G952), .A2(G953), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT114), .Z(new_n854));
  OAI21_X1  g668(.A(new_n767), .B1(new_n852), .B2(new_n854), .ZN(G75));
  NOR2_X1   g669(.A1(new_n843), .A2(new_n316), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT56), .B1(new_n856), .B2(G210), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n450), .A2(new_n454), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n453), .A2(new_n456), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n457), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT55), .ZN(new_n862));
  NOR2_X1   g676(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n857), .B(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n430), .A2(G952), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n865), .A2(new_n866), .ZN(G51));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT116), .B1(new_n843), .B2(new_n833), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n832), .A2(new_n835), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n872), .A3(new_n844), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n365), .B(KEYINPUT57), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n676), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI211_X1 g691(.A(KEYINPUT117), .B(new_n676), .C1(new_n873), .C2(new_n874), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n843), .A2(new_n316), .A3(new_n745), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n866), .B1(new_n879), .B2(new_n880), .ZN(G54));
  NAND3_X1  g695(.A1(new_n856), .A2(KEYINPUT58), .A3(G475), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n577), .A2(new_n578), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n882), .B(new_n883), .Z(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n866), .ZN(G60));
  XNOR2_X1  g699(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n408), .A2(new_n316), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n886), .B(new_n887), .Z(new_n888));
  NAND2_X1  g702(.A1(new_n847), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n599), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n866), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n873), .A2(new_n599), .A3(new_n888), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n888), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n839), .B2(new_n846), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n892), .B(new_n893), .C1(new_n896), .C2(new_n599), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n894), .A2(new_n899), .ZN(G63));
  NOR2_X1   g714(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n901));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT60), .Z(new_n903));
  AOI21_X1  g717(.A(new_n557), .B1(new_n870), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n866), .ZN(new_n905));
  MUX2_X1   g719(.A(KEYINPUT121), .B(new_n901), .S(new_n905), .Z(new_n906));
  NAND3_X1  g720(.A1(new_n870), .A2(new_n623), .A3(new_n903), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT120), .Z(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n907), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n906), .A2(new_n908), .B1(KEYINPUT61), .B2(new_n909), .ZN(G66));
  XNOR2_X1  g724(.A(new_n828), .B(KEYINPUT122), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n430), .B1(new_n418), .B2(G224), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n912), .A2(new_n430), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT124), .Z(new_n917));
  OAI21_X1  g731(.A(new_n859), .B1(G898), .B2(new_n430), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  AOI21_X1  g733(.A(new_n759), .B1(new_n741), .B2(new_n753), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n720), .A2(new_n721), .ZN(new_n921));
  OR4_X1    g735(.A1(new_n633), .A2(new_n752), .A3(new_n647), .A4(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n817), .B(KEYINPUT125), .Z(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(new_n727), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n920), .A2(new_n922), .A3(new_n723), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n430), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n274), .A2(new_n275), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(new_n526), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n923), .A2(new_n665), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n762), .B1(new_n658), .B2(new_n291), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n934), .A2(new_n651), .A3(new_n712), .A4(new_n804), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n935), .A3(new_n920), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n928), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n430), .ZN(new_n939));
  INV_X1    g753(.A(G900), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n351), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n926), .A2(G900), .A3(new_n929), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n939), .A2(KEYINPUT126), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n945));
  AOI21_X1  g759(.A(G953), .B1(new_n930), .B2(new_n937), .ZN(new_n946));
  INV_X1    g760(.A(new_n942), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n943), .A2(new_n948), .ZN(G72));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT63), .Z(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n936), .B2(new_n912), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n277), .B(KEYINPUT127), .Z(new_n953));
  NAND3_X1  g767(.A1(new_n952), .A2(new_n269), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n279), .A2(new_n292), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n840), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n951), .B1(new_n925), .B2(new_n912), .ZN(new_n957));
  INV_X1    g771(.A(new_n953), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n278), .A3(new_n958), .ZN(new_n959));
  AND4_X1   g773(.A1(new_n892), .A2(new_n954), .A3(new_n956), .A4(new_n959), .ZN(G57));
endmodule


