//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(G1gat), .ZN(new_n209));
  OAI21_X1  g008(.A(G8gat), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(new_n211), .C1(G1gat), .C2(new_n205), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n214));
  INV_X1    g013(.A(G57gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G64gat), .ZN(new_n216));
  INV_X1    g015(.A(G64gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G57gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT93), .ZN(new_n220));
  NAND2_X1  g019(.A1(G71gat), .A2(G78gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G71gat), .A2(G78gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(G71gat), .A2(G78gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT93), .A3(new_n221), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n219), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT92), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(KEYINPUT92), .A2(G71gat), .A3(G78gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G57gat), .B(G64gat), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n231), .B(new_n225), .C1(new_n232), .C2(new_n214), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT94), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT94), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n227), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n213), .B1(new_n238), .B2(KEYINPUT21), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G183gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G183gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n239), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n242), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n204), .B1(new_n243), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n250));
  NAND2_X1  g049(.A1(G231gat), .A2(G233gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  NAND3_X1  g051(.A1(new_n243), .A2(new_n247), .A3(new_n204), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n249), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n252), .ZN(new_n255));
  INV_X1    g054(.A(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(G29gat), .A2(G36gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT14), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G29gat), .A2(G36gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G43gat), .B(G50gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT15), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G43gat), .B(G50gat), .Z(new_n269));
  INV_X1    g068(.A(KEYINPUT15), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT88), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n263), .B(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n271), .A2(new_n262), .A3(new_n266), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT17), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT17), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n268), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G99gat), .ZN(new_n280));
  INV_X1    g079(.A(G106gat), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT8), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT96), .B(G92gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(G85gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(G85gat), .A2(G92gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT7), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G99gat), .B(G106gat), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n288), .A2(KEYINPUT97), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n284), .B2(new_n287), .ZN(new_n292));
  XOR2_X1   g091(.A(KEYINPUT96), .B(G92gat), .Z(new_n293));
  INV_X1    g092(.A(G85gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n285), .B(KEYINPUT7), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n295), .A2(new_n290), .A3(new_n282), .A4(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT97), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n279), .A2(new_n291), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n291), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n275), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G134gat), .B(G162gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G190gat), .B(G218gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT98), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n308), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n259), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n317), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT23), .ZN(new_n320));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n318), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT24), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n328), .A2(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n324), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n244), .A2(KEYINPUT66), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT66), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G183gat), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n329), .B(new_n327), .C1(new_n339), .C2(G190gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(KEYINPUT25), .A3(new_n324), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n343));
  OR2_X1    g142(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n345));
  AOI21_X1  g144(.A(G190gat), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT28), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n325), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT27), .ZN(new_n349));
  AOI21_X1  g148(.A(G190gat), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(KEYINPUT67), .B(new_n319), .C1(new_n318), .C2(KEYINPUT26), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n319), .A2(KEYINPUT26), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(new_n321), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n343), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n349), .A2(new_n344), .ZN(new_n359));
  INV_X1    g158(.A(G190gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n359), .A2(new_n347), .A3(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT27), .B(G183gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n360), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n326), .B1(new_n363), .B2(KEYINPUT28), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n361), .A2(new_n364), .A3(new_n357), .A4(new_n343), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n342), .B1(new_n358), .B2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G127gat), .B(G134gat), .Z(new_n368));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n368), .B1(KEYINPUT1), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT69), .ZN(new_n371));
  INV_X1    g170(.A(G120gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(G113gat), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n374), .A2(G120gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n368), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT1), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n373), .B2(new_n375), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(new_n377), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n370), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n367), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n361), .A2(new_n364), .A3(new_n357), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT68), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n390), .A2(new_n365), .B1(new_n335), .B2(new_n341), .ZN(new_n391));
  INV_X1    g190(.A(new_n386), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(new_n388), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n395));
  NOR2_X1   g194(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT73), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT73), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n394), .A2(new_n400), .A3(new_n395), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G71gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(new_n280), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT71), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT33), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n406), .B2(new_n405), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n393), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n388), .B(KEYINPUT64), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI221_X4 g210(.A(new_n386), .B1(new_n335), .B2(new_n341), .C1(new_n390), .C2(new_n365), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n365), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n392), .B1(new_n413), .B2(new_n342), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n410), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(KEYINPUT32), .A2(new_n411), .B1(new_n419), .B2(new_n405), .ZN(new_n420));
  OR3_X1    g219(.A1(new_n409), .A2(KEYINPUT34), .A3(new_n410), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n402), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n402), .B2(new_n421), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(G211gat), .A2(G218gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(G211gat), .A2(G218gat), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT75), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(G211gat), .ZN(new_n428));
  INV_X1    g227(.A(G218gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT75), .ZN(new_n431));
  NAND2_X1  g230(.A1(G211gat), .A2(G218gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT74), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT22), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G197gat), .B(G204gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT29), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n427), .A2(new_n433), .A3(new_n439), .A4(new_n440), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT3), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G155gat), .ZN(new_n448));
  INV_X1    g247(.A(G162gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR3_X1   g249(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n451));
  INV_X1    g250(.A(G141gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(G148gat), .ZN(new_n453));
  INV_X1    g252(.A(G148gat), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n454), .A2(G141gat), .ZN(new_n455));
  OAI22_X1  g254(.A1(new_n450), .A2(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n450), .ZN(new_n457));
  XNOR2_X1  g256(.A(G141gat), .B(G148gat), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n457), .B1(new_n458), .B2(KEYINPUT2), .ZN(new_n459));
  NOR2_X1   g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT79), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n456), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n446), .B(new_n456), .C1(new_n459), .C2(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n443), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT76), .ZN(new_n466));
  AND4_X1   g265(.A1(new_n427), .A2(new_n433), .A3(new_n439), .A4(new_n440), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n427), .A2(new_n433), .B1(new_n439), .B2(new_n440), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n442), .A2(KEYINPUT76), .A3(new_n444), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G228gat), .ZN(new_n472));
  INV_X1    g271(.A(G233gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n463), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n463), .A2(new_n471), .A3(new_n477), .A4(new_n474), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n467), .A2(new_n468), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n443), .B2(new_n464), .ZN(new_n481));
  INV_X1    g280(.A(new_n451), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n458), .B1(new_n457), .B2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G141gat), .B(G148gat), .Z(new_n484));
  INV_X1    g283(.A(KEYINPUT2), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n450), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n461), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n445), .B2(new_n446), .ZN(new_n489));
  OAI22_X1  g288(.A1(new_n481), .A2(new_n489), .B1(new_n472), .B2(new_n473), .ZN(new_n490));
  INV_X1    g289(.A(G22gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT83), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n479), .A2(KEYINPUT84), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G78gat), .B(G106gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT31), .ZN(new_n496));
  INV_X1    g295(.A(G50gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n476), .A2(new_n491), .A3(new_n490), .A4(new_n478), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n476), .A2(new_n490), .A3(new_n478), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n492), .B1(new_n502), .B2(new_n500), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(G22gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n499), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n498), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT85), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n424), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT35), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(new_n386), .B2(new_n462), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n384), .A2(new_n377), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n368), .B1(new_n384), .B2(new_n377), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n383), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(new_n488), .A3(KEYINPUT4), .A4(new_n370), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n386), .A2(new_n523), .A3(new_n464), .ZN(new_n524));
  NAND2_X1  g323(.A1(G225gat), .A2(G233gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n522), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n386), .B2(new_n462), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n517), .A2(new_n529), .A3(new_n521), .A4(new_n524), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n386), .A2(new_n462), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n488), .B1(new_n520), .B2(new_n370), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n526), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT80), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT80), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n530), .A2(new_n533), .A3(new_n536), .A4(KEYINPUT5), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n528), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539));
  XOR2_X1   g338(.A(G1gat), .B(G29gat), .Z(new_n540));
  XNOR2_X1  g339(.A(G57gat), .B(G85gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  NOR3_X1   g343(.A1(new_n538), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n538), .A2(new_n544), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT6), .B1(new_n538), .B2(new_n544), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AND2_X1   g348(.A1(G226gat), .A2(G233gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(KEYINPUT29), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n367), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n469), .A2(new_n470), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n342), .A2(new_n550), .A3(new_n389), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n552), .A2(KEYINPUT77), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n551), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n553), .B(new_n554), .C1(new_n391), .C2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT77), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n413), .A2(new_n550), .A3(new_n342), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n556), .B1(new_n342), .B2(new_n389), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n480), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G8gat), .B(G36gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n217), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n555), .A2(new_n559), .A3(new_n562), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT30), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT78), .ZN(new_n571));
  INV_X1    g370(.A(new_n568), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT30), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n559), .A3(new_n562), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n566), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n568), .A2(new_n576), .A3(new_n569), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n571), .A2(new_n573), .A3(new_n575), .A4(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n549), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  INV_X1    g379(.A(new_n544), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n581), .B1(new_n538), .B2(KEYINPUT86), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT86), .ZN(new_n583));
  AOI211_X1 g382(.A(new_n583), .B(new_n528), .C1(new_n535), .C2(new_n537), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n548), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n545), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n424), .A2(new_n512), .A3(new_n580), .A4(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n515), .A2(new_n579), .B1(new_n514), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n582), .A2(new_n584), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n522), .A2(new_n524), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n526), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n544), .B1(new_n592), .B2(KEYINPUT39), .ZN(new_n593));
  OR3_X1    g392(.A1(new_n531), .A2(new_n532), .A3(new_n526), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(KEYINPUT39), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n596), .A2(KEYINPUT40), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(KEYINPUT40), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n578), .A2(new_n590), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n574), .A2(KEYINPUT37), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n555), .A2(new_n559), .A3(new_n562), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n566), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n572), .B1(new_n603), .B2(KEYINPUT38), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n560), .A2(new_n480), .A3(new_n561), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n553), .B1(new_n552), .B2(new_n554), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT37), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n607), .A2(new_n602), .A3(new_n608), .A4(new_n566), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n604), .A2(new_n585), .A3(new_n586), .A4(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n599), .A2(new_n610), .A3(new_n512), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n510), .B(new_n511), .C1(new_n549), .C2(new_n578), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n422), .B2(new_n423), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n412), .A2(new_n414), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n396), .B1(new_n615), .B2(new_n388), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n400), .B1(new_n616), .B2(new_n395), .ZN(new_n617));
  INV_X1    g416(.A(new_n401), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n421), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n420), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n402), .A2(new_n420), .A3(new_n421), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(KEYINPUT36), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n611), .A2(new_n612), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n315), .B1(new_n589), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G204gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G176gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT101), .Z(new_n631));
  NAND4_X1  g430(.A1(new_n299), .A2(new_n235), .A3(new_n291), .A4(new_n237), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n292), .A2(new_n297), .A3(new_n233), .A4(new_n227), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n302), .A2(KEYINPUT10), .A3(new_n238), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(KEYINPUT102), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n638), .B1(new_n632), .B2(new_n634), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n631), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n630), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n647), .B(new_n639), .C1(new_n646), .C2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n213), .ZN(new_n650));
  INV_X1    g449(.A(new_n278), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n277), .B1(new_n268), .B2(new_n274), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G229gat), .A2(G233gat), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n210), .A2(new_n212), .B1(new_n268), .B2(new_n274), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(KEYINPUT89), .A2(KEYINPUT18), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n653), .A2(new_n654), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(KEYINPUT89), .A2(KEYINPUT18), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n655), .B1(new_n279), .B2(new_n650), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n661), .A2(KEYINPUT89), .A3(KEYINPUT18), .A4(new_n654), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n213), .A2(new_n275), .A3(KEYINPUT90), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT90), .B1(new_n213), .B2(new_n275), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n656), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n654), .B(KEYINPUT13), .Z(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n660), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT12), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT11), .B(G169gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G197gat), .ZN(new_n671));
  XOR2_X1   g470(.A(G113gat), .B(G141gat), .Z(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT87), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n669), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n678), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n676), .A3(KEYINPUT12), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n660), .A2(new_n662), .A3(new_n667), .A4(new_n682), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(KEYINPUT91), .A3(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT91), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n668), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n649), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n626), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n549), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT103), .B(G1gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT104), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n693), .B(new_n695), .ZN(G1324gat));
  NOR2_X1   g495(.A1(new_n691), .A2(new_n580), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n206), .A2(new_n211), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n206), .A2(new_n211), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n703), .B(new_n704), .C1(new_n211), .C2(new_n697), .ZN(G1325gat));
  INV_X1    g504(.A(new_n691), .ZN(new_n706));
  INV_X1    g505(.A(new_n624), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n707), .A2(KEYINPUT105), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(KEYINPUT105), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  AND3_X1   g510(.A1(new_n706), .A2(G15gat), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(G15gat), .B1(new_n706), .B2(new_n424), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(G1326gat));
  NOR2_X1   g513(.A1(new_n691), .A2(new_n512), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT43), .B(G22gat), .Z(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  AOI21_X1  g516(.A(new_n314), .B1(new_n589), .B2(new_n625), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n690), .A2(new_n258), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n721), .A2(G29gat), .A3(new_n692), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT45), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n588), .A2(new_n514), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n579), .A2(KEYINPUT35), .A3(new_n512), .A4(new_n424), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n599), .A2(new_n610), .A3(new_n512), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n624), .A2(new_n612), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n724), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n313), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(KEYINPUT44), .A3(new_n313), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n720), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n692), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n723), .A2(new_n735), .ZN(G1328gat));
  NOR3_X1   g535(.A1(new_n721), .A2(G36gat), .A3(new_n580), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n734), .B2(new_n580), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(new_n424), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n721), .A2(G43gat), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n731), .A2(new_n707), .A3(new_n732), .A4(new_n720), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(KEYINPUT106), .ZN(new_n744));
  OAI21_X1  g543(.A(G43gat), .B1(new_n743), .B2(KEYINPUT106), .ZN(new_n745));
  OAI211_X1 g544(.A(KEYINPUT47), .B(new_n742), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n711), .A3(new_n732), .A4(new_n720), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G43gat), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n748), .A2(new_n742), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(KEYINPUT47), .B2(new_n749), .ZN(G1330gat));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n721), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n512), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n718), .A2(KEYINPUT107), .A3(new_n720), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n497), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n733), .A2(G50gat), .A3(new_n753), .A4(new_n720), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT48), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n760), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1331gat));
  INV_X1    g561(.A(new_n649), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n589), .B2(new_n625), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n686), .A2(new_n688), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n258), .A2(new_n313), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n549), .B(KEYINPUT108), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(new_n215), .ZN(G1332gat));
  INV_X1    g570(.A(new_n767), .ZN(new_n772));
  NAND2_X1  g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(new_n578), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n775));
  NOR2_X1   g574(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n774), .B(new_n777), .ZN(G1333gat));
  NAND3_X1  g577(.A1(new_n772), .A2(G71gat), .A3(new_n711), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n767), .A2(new_n741), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(G71gat), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n753), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g583(.A1(new_n259), .A2(new_n763), .A3(new_n765), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n733), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n786), .A2(new_n294), .A3(new_n692), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n259), .A2(new_n765), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT51), .B1(new_n718), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n728), .A2(KEYINPUT51), .A3(new_n313), .A4(new_n788), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n649), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n792), .A2(new_n692), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n787), .B1(new_n793), .B2(new_n294), .ZN(G1336gat));
  NAND4_X1  g593(.A1(new_n731), .A2(new_n578), .A3(new_n732), .A4(new_n785), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(new_n795), .B2(new_n283), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n578), .A2(new_n565), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n795), .A2(KEYINPUT111), .A3(new_n283), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT111), .B1(new_n795), .B2(new_n283), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n728), .A2(new_n313), .A3(new_n788), .ZN(new_n801));
  XNOR2_X1  g600(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n763), .B(new_n797), .C1(new_n803), .C2(new_n790), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n799), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n798), .B1(new_n805), .B2(new_n806), .ZN(G1337gat));
  XOR2_X1   g606(.A(KEYINPUT113), .B(G99gat), .Z(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n786), .B2(new_n710), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n741), .A2(new_n808), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n792), .B2(new_n810), .ZN(G1338gat));
  AOI21_X1  g610(.A(new_n763), .B1(new_n803), .B2(new_n790), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n512), .A2(G106gat), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n731), .A2(new_n753), .A3(new_n732), .A4(new_n785), .ZN(new_n814));
  XOR2_X1   g613(.A(KEYINPUT114), .B(G106gat), .Z(new_n815));
  AOI22_X1  g614(.A1(new_n812), .A2(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT115), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n812), .A2(new_n813), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n815), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n823));
  XNOR2_X1  g622(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n824));
  INV_X1    g623(.A(new_n813), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n820), .B(new_n824), .C1(new_n792), .C2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n818), .A2(new_n823), .A3(new_n826), .ZN(G1339gat));
  NAND4_X1  g626(.A1(new_n259), .A2(new_n314), .A3(new_n763), .A4(new_n689), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n635), .A2(G230gat), .A3(G233gat), .A4(new_n636), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n639), .A2(new_n830), .A3(KEYINPUT54), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n639), .A2(new_n830), .A3(KEYINPUT117), .A4(KEYINPUT54), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n640), .B2(new_n642), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n630), .A4(new_n837), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n648), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n673), .A2(new_n675), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n665), .A2(new_n666), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n661), .A2(new_n654), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n685), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n835), .A2(new_n630), .A3(new_n837), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n839), .A2(new_n313), .A3(new_n845), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n645), .B2(new_n648), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n689), .B1(new_n847), .B2(new_n846), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n839), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n852), .B2(new_n313), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n829), .B1(new_n853), .B2(new_n258), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n854), .A2(new_n578), .A3(new_n769), .ZN(new_n855));
  INV_X1    g654(.A(new_n513), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n374), .A3(new_n765), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n854), .A2(new_n513), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n549), .A3(new_n580), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n689), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(G1340gat));
  OAI21_X1  g662(.A(G120gat), .B1(new_n861), .B2(new_n763), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n649), .A2(new_n372), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n857), .B2(new_n865), .ZN(G1341gat));
  INV_X1    g665(.A(G127gat), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n861), .A2(new_n867), .A3(new_n258), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n858), .A2(new_n259), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(new_n867), .ZN(G1342gat));
  OR2_X1    g669(.A1(new_n314), .A2(G134gat), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n857), .A2(KEYINPUT56), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n861), .B2(new_n314), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT56), .B1(new_n857), .B2(new_n871), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  AOI21_X1  g674(.A(new_n512), .B1(new_n708), .B2(new_n709), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n855), .A2(new_n765), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n452), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(new_n852), .B2(new_n313), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n848), .A2(new_n765), .A3(new_n648), .A4(new_n838), .ZN(new_n881));
  INV_X1    g680(.A(new_n850), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(KEYINPUT118), .A3(new_n314), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n884), .A3(new_n849), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n829), .B1(new_n885), .B2(new_n258), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n512), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n707), .A2(new_n692), .A3(new_n578), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n883), .A2(new_n314), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n259), .B1(new_n890), .B2(new_n849), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n889), .B(new_n753), .C1(new_n891), .C2(new_n829), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n887), .A2(G141gat), .A3(new_n888), .A4(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n878), .B1(new_n893), .B2(new_n689), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT58), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g695(.A(KEYINPUT58), .B(new_n878), .C1(new_n893), .C2(new_n689), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1344gat));
  NAND4_X1  g697(.A1(new_n887), .A2(new_n649), .A3(new_n888), .A4(new_n892), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(G148gat), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT57), .B1(new_n854), .B2(new_n512), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n828), .A2(KEYINPUT119), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n766), .A2(new_n905), .A3(new_n763), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n889), .B(new_n753), .C1(new_n891), .C2(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n903), .A2(new_n908), .A3(new_n649), .A4(new_n888), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G148gat), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n902), .B1(new_n910), .B2(KEYINPUT59), .ZN(new_n911));
  AOI211_X1 g710(.A(KEYINPUT120), .B(new_n900), .C1(new_n909), .C2(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n855), .A2(new_n876), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n454), .A3(new_n649), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1345gat));
  AOI21_X1  g715(.A(G155gat), .B1(new_n914), .B2(new_n259), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n448), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n917), .B1(new_n919), .B2(new_n259), .ZN(G1346gat));
  AOI21_X1  g719(.A(G162gat), .B1(new_n914), .B2(new_n313), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n918), .A2(new_n449), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n313), .ZN(G1347gat));
  NOR4_X1   g722(.A1(new_n854), .A2(new_n549), .A3(new_n580), .A4(new_n513), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n316), .A3(new_n765), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n768), .A2(new_n580), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n860), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(new_n765), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(new_n316), .ZN(G1348gat));
  AOI21_X1  g728(.A(G176gat), .B1(new_n924), .B2(new_n649), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n763), .A2(new_n317), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n927), .B2(new_n931), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n860), .A2(new_n259), .A3(new_n926), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT121), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n860), .A2(new_n935), .A3(new_n259), .A4(new_n926), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n339), .A3(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT60), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n259), .A3(new_n362), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n937), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1350gat));
  NAND3_X1  g742(.A1(new_n924), .A2(new_n360), .A3(new_n313), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT123), .Z(new_n945));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n313), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n947), .B2(G190gat), .ZN(new_n948));
  AOI211_X1 g747(.A(KEYINPUT61), .B(new_n360), .C1(new_n927), .C2(new_n313), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G1351gat));
  AND2_X1   g749(.A1(new_n903), .A2(new_n908), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n710), .A3(new_n926), .ZN(new_n952));
  OAI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n689), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n854), .A2(new_n549), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n578), .A3(new_n876), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n955), .A2(G197gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n689), .B2(new_n956), .ZN(G1352gat));
  NOR2_X1   g756(.A1(new_n763), .A2(G204gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n954), .A2(new_n578), .A3(new_n876), .A4(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n951), .A2(new_n649), .A3(new_n710), .A4(new_n926), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(G204gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n962), .A2(new_n964), .A3(new_n967), .ZN(G1353gat));
  OR3_X1    g767(.A1(new_n955), .A2(G211gat), .A3(new_n258), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n951), .A2(new_n259), .A3(new_n710), .A4(new_n926), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  OAI21_X1  g772(.A(new_n429), .B1(new_n955), .B2(new_n314), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT126), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n976), .B(new_n429), .C1(new_n955), .C2(new_n314), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n951), .A2(new_n979), .A3(new_n710), .A4(new_n926), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(G218gat), .A3(new_n313), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n952), .A2(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1355gat));
endmodule


