//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G902), .ZN(new_n193));
  AOI211_X1 g007(.A(new_n193), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT21), .B(G898), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT1), .B1(new_n197), .B2(G146), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n197), .A2(G146), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  OAI211_X1 g015(.A(G128), .B(new_n198), .C1(new_n199), .C2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n203), .B(new_n204), .C1(KEYINPUT1), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n203), .A2(new_n204), .A3(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(G143), .B(G146), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT0), .B(G128), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G224), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G953), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n218), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n209), .A2(new_n220), .A3(new_n215), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n224));
  INV_X1    g038(.A(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G107), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT3), .A3(G104), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(G107), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT79), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G101), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n226), .A2(new_n228), .B1(new_n225), .B2(G107), .ZN(new_n234));
  INV_X1    g048(.A(G101), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT79), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT80), .B(G101), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n237), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n233), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n243), .A3(new_n244), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G116), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G116), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(new_n256), .A3(G119), .ZN(new_n257));
  INV_X1    g071(.A(G119), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G116), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n247), .A2(new_n251), .B1(new_n257), .B2(new_n259), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n231), .A2(G101), .ZN(new_n263));
  OAI22_X1  g077(.A1(new_n261), .A2(new_n262), .B1(new_n263), .B2(KEYINPUT4), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n259), .B2(KEYINPUT5), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n267), .A2(new_n258), .A3(KEYINPUT84), .A4(G116), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n266), .A2(G113), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n257), .A2(KEYINPUT5), .A3(new_n259), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n257), .A2(new_n259), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n245), .A2(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT81), .B1(new_n227), .B2(G104), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n225), .A3(G107), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n227), .A2(G104), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G101), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n234), .A2(new_n238), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(KEYINPUT82), .A3(G101), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  OAI22_X1  g100(.A1(new_n241), .A2(new_n264), .B1(new_n275), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(G110), .B(G122), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT86), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n252), .A2(new_n260), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n234), .A2(new_n235), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n274), .A2(new_n291), .B1(new_n292), .B2(new_n237), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n240), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n269), .A2(new_n270), .B1(new_n272), .B2(new_n273), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(new_n283), .A3(new_n284), .A4(new_n285), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n294), .A2(new_n296), .A3(new_n297), .A4(new_n288), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n290), .A2(KEYINPUT6), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT85), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT6), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n286), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n304), .A2(new_n295), .B1(new_n293), .B2(new_n240), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n305), .B2(new_n288), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n287), .A2(new_n289), .A3(new_n302), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n223), .B1(new_n299), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G210), .B1(G237), .B2(G902), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n290), .A2(new_n298), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT7), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n220), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n219), .A2(new_n221), .A3(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n209), .A2(new_n312), .A3(new_n220), .A4(new_n215), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n270), .A2(KEYINPUT87), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n269), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n270), .A2(KEYINPUT87), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n274), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n304), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n288), .B(KEYINPUT8), .Z(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n286), .B2(new_n295), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n314), .A2(new_n315), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n311), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n309), .A2(new_n310), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(new_n310), .ZN(new_n326));
  AOI211_X1 g140(.A(new_n288), .B(new_n303), .C1(new_n294), .C2(new_n296), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n302), .B1(new_n287), .B2(new_n289), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n290), .A2(KEYINPUT6), .A3(new_n298), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n222), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n297), .B1(new_n305), .B2(new_n288), .ZN(new_n332));
  INV_X1    g146(.A(new_n298), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n323), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n193), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n326), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G214), .B1(G237), .B2(G902), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT88), .ZN(new_n340));
  INV_X1    g154(.A(new_n338), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n325), .B2(new_n336), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT88), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n196), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G469), .ZN(new_n346));
  XNOR2_X1  g160(.A(G110), .B(G140), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n187), .A2(G227), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G137), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G134), .ZN(new_n352));
  INV_X1    g166(.A(G134), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT11), .B1(new_n353), .B2(G137), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT11), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n351), .A3(G134), .ZN(new_n356));
  AOI211_X1 g170(.A(G131), .B(new_n352), .C1(new_n354), .C2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G131), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n354), .A2(new_n356), .ZN(new_n359));
  INV_X1    g173(.A(new_n352), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n214), .B1(new_n292), .B2(new_n237), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n240), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT69), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n207), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n202), .A2(KEYINPUT69), .A3(new_n206), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(KEYINPUT10), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n286), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n207), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(new_n283), .A3(new_n284), .A4(new_n285), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n363), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(KEYINPUT83), .B(new_n363), .C1(new_n370), .C2(new_n375), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n202), .A2(KEYINPUT69), .A3(new_n206), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT69), .B1(new_n202), .B2(new_n206), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n383), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n384), .A2(new_n362), .A3(new_n374), .A4(new_n365), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n350), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n286), .A2(new_n207), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n372), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT12), .B1(new_n388), .B2(new_n363), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT12), .ZN(new_n390));
  AOI211_X1 g204(.A(new_n390), .B(new_n362), .C1(new_n387), .C2(new_n372), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n350), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n346), .B(new_n193), .C1(new_n386), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n393), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n380), .A2(new_n396), .B1(new_n349), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G469), .B1(new_n398), .B2(G902), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G221), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT9), .B(G234), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n403), .B2(new_n193), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G140), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G125), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n208), .A2(G140), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT74), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n208), .A2(KEYINPUT74), .A3(G140), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n208), .A2(G140), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(G146), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n200), .B1(new_n412), .B2(new_n414), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n190), .A2(new_n187), .A3(G214), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT90), .A2(G143), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(KEYINPUT90), .A2(G143), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OR2_X1    g237(.A1(KEYINPUT90), .A2(G143), .ZN(new_n424));
  NOR2_X1   g238(.A1(G237), .A2(G953), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G214), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n358), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT17), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n424), .A2(new_n420), .B1(new_n425), .B2(G214), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n419), .A2(new_n422), .ZN(new_n430));
  OAI21_X1  g244(.A(G131), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n423), .A2(new_n358), .A3(new_n426), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n418), .B(new_n428), .C1(KEYINPUT17), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n410), .A2(new_n411), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT92), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(G146), .A3(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n407), .A2(G125), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT75), .B1(new_n413), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT75), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n408), .A2(new_n409), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n200), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT76), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n441), .A2(KEYINPUT76), .A3(new_n200), .A4(new_n443), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n439), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT18), .A2(G131), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n423), .A2(new_n426), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(KEYINPUT91), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n423), .A2(new_n453), .A3(new_n426), .ZN(new_n454));
  INV_X1    g268(.A(new_n451), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n450), .B(KEYINPUT93), .Z(new_n456));
  AOI22_X1  g270(.A1(new_n452), .A2(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n449), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n434), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(new_n225), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n434), .A2(new_n458), .A3(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n193), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n466), .A2(G475), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n437), .A2(KEYINPUT19), .A3(new_n438), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n441), .A2(new_n443), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n200), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n417), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT94), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT94), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n423), .A2(new_n358), .A3(new_n426), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n427), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n458), .A3(KEYINPUT96), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n462), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT96), .B1(new_n478), .B2(new_n458), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT97), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n472), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n473), .A3(new_n474), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n410), .A2(KEYINPUT92), .A3(new_n411), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT92), .B1(new_n410), .B2(new_n411), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n444), .A2(new_n445), .ZN(new_n488));
  AOI22_X1  g302(.A1(G146), .A2(new_n487), .B1(new_n488), .B2(new_n447), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT91), .B1(new_n429), .B2(new_n430), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n490), .A2(new_n454), .A3(KEYINPUT18), .A4(G131), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n455), .A2(new_n456), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n483), .A2(new_n484), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT97), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n462), .A4(new_n479), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n464), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT20), .ZN(new_n500));
  NOR2_X1   g314(.A1(G475), .A2(G902), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n499), .B2(new_n501), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n468), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G217), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n402), .A2(new_n506), .A3(G953), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT99), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT14), .A4(G122), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G107), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n254), .A2(new_n256), .A3(G122), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n253), .A2(G122), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n512), .A2(new_n227), .A3(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n197), .A2(G128), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n205), .A2(G143), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n519), .A3(G134), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n353), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT98), .B1(new_n516), .B2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n517), .A2(new_n520), .A3(new_n522), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT98), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n512), .A2(new_n513), .ZN(new_n527));
  OAI211_X1 g341(.A(G107), .B(new_n510), .C1(new_n527), .C2(KEYINPUT14), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT13), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n519), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n521), .A2(new_n532), .A3(G134), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n518), .B(new_n519), .C1(new_n531), .C2(new_n353), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n527), .A2(G107), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n517), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n509), .B1(new_n530), .B2(new_n538), .ZN(new_n539));
  AOI211_X1 g353(.A(KEYINPUT99), .B(new_n537), .C1(new_n524), .C2(new_n529), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n508), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n516), .A2(KEYINPUT98), .A3(new_n523), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n526), .B1(new_n525), .B2(new_n528), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n538), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT99), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n530), .A2(new_n509), .A3(new_n538), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n507), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(KEYINPUT100), .A3(new_n193), .ZN(new_n549));
  INV_X1    g363(.A(G478), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(G902), .B1(new_n541), .B2(new_n547), .ZN(new_n553));
  INV_X1    g367(.A(new_n551), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT100), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n406), .A2(new_n505), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n506), .B1(G234), .B2(new_n193), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n258), .A2(G128), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n205), .A2(KEYINPUT23), .A3(G119), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n258), .A2(G128), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G110), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT24), .B(G110), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n258), .A2(KEYINPUT73), .A3(G128), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n568), .B(new_n569), .C1(new_n258), .C2(G128), .ZN(new_n570));
  OAI221_X1 g384(.A(new_n565), .B1(new_n566), .B2(new_n570), .C1(new_n416), .C2(new_n417), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n566), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(G110), .B2(new_n564), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n573), .B(new_n473), .C1(new_n446), .C2(new_n448), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n401), .A2(new_n189), .A3(G953), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n575), .B(new_n576), .Z(new_n577));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n571), .B2(new_n574), .ZN(new_n580));
  OR3_X1    g394(.A1(new_n579), .A2(KEYINPUT78), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT78), .B1(new_n579), .B2(new_n580), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n560), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n580), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n193), .A3(new_n578), .ZN(new_n585));
  NOR2_X1   g399(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n586), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n583), .B1(new_n590), .B2(new_n558), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G472), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n193), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT31), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n274), .A2(new_n291), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n214), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n357), .B2(new_n361), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT68), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n598), .B(KEYINPUT68), .C1(new_n357), .C2(new_n361), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT64), .B1(new_n351), .B2(G134), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT64), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n605), .A2(new_n353), .A3(G137), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n351), .A2(G134), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G131), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n359), .A2(new_n358), .A3(new_n360), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n367), .A3(new_n368), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT70), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n383), .A2(KEYINPUT70), .A3(new_n611), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n603), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT30), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n611), .A2(new_n371), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n599), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(KEYINPUT30), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n597), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n603), .A2(new_n614), .A3(new_n615), .A4(new_n597), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n425), .A2(G210), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT27), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT26), .B(G101), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n595), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n628), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n620), .B1(new_n616), .B2(KEYINPUT30), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n630), .B(KEYINPUT31), .C1(new_n631), .C2(new_n597), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n623), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n610), .A2(new_n609), .A3(new_n206), .A4(new_n202), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n359), .A2(new_n360), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(G131), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n214), .B1(new_n637), .B2(new_n610), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n596), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT71), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT71), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n619), .A2(new_n641), .A3(new_n596), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT28), .B1(new_n634), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n612), .A2(new_n597), .A3(new_n599), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT28), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n627), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n594), .B1(new_n633), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n616), .A2(new_n596), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT72), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n623), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n616), .A2(KEYINPUT72), .A3(new_n596), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(KEYINPUT28), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n647), .A2(new_n627), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT29), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n617), .A2(new_n621), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n596), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n627), .B1(new_n662), .B2(new_n623), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n640), .A2(new_n642), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n646), .B1(new_n664), .B2(new_n623), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n658), .B1(new_n665), .B2(new_n657), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n193), .B(new_n660), .C1(new_n663), .C2(new_n666), .ZN(new_n667));
  AOI22_X1  g481(.A1(KEYINPUT32), .A2(new_n651), .B1(new_n667), .B2(G472), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT32), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n629), .A2(new_n632), .B1(new_n648), .B2(new_n649), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n669), .B1(new_n670), .B2(new_n594), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n592), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n345), .A2(new_n557), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(new_n238), .Z(G3));
  NAND2_X1  g488(.A1(new_n498), .A2(new_n464), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n477), .A2(new_n473), .A3(new_n474), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n676), .A2(new_n472), .B1(new_n449), .B2(new_n457), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n461), .B1(new_n677), .B2(KEYINPUT96), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n497), .B1(new_n678), .B2(new_n496), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n501), .B1(new_n675), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n503), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n467), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT33), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n548), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n541), .A2(new_n547), .A3(KEYINPUT33), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n550), .A2(G902), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(G478), .B2(new_n553), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT102), .B1(new_n684), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n505), .A2(new_n693), .A3(new_n690), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n339), .A2(new_n196), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n400), .A2(new_n591), .A3(new_n405), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n698), .B(G472), .C1(new_n670), .C2(G902), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n633), .A2(new_n650), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(G472), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n193), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n695), .A2(new_n696), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT34), .B(G104), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G6));
  NOR2_X1   g521(.A1(new_n680), .A2(new_n681), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n468), .B1(new_n708), .B2(new_n504), .ZN(new_n709));
  INV_X1    g523(.A(new_n556), .ZN(new_n710));
  NOR4_X1   g524(.A1(new_n709), .A2(new_n339), .A3(new_n710), .A4(new_n196), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n704), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT35), .B(G107), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G9));
  INV_X1    g528(.A(new_n703), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n590), .A2(new_n558), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n571), .A2(new_n574), .ZN(new_n717));
  INV_X1    g531(.A(new_n577), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT36), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n717), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n559), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n345), .A2(new_n557), .A3(new_n715), .A4(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT37), .B(G110), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G12));
  NAND2_X1  g539(.A1(new_n651), .A2(KEYINPUT32), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n667), .A2(G472), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n671), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n404), .B1(new_n395), .B2(new_n399), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n728), .A2(new_n342), .A3(new_n729), .A4(new_n722), .ZN(new_n730));
  INV_X1    g544(.A(G900), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n194), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n191), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n468), .B(new_n733), .C1(new_n708), .C2(new_n504), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n710), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT103), .B(G128), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G30));
  XNOR2_X1  g552(.A(new_n733), .B(KEYINPUT39), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n729), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT40), .Z(new_n741));
  AND2_X1   g555(.A1(new_n654), .A2(new_n655), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n193), .B1(new_n742), .B2(new_n627), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n627), .B1(new_n622), .B2(new_n634), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(G472), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n726), .A2(new_n671), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n337), .B(new_n748), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n684), .A2(new_n722), .A3(new_n341), .A4(new_n710), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n741), .A2(new_n747), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G143), .ZN(G45));
  INV_X1    g566(.A(new_n733), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n684), .A2(new_n691), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n730), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G146), .ZN(G48));
  OAI21_X1  g570(.A(new_n193), .B1(new_n386), .B2(new_n394), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(G469), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n395), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n404), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n695), .A2(new_n672), .A3(new_n696), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT41), .B(G113), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G15));
  NAND3_X1  g577(.A1(new_n711), .A2(new_n672), .A3(new_n760), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  INV_X1    g579(.A(new_n722), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n668), .B2(new_n671), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n342), .A2(new_n758), .A3(new_n405), .A4(new_n395), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n505), .A2(new_n196), .A3(new_n556), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G119), .ZN(G21));
  NOR3_X1   g586(.A1(new_n684), .A2(new_n339), .A3(new_n710), .ZN(new_n773));
  INV_X1    g587(.A(new_n633), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n627), .B1(new_n656), .B2(new_n647), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n593), .B(new_n193), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(G472), .B1(new_n670), .B2(G902), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n776), .A2(new_n777), .A3(new_n591), .ZN(new_n778));
  INV_X1    g592(.A(new_n196), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n773), .A2(new_n778), .A3(new_n779), .A4(new_n760), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  NAND3_X1  g595(.A1(new_n505), .A2(new_n690), .A3(new_n733), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n722), .A2(new_n776), .A3(new_n777), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n782), .A2(new_n783), .A3(new_n768), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n208), .ZN(G27));
  NAND3_X1  g599(.A1(new_n325), .A2(new_n336), .A3(new_n338), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n325), .A2(new_n336), .A3(KEYINPUT106), .A4(new_n338), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n788), .B(new_n789), .C1(new_n729), .C2(KEYINPUT105), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n729), .A2(KEYINPUT105), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n672), .A3(new_n754), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT42), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT107), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n651), .B2(KEYINPUT32), .ZN(new_n798));
  OAI211_X1 g612(.A(KEYINPUT107), .B(new_n669), .C1(new_n670), .C2(new_n594), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n726), .A3(new_n727), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(KEYINPUT42), .A3(new_n591), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT105), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n802), .B(new_n404), .C1(new_n395), .C2(new_n399), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n790), .A2(new_n782), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n796), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n788), .A2(new_n789), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n406), .A2(new_n802), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n754), .A2(new_n806), .A3(new_n807), .A4(new_n792), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n800), .A2(KEYINPUT42), .A3(new_n591), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT108), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n795), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g625(.A(KEYINPUT109), .B(G131), .Z(new_n812));
  XNOR2_X1  g626(.A(new_n811), .B(new_n812), .ZN(G33));
  NAND4_X1  g627(.A1(new_n791), .A2(new_n672), .A3(new_n735), .A4(new_n792), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G134), .ZN(G36));
  OR2_X1    g629(.A1(new_n398), .A2(KEYINPUT45), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n398), .A2(KEYINPUT45), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(G469), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(G469), .A2(G902), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT46), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(new_n822), .B(KEYINPUT110), .Z(new_n823));
  INV_X1    g637(.A(new_n395), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n820), .B2(new_n821), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n404), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n788), .A2(new_n789), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n684), .A2(new_n690), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(KEYINPUT43), .Z(new_n829));
  NOR2_X1   g643(.A1(new_n715), .A2(new_n766), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT44), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(KEYINPUT44), .A3(new_n830), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n826), .A2(new_n833), .A3(new_n739), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  NOR4_X1   g650(.A1(new_n728), .A2(new_n782), .A3(new_n827), .A4(new_n591), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n826), .A2(KEYINPUT47), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n826), .A2(KEYINPUT47), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  OR2_X1    g656(.A1(new_n747), .A2(new_n828), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n759), .B(KEYINPUT49), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n591), .A2(new_n338), .A3(new_n405), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n843), .A2(new_n844), .A3(new_n749), .A4(new_n845), .ZN(new_n846));
  XOR2_X1   g660(.A(new_n846), .B(KEYINPUT111), .Z(new_n847));
  AND2_X1   g661(.A1(new_n829), .A2(new_n192), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n778), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n839), .A2(new_n840), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n759), .A2(new_n405), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n806), .B(new_n849), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n760), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n827), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n783), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n747), .A2(new_n592), .A3(new_n191), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n854), .A2(new_n684), .A3(new_n691), .A4(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n852), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n853), .A2(new_n338), .A3(new_n749), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n849), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT50), .Z(new_n863));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n849), .A2(new_n769), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n854), .A2(new_n695), .A3(new_n858), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n188), .A3(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n800), .A2(new_n591), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(KEYINPUT115), .B2(KEYINPUT48), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n855), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(new_n868), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n852), .A2(KEYINPUT51), .A3(new_n863), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n857), .A2(new_n859), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT114), .Z(new_n876));
  OAI211_X1 g690(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n556), .B(new_n468), .C1(new_n502), .C2(new_n504), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT112), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n505), .A2(new_n690), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n682), .A2(new_n683), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(KEYINPUT112), .A3(new_n468), .A4(new_n556), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n345), .A3(new_n704), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n761), .A2(new_n886), .A3(new_n673), .A4(new_n780), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n723), .A2(new_n771), .A3(new_n764), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n791), .A2(new_n754), .A3(new_n856), .A4(new_n792), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n827), .A2(new_n734), .A3(new_n556), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n767), .A3(new_n729), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n814), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n811), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n784), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n406), .A2(new_n722), .A3(new_n753), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n747), .A3(new_n773), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n736), .A2(new_n755), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT52), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n784), .B1(new_n730), .B2(new_n735), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(new_n755), .A4(new_n898), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n878), .B1(new_n895), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n801), .A2(new_n804), .A3(new_n796), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT108), .B1(new_n808), .B2(new_n809), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n893), .B1(new_n908), .B2(new_n795), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n889), .A3(new_n900), .A4(new_n903), .ZN(new_n910));
  OR2_X1    g724(.A1(new_n901), .A2(new_n902), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n878), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n905), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT54), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(KEYINPUT53), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT113), .B(new_n878), .C1(new_n895), .C2(new_n904), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT113), .B1(new_n910), .B2(new_n878), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n915), .B1(new_n921), .B2(KEYINPUT54), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n864), .A2(new_n877), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(G952), .A2(G953), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n847), .B1(new_n923), .B2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n910), .A2(new_n916), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT113), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n905), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n926), .B1(new_n928), .B2(new_n918), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n193), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(G210), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n329), .A2(new_n330), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT116), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT117), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n223), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n931), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n937), .B1(new_n931), .B2(new_n932), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n187), .A2(G952), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(G51));
  XNOR2_X1  g755(.A(new_n921), .B(KEYINPUT54), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n819), .B(KEYINPUT57), .Z(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n386), .B2(new_n394), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n818), .B(KEYINPUT118), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n930), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n940), .B1(new_n945), .B2(new_n947), .ZN(G54));
  NAND3_X1  g762(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n949));
  INV_X1    g763(.A(new_n499), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n949), .A2(new_n950), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n951), .A2(new_n952), .A3(new_n940), .ZN(G60));
  AND2_X1   g767(.A1(new_n686), .A2(new_n687), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT119), .ZN(new_n955));
  XNOR2_X1  g769(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n550), .A2(new_n193), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n955), .B1(new_n922), .B2(new_n958), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n955), .A2(new_n958), .ZN(new_n960));
  AOI211_X1 g774(.A(new_n940), .B(new_n959), .C1(new_n942), .C2(new_n960), .ZN(G63));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT60), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n929), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n964), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n581), .A2(new_n582), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n940), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n720), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n965), .B2(new_n967), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT122), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n971), .B(new_n974), .C1(new_n975), .C2(KEYINPUT61), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n969), .A2(new_n975), .A3(new_n970), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n969), .A2(new_n970), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n977), .B(new_n978), .C1(new_n979), .C2(new_n973), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n976), .A2(new_n980), .ZN(G66));
  OAI21_X1  g795(.A(G953), .B1(new_n195), .B2(new_n217), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n889), .B2(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n934), .B1(G898), .B2(new_n187), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G69));
  NAND2_X1  g799(.A1(new_n469), .A2(new_n471), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT123), .Z(new_n987));
  XNOR2_X1  g801(.A(new_n661), .B(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(G900), .B2(G953), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  INV_X1    g805(.A(new_n869), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n773), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n826), .A2(new_n739), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT126), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n826), .A2(new_n997), .A3(new_n739), .A4(new_n994), .ZN(new_n998));
  AOI22_X1  g812(.A1(new_n996), .A2(new_n998), .B1(new_n795), .B2(new_n908), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n835), .A2(new_n814), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n901), .A2(new_n755), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n841), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n991), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n841), .A2(new_n1002), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1005), .A2(new_n999), .A3(new_n1001), .A4(KEYINPUT127), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n990), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1002), .A2(new_n751), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1010));
  NOR2_X1   g824(.A1(new_n827), .A2(new_n740), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n885), .A2(new_n1011), .A3(new_n672), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n835), .A2(KEYINPUT124), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(KEYINPUT124), .B1(new_n835), .B2(new_n1012), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n1010), .B(new_n841), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n187), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n989), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT125), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1017), .A2(KEYINPUT125), .A3(new_n989), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1008), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n187), .B1(G227), .B2(G900), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1023), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1008), .A2(new_n1020), .A3(new_n1025), .A4(new_n1021), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1024), .A2(new_n1026), .ZN(G72));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  INV_X1    g843(.A(new_n889), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1016), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n745), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n622), .A2(new_n628), .ZN(new_n1033));
  OAI211_X1 g847(.A(new_n914), .B(new_n1029), .C1(new_n1033), .C2(new_n663), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1032), .A2(new_n970), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1029), .B1(new_n1007), .B2(new_n1030), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n662), .A2(new_n623), .A3(new_n649), .ZN(new_n1037));
  INV_X1    g851(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1035), .B1(new_n1036), .B2(new_n1038), .ZN(G57));
endmodule


