//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT92), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n205), .A2(new_n208), .A3(G43gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n204), .B1(new_n210), .B2(KEYINPUT93), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT14), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n214), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(new_n215), .B2(new_n212), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n206), .A2(new_n218), .A3(new_n207), .A4(new_n209), .ZN(new_n219));
  INV_X1    g018(.A(new_n216), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n204), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT17), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n223), .B(new_n224), .C1(new_n216), .C2(new_n211), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(G1gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G1gat), .B2(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n222), .A2(new_n225), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n217), .A2(new_n221), .ZN(new_n233));
  INV_X1    g032(.A(new_n231), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n236), .A2(KEYINPUT94), .B1(G229gat), .B2(G233gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n232), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n236), .A2(KEYINPUT94), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT13), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n235), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n233), .A2(new_n234), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n232), .A2(new_n235), .A3(new_n239), .A4(new_n237), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n241), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT91), .ZN(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G197gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT11), .ZN(new_n253));
  INV_X1    g052(.A(G169gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT12), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n249), .A2(new_n250), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n249), .B2(new_n250), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT24), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(G183gat), .A3(G190gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(G183gat), .A2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT24), .ZN(new_n265));
  NOR2_X1   g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT66), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(G169gat), .A3(G176gat), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n269), .A2(new_n272), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n278), .B(new_n263), .C1(new_n265), .C2(new_n266), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n268), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n277), .A2(KEYINPUT25), .ZN(new_n283));
  INV_X1    g082(.A(new_n267), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT27), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT28), .B1(new_n288), .B2(KEYINPUT67), .ZN(new_n289));
  INV_X1    g088(.A(G190gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n289), .B(new_n290), .C1(KEYINPUT67), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n290), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n292), .A2(new_n294), .A3(new_n264), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n276), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n297), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT69), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n270), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n296), .A2(new_n305), .A3(new_n298), .A4(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n295), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n261), .B1(new_n286), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT75), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n260), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n295), .A2(new_n307), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n281), .A2(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n311), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n282), .A2(new_n285), .B1(new_n295), .B2(new_n307), .ZN(new_n317));
  OAI211_X1 g116(.A(KEYINPUT77), .B(new_n316), .C1(new_n317), .C2(new_n261), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n312), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n320), .B(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G197gat), .B(G204gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G211gat), .B(G218gat), .Z(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n325), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n327), .A3(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n316), .B1(new_n317), .B2(KEYINPUT29), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n329), .A3(new_n315), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT78), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n332), .A2(new_n335), .A3(new_n329), .A4(new_n315), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G8gat), .B(G36gat), .Z(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(G64gat), .ZN(new_n339));
  INV_X1    g138(.A(G92gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n316), .B1(new_n286), .B2(new_n308), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n313), .B2(new_n314), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n345), .B2(new_n316), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n335), .B1(new_n346), .B2(new_n329), .ZN(new_n347));
  AND4_X1   g146(.A1(new_n335), .A2(new_n332), .A3(new_n329), .A4(new_n315), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n341), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(new_n331), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n351), .A3(KEYINPUT30), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n337), .A2(KEYINPUT30), .A3(new_n341), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  INV_X1    g154(.A(G134gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G127gat), .ZN(new_n357));
  INV_X1    g156(.A(G127gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G134gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT71), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT1), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G113gat), .ZN(new_n366));
  OR3_X1    g165(.A1(new_n366), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT70), .B1(new_n366), .B2(G120gat), .ZN(new_n368));
  INV_X1    g167(.A(G120gat), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n367), .B(new_n368), .C1(G113gat), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n366), .A2(G120gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n369), .A2(G113gat), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n365), .A2(new_n370), .B1(new_n374), .B2(new_n360), .ZN(new_n375));
  INV_X1    g174(.A(G155gat), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G141gat), .B(G148gat), .Z(new_n381));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  INV_X1    g183(.A(new_n379), .ZN(new_n385));
  NOR2_X1   g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G141gat), .B(G148gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n379), .B1(new_n378), .B2(KEYINPUT2), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n381), .A3(KEYINPUT79), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n383), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n355), .B1(new_n375), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n360), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n362), .A2(new_n364), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n371), .A3(new_n370), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n392), .A2(new_n355), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT81), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n375), .A2(new_n392), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n379), .B(new_n378), .C1(new_n388), .C2(KEYINPUT2), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n387), .A2(new_n384), .A3(new_n388), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT79), .B1(new_n390), .B2(new_n381), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n403), .B1(new_n407), .B2(KEYINPUT3), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n392), .A2(KEYINPUT80), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n375), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(KEYINPUT3), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n400), .A2(new_n402), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  NAND2_X1  g213(.A1(G225gat), .A2(G233gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n408), .A2(new_n410), .ZN(new_n417));
  INV_X1    g216(.A(new_n375), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n418), .A3(new_n412), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n394), .A2(new_n398), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n418), .A2(new_n407), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n401), .ZN(new_n423));
  INV_X1    g222(.A(new_n415), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n414), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT0), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(G57gat), .ZN(new_n430));
  INV_X1    g229(.A(G85gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n432), .A3(new_n426), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n354), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G78gat), .B(G106gat), .Z(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(KEYINPUT31), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(new_n208), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT83), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n261), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n329), .B1(new_n417), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n322), .A2(KEYINPUT82), .A3(new_n327), .A4(new_n323), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n447), .B(new_n449), .C1(new_n329), .C2(KEYINPUT82), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n392), .B1(new_n450), .B2(new_n409), .ZN(new_n451));
  INV_X1    g250(.A(G228gat), .ZN(new_n452));
  INV_X1    g251(.A(G233gat), .ZN(new_n453));
  OAI22_X1  g252(.A1(new_n448), .A2(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT29), .B1(new_n326), .B2(new_n328), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n407), .B1(new_n456), .B2(KEYINPUT3), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n261), .B1(new_n408), .B2(new_n410), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n455), .B(new_n457), .C1(new_n458), .C2(new_n329), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n444), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(G22gat), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G22gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n454), .A2(new_n463), .A3(new_n459), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n446), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n454), .A2(new_n463), .A3(new_n459), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n463), .B1(new_n454), .B2(new_n459), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n466), .A2(new_n467), .A3(new_n445), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n441), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n375), .B1(new_n313), .B2(new_n314), .ZN(new_n472));
  INV_X1    g271(.A(G227gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n453), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n286), .A2(new_n418), .A3(new_n308), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT32), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G43gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(G71gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(G99gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT33), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n476), .A2(KEYINPUT72), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT72), .B1(new_n476), .B2(new_n482), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n477), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n476), .B(KEYINPUT32), .C1(new_n482), .C2(new_n480), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n475), .ZN(new_n488));
  INV_X1    g287(.A(new_n474), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI211_X1 g289(.A(KEYINPUT34), .B(new_n474), .C1(new_n472), .C2(new_n475), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n485), .B2(new_n486), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(KEYINPUT36), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n485), .A2(new_n486), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT73), .ZN(new_n498));
  INV_X1    g297(.A(new_n492), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n492), .A3(new_n486), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT73), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n496), .B1(new_n504), .B2(KEYINPUT36), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n349), .B2(new_n331), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n506), .B1(new_n508), .B2(new_n350), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n331), .A2(new_n507), .A3(new_n334), .A4(new_n336), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n319), .A2(new_n330), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n334), .A2(new_n336), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT37), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(KEYINPUT88), .A3(new_n341), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n509), .A2(KEYINPUT38), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n319), .A2(new_n329), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n346), .A2(new_n330), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT37), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n516), .A2(new_n517), .A3(new_n520), .A4(KEYINPUT37), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n519), .A2(new_n341), .A3(new_n521), .A4(new_n510), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT38), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n439), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n469), .B1(new_n525), .B2(new_n351), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT86), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n393), .B1(KEYINPUT81), .B2(new_n398), .ZN(new_n528));
  INV_X1    g327(.A(new_n402), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n419), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n424), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n422), .A2(new_n415), .A3(new_n401), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n531), .A2(KEYINPUT39), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n534), .A3(new_n424), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n432), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT85), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT85), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n535), .A2(new_n538), .A3(new_n432), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n533), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n527), .B1(new_n540), .B2(KEYINPUT40), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n531), .A2(KEYINPUT39), .A3(new_n532), .ZN(new_n542));
  INV_X1    g341(.A(new_n539), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n538), .B1(new_n535), .B2(new_n432), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT40), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(KEYINPUT86), .A3(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n541), .A2(new_n434), .A3(new_n547), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT84), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT84), .B1(new_n352), .B2(new_n353), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n540), .A2(KEYINPUT40), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI211_X1 g352(.A(new_n471), .B(new_n505), .C1(new_n526), .C2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n437), .A2(new_n438), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT89), .B(KEYINPUT35), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n500), .A2(new_n501), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n469), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n557), .B(new_n559), .C1(new_n549), .C2(new_n550), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT90), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n497), .A2(KEYINPUT73), .A3(new_n499), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n495), .B2(new_n498), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n564), .B2(new_n469), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n504), .A2(KEYINPUT90), .A3(new_n470), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n441), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n561), .B1(new_n567), .B2(KEYINPUT35), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n259), .B1(new_n554), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g370(.A(KEYINPUT95), .B(new_n259), .C1(new_n554), .C2(new_n568), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G85gat), .A2(G92gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT7), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(KEYINPUT8), .A2(new_n576), .B1(new_n431), .B2(new_n340), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G99gat), .B(G106gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(KEYINPUT97), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT9), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G57gat), .B(G64gat), .Z(new_n595));
  NAND3_X1  g394(.A1(new_n586), .A2(new_n591), .A3(new_n592), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n596), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n599), .A2(new_n588), .A3(new_n593), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(new_n589), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n582), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n590), .A2(new_n597), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n589), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT98), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n581), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n604), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n580), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n602), .A2(new_n605), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n611), .A2(KEYINPUT10), .A3(new_n580), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G230gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n453), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n606), .A2(new_n609), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n615), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  INV_X1    g420(.A(G176gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G204gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n617), .A2(new_n619), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(new_n358), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n234), .B1(new_n611), .B2(KEYINPUT21), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n631), .B(G127gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g438(.A(G155gat), .B(G183gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n635), .A2(new_n637), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(G211gat), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n642), .A2(new_n647), .A3(new_n644), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(G232gat), .A2(G233gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G162gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(G190gat), .B(G218gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n222), .A2(new_n225), .A3(new_n581), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n657), .A2(KEYINPUT99), .B1(KEYINPUT41), .B2(new_n652), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n233), .A2(new_n580), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT99), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n222), .A2(new_n225), .A3(new_n660), .A4(new_n581), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G134gat), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n658), .A2(new_n356), .A3(new_n659), .A4(new_n661), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n656), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(new_n664), .A3(new_n656), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n651), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n573), .A2(new_n630), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n555), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g472(.A(new_n230), .B1(new_n671), .B2(new_n551), .ZN(new_n674));
  INV_X1    g473(.A(new_n551), .ZN(new_n675));
  NOR2_X1   g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n227), .A2(new_n230), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n670), .A2(new_n675), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT42), .B1(new_n674), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(KEYINPUT42), .B2(new_n678), .ZN(G1325gat));
  AND3_X1   g479(.A1(new_n671), .A2(G15gat), .A3(new_n505), .ZN(new_n681));
  AOI21_X1  g480(.A(G15gat), .B1(new_n671), .B2(new_n495), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(G1326gat));
  NOR2_X1   g482(.A1(new_n670), .A2(new_n470), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT43), .B(G22gat), .Z(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(G1327gat));
  INV_X1    g485(.A(new_n668), .ZN(new_n687));
  INV_X1    g486(.A(new_n651), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n629), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI211_X1 g489(.A(new_n687), .B(new_n690), .C1(new_n571), .C2(new_n572), .ZN(new_n691));
  INV_X1    g490(.A(G29gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n555), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n695), .B(new_n668), .C1(new_n554), .C2(new_n568), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT100), .B(new_n668), .C1(new_n554), .C2(new_n568), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT44), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n259), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n690), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n439), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n694), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n694), .A2(KEYINPUT102), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1328gat));
  NAND2_X1  g511(.A1(new_n691), .A2(new_n551), .ZN(new_n713));
  OAI22_X1  g512(.A1(new_n713), .A2(G36gat), .B1(KEYINPUT103), .B2(KEYINPUT46), .ZN(new_n714));
  NAND2_X1  g513(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n714), .B(new_n715), .Z(new_n716));
  OAI21_X1  g515(.A(G36gat), .B1(new_n706), .B2(new_n675), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1329gat));
  AOI21_X1  g517(.A(KEYINPUT90), .B1(new_n504), .B2(new_n470), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n562), .B(new_n469), .C1(new_n502), .C2(new_n503), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n719), .A2(new_n720), .A3(new_n440), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT35), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n560), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n471), .ZN(new_n724));
  INV_X1    g523(.A(new_n505), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n514), .A2(new_n510), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n350), .B1(new_n337), .B2(KEYINPUT37), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT38), .B1(new_n728), .B2(KEYINPUT88), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n524), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n730), .A2(new_n555), .A3(new_n351), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n470), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n724), .B(new_n725), .C1(new_n726), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n723), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT95), .B1(new_n734), .B2(new_n259), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n570), .B(new_n704), .C1(new_n723), .C2(new_n733), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n668), .B(new_n689), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(G43gat), .A3(new_n558), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n703), .A2(new_n505), .A3(new_n705), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT47), .ZN(G1330gat));
  AOI22_X1  g540(.A1(new_n697), .A2(new_n696), .B1(new_n699), .B2(KEYINPUT44), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT44), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n469), .B(new_n705), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G50gat), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT48), .B1(new_n745), .B2(KEYINPUT105), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n573), .A2(new_n749), .A3(new_n668), .A4(new_n689), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n748), .A2(new_n208), .A3(new_n469), .A4(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n751), .A2(new_n752), .A3(new_n745), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(new_n745), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n747), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n469), .B1(new_n691), .B2(new_n749), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n750), .A2(new_n208), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n745), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT106), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n751), .A2(new_n752), .A3(new_n745), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n759), .A2(new_n746), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n755), .A2(new_n761), .ZN(G1331gat));
  NAND4_X1  g561(.A1(new_n734), .A2(new_n629), .A3(new_n704), .A4(new_n669), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n439), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(G57gat), .Z(G1332gat));
  AOI211_X1 g564(.A(new_n675), .B(new_n763), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT107), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n763), .B2(new_n725), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n495), .A2(new_n583), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n763), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g572(.A1(new_n763), .A2(new_n470), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(new_n584), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n688), .A2(new_n259), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n734), .A2(new_n668), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT108), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n782), .A2(new_n431), .A3(new_n555), .A4(new_n629), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n703), .A2(new_n629), .A3(new_n776), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n439), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1336gat));
  NAND4_X1  g585(.A1(new_n703), .A2(new_n629), .A3(new_n551), .A4(new_n776), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT109), .B1(new_n787), .B2(G92gat), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(KEYINPUT52), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n630), .B1(new_n779), .B2(new_n780), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n675), .A2(G92gat), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n787), .A2(G92gat), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n789), .B(new_n792), .ZN(G1337gat));
  NOR3_X1   g592(.A1(new_n558), .A2(G99gat), .A3(new_n630), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT110), .Z(new_n795));
  NAND2_X1  g594(.A1(new_n782), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(G99gat), .B1(new_n784), .B2(new_n725), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1338gat));
  OAI21_X1  g597(.A(G106gat), .B1(new_n784), .B2(new_n470), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n470), .A2(G106gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n802), .B(new_n803), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n256), .A2(new_n241), .A3(new_n247), .A4(new_n248), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n245), .A2(new_n246), .A3(new_n244), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n242), .B1(new_n232), .B2(new_n235), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n255), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n667), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(new_n665), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n610), .A2(new_n615), .A3(new_n612), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n617), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n615), .B1(new_n610), .B2(new_n612), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n627), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n628), .ZN(new_n819));
  AOI21_X1  g618(.A(KEYINPUT55), .B1(new_n814), .B2(new_n817), .ZN(new_n820));
  OR2_X1    g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n805), .B1(new_n812), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n819), .A2(new_n820), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n668), .A2(new_n823), .A3(KEYINPUT112), .A4(new_n810), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n629), .ZN(new_n826));
  INV_X1    g625(.A(new_n258), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n249), .A2(new_n250), .A3(new_n256), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n628), .A3(new_n828), .A4(new_n818), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n826), .B1(new_n829), .B2(new_n820), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n687), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n688), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  NOR4_X1   g631(.A1(new_n651), .A2(new_n668), .A3(new_n629), .A4(new_n259), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT113), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n669), .A2(new_n630), .A3(new_n704), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n822), .A2(new_n824), .B1(new_n830), .B2(new_n687), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n835), .B(new_n836), .C1(new_n837), .C2(new_n688), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(new_n555), .A3(new_n675), .A4(new_n559), .ZN(new_n840));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840), .B2(new_n704), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n839), .A2(new_n555), .A3(new_n565), .A4(new_n566), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n675), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n259), .A2(new_n366), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(G1340gat));
  OAI21_X1  g645(.A(G120gat), .B1(new_n840), .B2(new_n630), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n629), .A2(new_n369), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n844), .B2(new_n848), .ZN(G1341gat));
  NOR3_X1   g648(.A1(new_n840), .A2(new_n358), .A3(new_n651), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n675), .A3(new_n688), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n358), .ZN(G1342gat));
  NOR3_X1   g651(.A1(new_n844), .A2(G134gat), .A3(new_n687), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n840), .B2(new_n687), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  AND2_X1   g657(.A1(new_n839), .A2(new_n469), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n725), .A2(new_n555), .A3(new_n675), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(G141gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n864), .A3(new_n259), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n859), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n822), .A2(new_n824), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n814), .A2(new_n817), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT115), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT55), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n814), .A2(new_n872), .A3(new_n817), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n819), .A2(new_n257), .A3(new_n258), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n871), .A4(new_n873), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n668), .B1(new_n879), .B2(new_n826), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n651), .B1(new_n868), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT117), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n835), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n866), .B1(new_n883), .B2(new_n469), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n860), .A3(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n259), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n865), .B1(new_n886), .B2(new_n864), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n865), .B2(KEYINPUT118), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n887), .B(new_n889), .ZN(G1344gat));
  INV_X1    g689(.A(G148gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n863), .A2(new_n891), .A3(new_n629), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n891), .C1(new_n885), .C2(new_n629), .ZN(new_n893));
  XNOR2_X1  g692(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n834), .A2(new_n838), .A3(KEYINPUT57), .A4(new_n469), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n812), .A2(new_n821), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n651), .B1(new_n880), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n835), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(KEYINPUT121), .A3(new_n835), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n469), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n866), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n903), .B2(new_n866), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n629), .A3(new_n861), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n894), .B1(new_n908), .B2(G148gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n909), .ZN(G1345gat));
  INV_X1    g709(.A(new_n885), .ZN(new_n911));
  OAI21_X1  g710(.A(G155gat), .B1(new_n911), .B2(new_n651), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n863), .A2(new_n376), .A3(new_n688), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1346gat));
  OAI21_X1  g713(.A(G162gat), .B1(new_n911), .B2(new_n687), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n863), .A2(new_n377), .A3(new_n668), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n675), .A2(new_n555), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n839), .A2(new_n559), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919), .B2(new_n704), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(KEYINPUT123), .Z(new_n921));
  AND4_X1   g720(.A1(new_n565), .A2(new_n839), .A3(new_n566), .A4(new_n918), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n254), .A3(new_n259), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1348gat));
  NOR3_X1   g723(.A1(new_n919), .A2(new_n622), .A3(new_n630), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n922), .A2(new_n629), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(new_n622), .ZN(G1349gat));
  OR3_X1    g726(.A1(new_n919), .A2(KEYINPUT124), .A3(new_n651), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT124), .B1(new_n919), .B2(new_n651), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(G183gat), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n922), .A2(new_n291), .A3(new_n688), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n919), .B2(new_n687), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n922), .A2(new_n290), .A3(new_n668), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(new_n937), .ZN(G1351gat));
  INV_X1    g737(.A(new_n907), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n918), .A2(new_n725), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n939), .A2(new_n704), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(G197gat), .ZN(new_n942));
  INV_X1    g741(.A(new_n940), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n859), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n259), .A2(new_n942), .ZN(new_n945));
  OAI22_X1  g744(.A1(new_n941), .A2(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  NOR3_X1   g745(.A1(new_n944), .A2(G204gat), .A3(new_n630), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n939), .A2(new_n630), .A3(new_n940), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n624), .ZN(G1353gat));
  OR3_X1    g749(.A1(new_n944), .A2(G211gat), .A3(new_n651), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n907), .A2(new_n688), .A3(new_n943), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n907), .A2(KEYINPUT126), .A3(new_n688), .A4(new_n943), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(G211gat), .A3(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(G1354gat));
  INV_X1    g759(.A(G218gat), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n961), .B1(new_n944), .B2(new_n687), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT127), .Z(new_n963));
  NOR2_X1   g762(.A1(new_n939), .A2(new_n940), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n687), .A2(new_n961), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(G1355gat));
endmodule


