//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  AOI21_X1  g008(.A(G128), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(KEYINPUT1), .A3(G146), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n192), .A3(new_n194), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT0), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(new_n200), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n209), .A2(new_n210), .B1(KEYINPUT0), .B2(G128), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n206), .B(G125), .C1(new_n211), .C2(new_n204), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT84), .B1(new_n203), .B2(new_n212), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n212), .A2(KEYINPUT84), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G224), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(G224), .B(new_n216), .C1(new_n213), .C2(new_n214), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(G110), .B(G122), .ZN(new_n222));
  XOR2_X1   g036(.A(new_n222), .B(KEYINPUT81), .Z(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G113), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G119), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n225), .B(new_n227), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n225), .A2(new_n227), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n239));
  INV_X1    g053(.A(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G104), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(G107), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G101), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(G101), .B1(new_n237), .B2(G107), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n238), .A2(new_n247), .A3(new_n241), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT78), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n238), .A2(new_n247), .A3(new_n241), .A4(KEYINPUT78), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n244), .B1(new_n243), .B2(G101), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n246), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n240), .A2(G104), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n242), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n256), .A2(G101), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(new_n250), .B2(new_n251), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n224), .B1(new_n229), .B2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n259), .A2(new_n261), .B1(new_n234), .B2(new_n233), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n223), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT6), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n252), .A2(new_n253), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n236), .A2(new_n245), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n266), .A2(new_n267), .B1(new_n258), .B2(new_n262), .ZN(new_n268));
  INV_X1    g082(.A(new_n223), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT82), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(new_n268), .B2(new_n222), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT82), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n223), .C1(new_n254), .C2(new_n263), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT83), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n270), .A2(new_n272), .A3(new_n274), .A4(new_n277), .ZN(new_n278));
  AOI211_X1 g092(.A(new_n221), .B(new_n265), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n217), .A2(KEYINPUT7), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n213), .A2(new_n214), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(KEYINPUT87), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n268), .A2(new_n222), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n203), .A2(new_n212), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n280), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n222), .B(KEYINPUT8), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n257), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n252), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT86), .B1(new_n291), .B2(KEYINPUT85), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n262), .B1(new_n258), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(KEYINPUT86), .B(new_n262), .C1(new_n291), .C2(KEYINPUT85), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n295), .A2(new_n296), .B1(new_n281), .B2(KEYINPUT87), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n287), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n190), .B1(new_n279), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n276), .A2(new_n278), .ZN(new_n301));
  INV_X1    g115(.A(new_n265), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n220), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n298), .A3(new_n189), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n188), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  OAI21_X1  g120(.A(G221), .B1(new_n306), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n198), .B2(new_n202), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n258), .A2(new_n309), .A3(KEYINPUT80), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT80), .B1(new_n258), .B2(new_n309), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G134), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G134), .ZN(new_n316));
  INV_X1    g130(.A(G137), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT11), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(KEYINPUT66), .A2(G131), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(KEYINPUT11), .A3(G134), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n319), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n325), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n320), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT79), .B1(new_n195), .B2(new_n197), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(new_n196), .C1(new_n204), .C2(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n202), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n258), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n206), .B1(new_n211), .B2(new_n204), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n336), .A2(new_n245), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n335), .A2(new_n308), .B1(new_n337), .B2(new_n266), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n312), .A2(new_n330), .A3(new_n338), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n202), .B(new_n196), .C1(G128), .C2(new_n204), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n291), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n335), .ZN(new_n343));
  INV_X1    g157(.A(new_n330), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT12), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT12), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n346), .B(new_n330), .C1(new_n342), .C2(new_n335), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n339), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G110), .B(G140), .ZN(new_n349));
  INV_X1    g163(.A(G227), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G953), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n335), .A2(new_n308), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n258), .A2(new_n309), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT80), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n337), .A2(new_n266), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n258), .A2(new_n309), .A3(KEYINPUT80), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n354), .A2(new_n357), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n344), .ZN(new_n361));
  INV_X1    g175(.A(new_n352), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n339), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(G469), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(G469), .A2(G902), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n360), .A2(new_n344), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n330), .B1(new_n312), .B2(new_n338), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n352), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n339), .B(new_n362), .C1(new_n345), .C2(new_n347), .ZN(new_n370));
  AOI211_X1 g184(.A(G469), .B(G902), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n307), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G902), .ZN(new_n374));
  XNOR2_X1  g188(.A(G125), .B(G140), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT75), .B1(new_n375), .B2(new_n191), .ZN(new_n376));
  INV_X1    g190(.A(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G125), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n199), .A2(G140), .ZN(new_n379));
  AND4_X1   g193(.A1(KEYINPUT75), .A2(new_n378), .A3(new_n379), .A4(new_n191), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(KEYINPUT72), .ZN(new_n381));
  OR3_X1    g195(.A1(new_n377), .A2(KEYINPUT72), .A3(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  OAI22_X1  g197(.A1(new_n376), .A2(new_n380), .B1(new_n383), .B2(new_n191), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n193), .A2(KEYINPUT88), .ZN(new_n385));
  NOR2_X1   g199(.A1(G237), .A2(G953), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n385), .A2(G214), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT88), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G143), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n389), .A2(new_n385), .B1(new_n386), .B2(G214), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT18), .B(G131), .C1(new_n387), .C2(new_n390), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n386), .A2(G214), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n385), .ZN(new_n393));
  NAND2_X1  g207(.A1(KEYINPUT18), .A2(G131), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n389), .A2(new_n385), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n393), .B(new_n394), .C1(new_n395), .C2(new_n392), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n384), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n384), .A2(KEYINPUT89), .A3(new_n391), .A4(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n378), .A2(KEYINPUT16), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT16), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n381), .B2(new_n382), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n405), .B2(KEYINPUT73), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n377), .A2(KEYINPUT72), .A3(G125), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n375), .B2(KEYINPUT72), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT73), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n408), .A2(new_n409), .A3(new_n404), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n191), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n409), .B1(new_n408), .B2(new_n404), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n383), .A2(KEYINPUT73), .A3(KEYINPUT16), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n412), .A2(G146), .A3(new_n413), .A4(new_n403), .ZN(new_n414));
  OAI21_X1  g228(.A(G131), .B1(new_n387), .B2(new_n390), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT17), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G131), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n393), .B(new_n418), .C1(new_n395), .C2(new_n392), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n415), .A3(new_n416), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n411), .A2(new_n414), .A3(new_n417), .A4(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n237), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n401), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n401), .B2(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n374), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G475), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT74), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n414), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n383), .A2(KEYINPUT16), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n402), .B1(new_n431), .B2(new_n409), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n432), .A2(KEYINPUT74), .A3(G146), .A4(new_n413), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n383), .A2(KEYINPUT19), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(KEYINPUT19), .B2(new_n375), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n435), .A2(new_n191), .B1(new_n419), .B2(new_n415), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n430), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n401), .ZN(new_n438));
  INV_X1    g252(.A(new_n423), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n401), .A2(new_n421), .A3(new_n423), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n428), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n423), .B1(new_n437), .B2(new_n401), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n428), .B(new_n443), .C1(new_n424), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n427), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT90), .B1(new_n193), .B2(G128), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT90), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n200), .A3(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n193), .A2(G128), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n314), .A2(new_n316), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n449), .A2(new_n451), .B1(G128), .B2(new_n193), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT65), .B(G134), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G122), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G116), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT14), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n228), .A2(G122), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n461), .A2(G116), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n463), .B(G107), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n228), .A2(G122), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n462), .B(new_n467), .C1(KEYINPUT14), .C2(new_n240), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G107), .B1(new_n464), .B2(new_n465), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n462), .A2(new_n467), .A3(new_n240), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n457), .A2(new_n458), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n453), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n193), .A2(KEYINPUT13), .A3(G128), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n452), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G134), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n460), .A2(new_n469), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G217), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n306), .A2(new_n479), .A3(G953), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT92), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n482));
  INV_X1    g296(.A(new_n480), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n472), .A2(new_n477), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n466), .A2(new_n468), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n459), .B2(new_n456), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n482), .B(new_n483), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT91), .B1(new_n478), .B2(new_n480), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n452), .A2(new_n453), .A3(new_n458), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n458), .B1(new_n452), .B2(new_n453), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n468), .B(new_n466), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  AND4_X1   g306(.A1(KEYINPUT91), .A2(new_n492), .A3(new_n484), .A4(new_n480), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n481), .B(new_n488), .C1(new_n489), .C2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n495));
  NOR2_X1   g309(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n496));
  OAI21_X1  g310(.A(G478), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n494), .A2(new_n374), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n494), .B2(new_n374), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G952), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n502), .A2(G953), .ZN(new_n503));
  NAND2_X1  g317(.A1(G234), .A2(G237), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT21), .B(G898), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n504), .A2(G902), .A3(G953), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT94), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n448), .A2(new_n501), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n305), .A2(new_n373), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G472), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n321), .B1(new_n319), .B2(new_n325), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n327), .A2(new_n320), .A3(new_n328), .ZN(new_n516));
  INV_X1    g330(.A(new_n210), .ZN(new_n517));
  NOR3_X1   g331(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n205), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n204), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n515), .A2(new_n516), .B1(new_n521), .B2(new_n206), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n418), .B1(G134), .B2(G137), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n455), .B2(G137), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n328), .A2(new_n418), .A3(new_n322), .A4(new_n324), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n340), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n522), .A2(new_n526), .A3(new_n236), .ZN(new_n527));
  INV_X1    g341(.A(new_n236), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n336), .B1(new_n326), .B2(new_n329), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n340), .A2(new_n525), .A3(new_n524), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT28), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n528), .A3(new_n530), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n533), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n386), .A2(G210), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT27), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT26), .B(G101), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT29), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n374), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n544), .A2(KEYINPUT69), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n522), .A2(new_n526), .A3(KEYINPUT30), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n529), .B2(new_n530), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n236), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n533), .ZN(new_n550));
  INV_X1    g364(.A(new_n542), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT29), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n533), .A2(new_n535), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n532), .A2(new_n553), .A3(new_n542), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n544), .A2(KEYINPUT69), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n514), .B1(new_n545), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n549), .A2(new_n533), .A3(new_n542), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT31), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n532), .A2(new_n553), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n551), .ZN(new_n561));
  OAI21_X1  g375(.A(KEYINPUT30), .B1(new_n522), .B2(new_n526), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n529), .A2(new_n547), .A3(new_n530), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n527), .B1(new_n564), .B2(new_n236), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n542), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n559), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(KEYINPUT32), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT67), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT32), .B1(new_n568), .B2(new_n569), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n569), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT32), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(KEYINPUT67), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n557), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT77), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n479), .B1(G234), .B2(new_n374), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n411), .A2(new_n414), .ZN(new_n583));
  XNOR2_X1  g397(.A(G119), .B(G128), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT70), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT24), .B(G110), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n230), .A2(G128), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n230), .A2(G128), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(KEYINPUT23), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G110), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT71), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n592), .A2(KEYINPUT71), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n587), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n583), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n376), .A2(new_n380), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n585), .A2(new_n586), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n591), .A2(G110), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n430), .A2(new_n433), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT22), .B(G137), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n596), .A2(new_n601), .A3(new_n605), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n374), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT25), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n607), .A2(KEYINPUT25), .A3(new_n374), .A4(new_n608), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n582), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n596), .A2(new_n601), .A3(new_n605), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n605), .B1(new_n596), .B2(new_n601), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n581), .A2(G902), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT76), .Z(new_n619));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n579), .A2(new_n580), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n566), .B1(new_n565), .B2(new_n542), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n528), .B1(new_n562), .B2(new_n563), .ZN(new_n624));
  NOR4_X1   g438(.A1(new_n624), .A2(KEYINPUT31), .A3(new_n527), .A4(new_n551), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n542), .B1(new_n532), .B2(new_n553), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n569), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n576), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n571), .A3(new_n570), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n556), .B1(new_n630), .B2(new_n577), .ZN(new_n631));
  AOI21_X1  g445(.A(KEYINPUT25), .B1(new_n616), .B2(new_n374), .ZN(new_n632));
  INV_X1    g446(.A(new_n612), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n581), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n620), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT77), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n513), .B1(new_n622), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(G101), .Z(G3));
  AOI21_X1  g453(.A(new_n189), .B1(new_n303), .B2(new_n298), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n188), .B1(new_n640), .B2(KEYINPUT95), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n478), .A2(new_n480), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT33), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n374), .A2(G478), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT96), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT33), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n494), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n646), .B1(new_n494), .B2(new_n647), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n644), .B(new_n645), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT97), .B(G478), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n494), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(G902), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n655), .A2(new_n448), .A3(new_n510), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT95), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n300), .A2(new_n657), .A3(new_n304), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n641), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n641), .A2(new_n656), .A3(new_n658), .A4(KEYINPUT98), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n568), .A2(new_n374), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n664), .A2(G472), .B1(new_n568), .B2(new_n569), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n621), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n372), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT34), .B(G104), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G6));
  NOR3_X1   g484(.A1(new_n448), .A2(new_n500), .A3(new_n511), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n641), .A2(new_n658), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n667), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT99), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT35), .B(G107), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n606), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n602), .B(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n619), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n634), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n681), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT100), .B1(new_n613), .B2(new_n683), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n682), .A2(new_n684), .A3(new_n665), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(new_n512), .A3(new_n305), .A4(new_n373), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT101), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n686), .B(new_n688), .ZN(G12));
  NAND2_X1  g503(.A1(new_n682), .A2(new_n684), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n631), .A2(new_n690), .A3(new_n372), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n641), .A2(new_n658), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n424), .A2(new_n445), .ZN(new_n694));
  INV_X1    g508(.A(new_n443), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT20), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(new_n446), .B1(G475), .B2(new_n426), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n501), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT102), .B(G900), .Z(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(new_n508), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n505), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n693), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G128), .ZN(G30));
  XNOR2_X1  g519(.A(new_n701), .B(KEYINPUT39), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n373), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT40), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n527), .A2(new_n531), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n374), .B1(new_n709), .B2(new_n542), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n550), .A2(new_n542), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n514), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n630), .B2(new_n577), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n613), .A2(new_n683), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n697), .A2(new_n500), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n187), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n300), .A2(new_n304), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(KEYINPUT38), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n708), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n193), .ZN(G45));
  NAND3_X1  g537(.A1(new_n655), .A2(new_n448), .A3(new_n701), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n693), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  NAND2_X1  g541(.A1(new_n630), .A2(new_n577), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n636), .B1(new_n728), .B2(new_n557), .ZN(new_n729));
  INV_X1    g543(.A(new_n370), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n362), .B1(new_n361), .B2(new_n339), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n374), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  INV_X1    g547(.A(G469), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n734), .B(new_n374), .C1(new_n730), .C2(new_n731), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n733), .A2(new_n307), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n661), .B2(new_n662), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT41), .B(G113), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND3_X1  g554(.A1(new_n729), .A2(new_n672), .A3(new_n736), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  AND2_X1   g556(.A1(new_n682), .A2(new_n684), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n579), .A2(new_n743), .A3(new_n512), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n641), .A2(new_n658), .A3(new_n736), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n641), .A2(new_n658), .A3(new_n736), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT103), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n744), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n230), .ZN(G21));
  NAND2_X1  g564(.A1(new_n664), .A2(G472), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n538), .A2(new_n551), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n559), .A3(new_n567), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n569), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n751), .A2(new_n634), .A3(new_n635), .A4(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n733), .A2(new_n510), .A3(new_n307), .A4(new_n735), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n658), .A3(new_n641), .A4(new_n717), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NAND2_X1  g573(.A1(new_n748), .A2(new_n746), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n751), .A2(new_n754), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n716), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n724), .A2(KEYINPUT104), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G125), .ZN(G27));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT105), .B1(new_n366), .B2(new_n371), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n735), .A2(new_n770), .A3(new_n365), .A4(new_n364), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n307), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n300), .A2(new_n187), .A3(new_n304), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n729), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n761), .A2(new_n764), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n768), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n556), .B1(KEYINPUT106), .B2(new_n573), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n570), .A2(KEYINPUT106), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n629), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n636), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n772), .A2(new_n768), .A3(new_n773), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n782), .A3(new_n764), .A4(new_n761), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G131), .ZN(G33));
  NAND3_X1  g599(.A1(new_n729), .A2(new_n774), .A3(new_n703), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  INV_X1    g601(.A(new_n307), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n339), .A2(new_n362), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g604(.A1(new_n790), .A2(new_n361), .B1(new_n348), .B2(new_n352), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT45), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(G469), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT46), .B1(new_n794), .B2(new_n365), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n371), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n365), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n788), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n706), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT107), .ZN(new_n800));
  INV_X1    g614(.A(new_n773), .ZN(new_n801));
  INV_X1    g615(.A(new_n655), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n448), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n804), .A2(KEYINPUT43), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(KEYINPUT43), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n716), .A2(new_n665), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT44), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n801), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n800), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  XNOR2_X1  g627(.A(new_n798), .B(KEYINPUT47), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n773), .A2(new_n724), .A3(new_n621), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n631), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n498), .A2(new_n499), .A3(new_n702), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n697), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n697), .B2(new_n819), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n773), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(new_n373), .A3(new_n579), .A4(new_n743), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n774), .A2(new_n763), .A3(new_n764), .A4(new_n761), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n786), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n777), .B2(new_n783), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n738), .A2(new_n749), .A3(new_n638), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n279), .A2(new_n299), .A3(new_n190), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n187), .B1(new_n828), .B2(new_n640), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n697), .A2(new_n501), .A3(new_n510), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT108), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT108), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n305), .A2(new_n832), .A3(new_n671), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n831), .A2(new_n667), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n741), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n666), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n305), .A3(new_n373), .A4(new_n656), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n686), .A2(new_n758), .A3(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n826), .A2(new_n827), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT110), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n691), .B(new_n692), .C1(new_n703), .C2(new_n725), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n766), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n641), .A2(new_n658), .A3(new_n717), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n716), .A2(new_n701), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n772), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n847), .A3(new_n715), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT111), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n613), .A2(new_n683), .A3(new_n702), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n307), .A3(new_n771), .A4(new_n769), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n714), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n845), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n842), .B1(new_n844), .B2(new_n855), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n853), .A2(new_n845), .A3(new_n847), .A4(new_n715), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n852), .B2(new_n845), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .A3(new_n766), .A4(new_n843), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n840), .A2(new_n841), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT110), .A4(new_n839), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT53), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n513), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n622), .A2(new_n637), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n579), .A2(new_n621), .A3(new_n736), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n864), .A2(new_n865), .B1(new_n663), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n749), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n839), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n825), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n784), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n856), .A2(new_n860), .ZN(new_n873));
  XOR2_X1   g687(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(KEYINPUT54), .B1(new_n863), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n856), .A2(new_n860), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n874), .B1(new_n879), .B2(new_n840), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT113), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n880), .A2(new_n885), .A3(new_n881), .A4(new_n882), .ZN(new_n886));
  INV_X1    g700(.A(new_n505), .ZN(new_n887));
  INV_X1    g701(.A(new_n755), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n805), .A2(new_n887), .A3(new_n888), .A4(new_n806), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n773), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n733), .A2(new_n735), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(new_n788), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n814), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n721), .A2(new_n188), .A3(new_n736), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT50), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n894), .A2(new_n889), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n894), .B2(new_n889), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n801), .A2(new_n736), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT114), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n714), .A2(new_n887), .A3(new_n621), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n655), .A2(new_n448), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n805), .A2(new_n887), .A3(new_n806), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n902), .A2(new_n903), .B1(new_n905), .B2(new_n763), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n893), .A2(new_n898), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT51), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n893), .A2(new_n898), .A3(KEYINPUT51), .A4(new_n906), .ZN(new_n910));
  INV_X1    g724(.A(new_n781), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n900), .A2(new_n904), .A3(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT48), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n802), .A2(new_n697), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n902), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n760), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n915), .B(new_n503), .C1(new_n916), .C2(new_n889), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n909), .A2(new_n910), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n878), .A2(new_n884), .A3(new_n886), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT115), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n841), .B1(new_n869), .B2(new_n871), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n922), .A2(new_n873), .A3(new_n862), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n876), .ZN(new_n926));
  AOI22_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .B1(new_n883), .B2(KEYINPUT113), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n927), .A2(new_n928), .A3(new_n886), .A4(new_n919), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n502), .A2(new_n216), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n921), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n891), .B(KEYINPUT49), .Z(new_n932));
  NOR2_X1   g746(.A1(new_n932), .A2(new_n804), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n636), .A2(new_n188), .A3(new_n788), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n714), .A3(new_n721), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n931), .A2(new_n935), .ZN(G75));
  AOI21_X1  g750(.A(new_n374), .B1(new_n880), .B2(new_n882), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(G210), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(KEYINPUT117), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(KEYINPUT117), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n301), .A2(new_n302), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n221), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n303), .ZN(new_n943));
  XOR2_X1   g757(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n945), .A2(KEYINPUT56), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n940), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n216), .A2(G952), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n938), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n948), .B1(new_n950), .B2(new_n945), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n947), .A2(new_n951), .ZN(G51));
  XOR2_X1   g766(.A(new_n794), .B(KEYINPUT119), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n937), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n365), .B(KEYINPUT57), .Z(new_n956));
  AND3_X1   g770(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT53), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n875), .B1(new_n872), .B2(new_n873), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT54), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n730), .A2(new_n731), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n955), .B1(new_n964), .B2(KEYINPUT118), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT118), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n961), .A2(new_n966), .A3(new_n963), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n948), .B1(new_n965), .B2(new_n967), .ZN(G54));
  INV_X1    g782(.A(new_n948), .ZN(new_n969));
  NAND2_X1  g783(.A1(KEYINPUT58), .A2(G475), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n937), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n969), .B1(new_n973), .B2(new_n442), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n442), .B2(new_n973), .ZN(G60));
  OR2_X1    g789(.A1(new_n648), .A2(new_n649), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n976), .A2(new_n644), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n878), .A2(new_n884), .A3(new_n886), .ZN(new_n978));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT59), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT120), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n977), .B(new_n980), .C1(new_n959), .C2(new_n960), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n969), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n977), .A2(new_n980), .ZN(new_n985));
  OAI21_X1  g799(.A(KEYINPUT54), .B1(new_n957), .B2(new_n958), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n985), .B1(new_n986), .B2(new_n883), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n987), .A2(KEYINPUT120), .A3(new_n948), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n981), .A2(new_n984), .A3(new_n988), .ZN(G63));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT121), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n957), .B2(new_n958), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n948), .B1(new_n993), .B2(new_n617), .ZN(new_n994));
  INV_X1    g808(.A(new_n679), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n994), .B1(new_n995), .B2(new_n993), .ZN(new_n996));
  XNOR2_X1  g810(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G66));
  AOI21_X1  g812(.A(new_n216), .B1(new_n507), .B2(G224), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT123), .Z(new_n1000));
  INV_X1    g814(.A(new_n869), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1000), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT124), .Z(new_n1003));
  OAI21_X1  g817(.A(new_n941), .B1(G898), .B2(new_n216), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  XOR2_X1   g819(.A(new_n564), .B(new_n435), .Z(new_n1006));
  AND2_X1   g820(.A1(new_n816), .A2(new_n786), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n781), .A2(new_n845), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n800), .B1(new_n811), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n844), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n1007), .A2(new_n1009), .A3(new_n784), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(G953), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n350), .A2(KEYINPUT126), .A3(G900), .ZN(new_n1013));
  OAI21_X1  g827(.A(G953), .B1(KEYINPUT126), .B2(G900), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n1006), .B(new_n1012), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n844), .A2(new_n722), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1018), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT125), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1020));
  OAI221_X1 g834(.A(new_n816), .B1(KEYINPUT62), .B2(new_n1018), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n914), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n773), .B(new_n707), .C1(new_n1022), .C2(new_n698), .ZN(new_n1023));
  AOI22_X1  g837(.A1(new_n800), .A2(new_n811), .B1(new_n865), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n216), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1017), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1016), .B1(new_n1026), .B2(new_n1006), .ZN(G72));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  OAI21_X1  g843(.A(new_n1029), .B1(new_n1011), .B2(new_n869), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n550), .A2(new_n542), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n948), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(new_n926), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1031), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1034), .A2(new_n712), .A3(new_n1029), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1032), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1024), .A2(new_n1001), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1029), .B1(new_n1021), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n712), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OR2_X1    g854(.A1(new_n1040), .A2(KEYINPUT127), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1040), .A2(KEYINPUT127), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(G57));
endmodule


