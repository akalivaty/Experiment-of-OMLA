//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(G228gat), .ZN(new_n205));
  INV_X1    g004(.A(G233gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  AND2_X1   g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G197gat), .A2(G204gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n211), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G211gat), .B(G218gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(G197gat), .B(G204gat), .ZN(new_n218));
  INV_X1    g017(.A(new_n215), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT71), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n216), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT71), .B(new_n211), .C1(new_n214), .C2(new_n215), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G155gat), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G162gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g031(.A(G141gat), .B(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n236), .A2(G148gat), .ZN(new_n237));
  INV_X1    g036(.A(G148gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(G141gat), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT74), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n231), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(G148gat), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n237), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n231), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT2), .B1(new_n249), .B2(new_n227), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n241), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n225), .B1(new_n226), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n216), .A2(new_n220), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT3), .B1(new_n255), .B2(new_n226), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n233), .A2(new_n234), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT74), .B1(new_n237), .B2(new_n239), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n232), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n259), .A2(new_n231), .B1(new_n246), .B2(new_n250), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n208), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n222), .A2(new_n226), .A3(new_n223), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT81), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT81), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n222), .A2(new_n265), .A3(new_n226), .A4(new_n223), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n252), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n241), .A2(new_n251), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n226), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n253), .A2(KEYINPUT83), .A3(new_n226), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n273), .A2(new_n224), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n270), .A2(new_n275), .A3(new_n207), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n204), .B(new_n262), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n267), .A2(new_n269), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT82), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n225), .B1(new_n271), .B2(new_n272), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n208), .B1(new_n282), .B2(new_n274), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n283), .A3(new_n270), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n204), .B1(new_n284), .B2(new_n262), .ZN(new_n285));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286));
  XOR2_X1   g085(.A(new_n286), .B(KEYINPUT80), .Z(new_n287));
  NOR3_X1   g086(.A1(new_n279), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n287), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n262), .B1(new_n276), .B2(new_n277), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G22gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n289), .B1(new_n291), .B2(new_n278), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n203), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n287), .B1(new_n279), .B2(new_n285), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n291), .A2(new_n289), .A3(new_n278), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n202), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G1gat), .B(G29gat), .Z(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT78), .B(KEYINPUT0), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G57gat), .B(G85gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G225gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G127gat), .B(G134gat), .Z(new_n306));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n306), .B(KEYINPUT68), .C1(KEYINPUT1), .C2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n309));
  INV_X1    g108(.A(G113gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G120gat), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G113gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT1), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT69), .ZN(new_n317));
  OR3_X1    g116(.A1(new_n312), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n315), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n308), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(KEYINPUT3), .B2(new_n269), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n305), .B1(new_n322), .B2(new_n253), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n316), .A3(new_n320), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT79), .B(KEYINPUT4), .C1(new_n269), .C2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT4), .B1(new_n269), .B2(new_n325), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n321), .A2(new_n260), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT79), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n323), .A2(new_n324), .A3(new_n326), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n329), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n325), .A3(new_n253), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n304), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(KEYINPUT77), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n323), .B2(new_n333), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n260), .B(new_n325), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT5), .B1(new_n341), .B2(new_n304), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n303), .B(new_n332), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n336), .A2(KEYINPUT77), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n323), .A2(new_n338), .A3(new_n333), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n332), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n302), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT6), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n343), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(KEYINPUT6), .B(new_n302), .C1(new_n346), .C2(new_n347), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(G169gat), .ZN(new_n358));
  INV_X1    g157(.A(G176gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT23), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n363), .A2(KEYINPUT23), .A3(new_n358), .A4(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n356), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n367), .B1(new_n369), .B2(KEYINPUT23), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n356), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT65), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n356), .A2(KEYINPUT65), .A3(new_n362), .A4(new_n370), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  XOR2_X1   g175(.A(KEYINPUT27), .B(G183gat), .Z(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n377), .B2(G190gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT67), .B(KEYINPUT28), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n376), .B(new_n379), .C1(new_n377), .C2(G190gat), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n360), .A2(KEYINPUT26), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n357), .B1(new_n360), .B2(KEYINPUT26), .ZN(new_n384));
  AOI22_X1  g183(.A1(new_n383), .A2(new_n384), .B1(G183gat), .B2(G190gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G226gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(new_n206), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n375), .B2(new_n386), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(new_n225), .C1(new_n389), .C2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n389), .B1(new_n387), .B2(new_n226), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n389), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n375), .B2(new_n386), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n393), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n392), .B1(new_n399), .B2(new_n225), .ZN(new_n400));
  XOR2_X1   g199(.A(G8gat), .B(G36gat), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT73), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n404), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n392), .B(new_n406), .C1(new_n399), .C2(new_n225), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(KEYINPUT30), .A3(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n393), .A2(new_n224), .A3(new_n397), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n397), .A2(KEYINPUT72), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n394), .B(new_n396), .C1(new_n375), .C2(new_n386), .ZN(new_n411));
  OAI22_X1  g210(.A1(new_n410), .A2(new_n411), .B1(new_n389), .B2(new_n391), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n412), .B2(new_n224), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n406), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n350), .A2(new_n351), .B1(new_n408), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n297), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n387), .A2(new_n321), .ZN(new_n418));
  INV_X1    g217(.A(G227gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n206), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n375), .A2(new_n325), .A3(new_n386), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT32), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G15gat), .B(G43gat), .Z(new_n426));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n422), .B(KEYINPUT32), .C1(new_n424), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT34), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n420), .B1(new_n418), .B2(new_n421), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT70), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n429), .A2(new_n431), .A3(new_n436), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n438), .A2(new_n435), .A3(new_n434), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n434), .A2(new_n435), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n429), .A2(new_n431), .A3(new_n436), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n436), .B1(new_n429), .B2(new_n431), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT36), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n444), .A3(KEYINPUT36), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n417), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n407), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT37), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n406), .B1(new_n413), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n412), .A2(new_n225), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n393), .A2(new_n397), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n455), .B2(new_n224), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT38), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n451), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n392), .B(new_n452), .C1(new_n399), .C2(new_n225), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n404), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n412), .A2(new_n224), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n452), .B1(new_n461), .B2(new_n392), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT38), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n458), .A2(new_n463), .A3(new_n350), .A4(new_n351), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n331), .A2(new_n335), .A3(new_n326), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n305), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT39), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n341), .B2(new_n304), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n467), .A3(new_n305), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n469), .A2(KEYINPUT40), .A3(new_n303), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n348), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n469), .A2(new_n303), .A3(new_n470), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT40), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n472), .A2(new_n415), .A3(new_n408), .A4(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n294), .A2(new_n202), .A3(new_n295), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n202), .B1(new_n294), .B2(new_n295), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n464), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n416), .B(new_n445), .C1(new_n477), .C2(new_n478), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n297), .A2(new_n482), .A3(new_n416), .A4(new_n445), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n450), .A2(new_n479), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT84), .ZN(new_n485));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G197gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT11), .B(G169gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n487), .B(new_n488), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT12), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  OR2_X1    g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(G43gat), .A2(G50gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n492), .B1(new_n495), .B2(KEYINPUT85), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT85), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n493), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G29gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n500), .A2(KEYINPUT14), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n500), .B2(KEYINPUT14), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n493), .A2(new_n492), .A3(new_n494), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n496), .A2(new_n498), .A3(new_n505), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n491), .B1(new_n510), .B2(KEYINPUT17), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n508), .A2(KEYINPUT86), .A3(new_n512), .A4(new_n509), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(G1gat), .ZN(new_n517));
  AND2_X1   g316(.A1(new_n517), .A2(KEYINPUT87), .ZN(new_n518));
  XOR2_X1   g317(.A(G15gat), .B(G22gat), .Z(new_n519));
  INV_X1    g318(.A(G1gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n517), .B2(KEYINPUT87), .ZN(new_n522));
  OAI21_X1  g321(.A(G8gat), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n517), .A2(KEYINPUT88), .ZN(new_n524));
  INV_X1    g323(.A(G8gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n515), .B(new_n526), .C1(new_n516), .C2(G1gat), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n524), .A2(new_n525), .A3(new_n521), .A4(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n510), .A2(KEYINPUT17), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n523), .A2(new_n528), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(new_n508), .A3(new_n509), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n532), .B(KEYINPUT13), .Z(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n510), .A2(new_n523), .A3(new_n537), .A4(new_n528), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n529), .B2(new_n510), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n529), .A2(new_n510), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n511), .A2(new_n513), .B1(KEYINPUT17), .B2(new_n510), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(new_n529), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT18), .B1(new_n545), .B2(new_n532), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n485), .B(new_n490), .C1(new_n542), .C2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n535), .A3(new_n541), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n490), .B1(new_n552), .B2(new_n485), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT90), .Z(new_n557));
  XOR2_X1   g356(.A(G57gat), .B(G64gat), .Z(new_n558));
  AOI22_X1  g357(.A1(new_n558), .A2(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G57gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G64gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n556), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n557), .A2(new_n559), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(G127gat), .Z(new_n572));
  OAI21_X1  g371(.A(new_n529), .B1(new_n568), .B2(new_n567), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n574), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT92), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT92), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(G85gat), .A3(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n584), .A3(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT8), .ZN(new_n590));
  OR2_X1    g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n590), .A2(KEYINPUT93), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT93), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n587), .B(new_n588), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G99gat), .B(G106gat), .Z(new_n595));
  OAI21_X1  g394(.A(new_n580), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n592), .A2(new_n593), .ZN(new_n597));
  INV_X1    g396(.A(new_n588), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT7), .B1(new_n582), .B2(new_n584), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n595), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n597), .A2(new_n600), .A3(KEYINPUT94), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n594), .A2(new_n595), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n594), .A2(KEYINPUT95), .A3(new_n595), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n510), .ZN(new_n609));
  AND2_X1   g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n609), .B1(KEYINPUT41), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n544), .A2(KEYINPUT96), .A3(new_n608), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT96), .B1(new_n544), .B2(new_n608), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G190gat), .B(G218gat), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G134gat), .B(G162gat), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n615), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n611), .B(new_n620), .C1(new_n612), .C2(new_n613), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n616), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n619), .B1(new_n616), .B2(new_n621), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n579), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n566), .A2(KEYINPUT10), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n608), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n604), .A3(new_n566), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT97), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT97), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n629), .A2(new_n604), .A3(new_n566), .A4(new_n632), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n608), .A2(new_n567), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G230gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT98), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n636), .A2(new_n638), .B1(new_n637), .B2(new_n634), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n608), .A2(new_n567), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n631), .A2(new_n633), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n635), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n628), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n637), .ZN(new_n650));
  INV_X1    g449(.A(new_n634), .ZN(new_n651));
  INV_X1    g450(.A(new_n637), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n643), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n644), .A2(new_n654), .ZN(new_n655));
  NOR4_X1   g454(.A1(new_n484), .A2(new_n555), .A3(new_n626), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n350), .A2(new_n351), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT99), .B(G1gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n408), .A2(new_n415), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  AND2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n664), .A2(new_n525), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT42), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(KEYINPUT42), .B2(new_n666), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n656), .A2(new_n670), .A3(new_n445), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n656), .A2(new_n449), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n670), .ZN(G1326gat));
  INV_X1    g472(.A(new_n297), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT100), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  NAND2_X1  g477(.A1(new_n481), .A2(new_n483), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n440), .A2(new_n444), .A3(KEYINPUT36), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT36), .B1(new_n440), .B2(new_n444), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n657), .A2(new_n662), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n296), .A3(new_n293), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n479), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n625), .B1(new_n679), .B2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n579), .A2(new_n555), .A3(new_n655), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n500), .A3(new_n658), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT101), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n293), .A2(new_n296), .B1(new_n440), .B2(new_n444), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n482), .B1(new_n692), .B2(new_n416), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n685), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n695), .A2(new_n624), .B1(KEYINPUT102), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n698));
  AOI211_X1 g497(.A(new_n625), .B(new_n698), .C1(new_n679), .C2(new_n685), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n687), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n657), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n691), .A2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n663), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n503), .B1(new_n705), .B2(KEYINPUT103), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(KEYINPUT103), .B2(new_n705), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n503), .A3(new_n663), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT46), .Z(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(G1329gat));
  NAND2_X1  g509(.A1(new_n704), .A2(new_n449), .ZN(new_n711));
  INV_X1    g510(.A(new_n445), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(G43gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n711), .A2(G43gat), .B1(new_n688), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g514(.A1(new_n704), .A2(G50gat), .A3(new_n674), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n688), .A2(new_n674), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(G50gat), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT48), .ZN(G1331gat));
  AOI22_X1  g518(.A1(new_n639), .A2(new_n643), .B1(new_n650), .B2(new_n653), .ZN(new_n720));
  NOR4_X1   g519(.A1(new_n484), .A2(new_n554), .A3(new_n626), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n658), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n663), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT49), .B(G64gat), .Z(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(G1333gat));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n449), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n712), .A2(G71gat), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n728), .A2(G71gat), .B1(new_n721), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n721), .A2(new_n674), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n579), .A2(new_n554), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n720), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n697), .B2(new_n699), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n739), .B(new_n736), .C1(new_n697), .C2(new_n699), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n738), .A2(new_n658), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(G85gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n695), .A2(new_n744), .A3(new_n624), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n734), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n686), .A2(new_n744), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n735), .B1(new_n686), .B2(new_n744), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT105), .B1(new_n484), .B2(new_n625), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT51), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n658), .A2(new_n742), .A3(new_n655), .ZN(new_n754));
  OAI22_X1  g553(.A1(new_n741), .A2(new_n742), .B1(new_n753), .B2(new_n754), .ZN(G1336gat));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n738), .A2(new_n663), .A3(new_n740), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G92gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n749), .A2(new_n750), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n743), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n761), .A3(KEYINPUT51), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n662), .A2(G92gat), .A3(new_n720), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n757), .B1(new_n759), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G92gat), .B1(new_n737), .B2(new_n662), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n757), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n749), .A2(KEYINPUT51), .A3(new_n750), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n749), .B2(new_n750), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT107), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n752), .A2(new_n774), .A3(new_n765), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n769), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n756), .B1(new_n767), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n769), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n774), .B1(new_n752), .B2(new_n765), .ZN(new_n779));
  INV_X1    g578(.A(new_n765), .ZN(new_n780));
  AOI211_X1 g579(.A(KEYINPUT107), .B(new_n780), .C1(new_n748), .C2(new_n751), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT51), .B1(new_n760), .B2(new_n761), .ZN(new_n783));
  AOI211_X1 g582(.A(KEYINPUT106), .B(new_n743), .C1(new_n749), .C2(new_n750), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n785), .A2(new_n765), .B1(new_n758), .B2(G92gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n782), .B(KEYINPUT108), .C1(new_n757), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n777), .A2(new_n787), .ZN(G1337gat));
  NAND3_X1  g587(.A1(new_n738), .A2(new_n449), .A3(new_n740), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT109), .B(G99gat), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n712), .A2(new_n720), .A3(new_n790), .ZN(new_n792));
  XOR2_X1   g591(.A(new_n792), .B(KEYINPUT110), .Z(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n753), .B2(new_n793), .ZN(G1338gat));
  NOR3_X1   g593(.A1(new_n297), .A2(G106gat), .A3(new_n720), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n763), .A2(new_n764), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n785), .A2(KEYINPUT111), .A3(new_n795), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n738), .A2(new_n674), .A3(new_n740), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(G106gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n700), .A2(new_n674), .A3(new_n736), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n804), .B2(G106gat), .ZN(new_n805));
  INV_X1    g604(.A(new_n795), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n753), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n803), .A2(new_n807), .ZN(G1339gat));
  INV_X1    g607(.A(new_n579), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT54), .B1(new_n636), .B2(new_n652), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n647), .A2(new_n648), .A3(new_n638), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT112), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n636), .A2(new_n638), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n650), .A2(new_n813), .A3(new_n814), .A4(KEYINPUT54), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n636), .A2(new_n638), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n642), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n812), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n812), .A2(new_n818), .A3(new_n815), .A4(KEYINPUT55), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n821), .A2(new_n554), .A3(new_n654), .A4(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n551), .A2(new_n535), .A3(new_n541), .A4(new_n490), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n545), .A2(new_n532), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n539), .A2(new_n540), .A3(new_n536), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n489), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n824), .B1(new_n830), .B2(new_n655), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n720), .A2(new_n829), .A3(KEYINPUT113), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n624), .B1(new_n823), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n821), .A2(new_n654), .A3(new_n822), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n624), .A2(new_n830), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n809), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n579), .A2(new_n555), .A3(new_n625), .A4(new_n720), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n657), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n692), .A2(new_n662), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(new_n555), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(new_n310), .ZN(G1340gat));
  NOR2_X1   g644(.A1(new_n843), .A2(new_n720), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(new_n312), .ZN(G1341gat));
  NOR2_X1   g646(.A1(new_n843), .A2(new_n809), .ZN(new_n848));
  NOR2_X1   g647(.A1(KEYINPUT114), .A2(G127gat), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(G1342gat));
  NAND3_X1  g649(.A1(new_n840), .A2(new_n624), .A3(new_n842), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n851), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT56), .B1(new_n851), .B2(G134gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(G134gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(G1343gat));
  AOI21_X1  g654(.A(new_n297), .B1(new_n838), .B2(new_n839), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT57), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n830), .A2(new_n655), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n624), .B1(new_n823), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n809), .B1(new_n859), .B2(new_n837), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n297), .B1(new_n860), .B2(new_n839), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n861), .B2(KEYINPUT57), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n839), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(KEYINPUT115), .A3(KEYINPUT57), .A4(new_n674), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n449), .A2(new_n657), .A3(new_n663), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n863), .A2(new_n868), .A3(new_n554), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n242), .A2(new_n243), .ZN(new_n870));
  AND4_X1   g669(.A1(new_n674), .A2(new_n840), .A3(new_n662), .A4(new_n682), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n555), .A2(G141gat), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n873), .A2(KEYINPUT116), .A3(KEYINPUT58), .ZN(new_n874));
  NOR2_X1   g673(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n875));
  AND2_X1   g674(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(new_n877), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n871), .A2(new_n238), .A3(new_n655), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n838), .A2(new_n839), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .A3(new_n674), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n882), .B(KEYINPUT117), .C1(KEYINPUT57), .C2(new_n861), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n856), .A2(new_n884), .A3(KEYINPUT57), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n883), .A2(new_n655), .A3(new_n866), .A4(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n880), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n880), .A2(G148gat), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n867), .B1(new_n857), .B2(new_n862), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n655), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n879), .B1(new_n887), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n893), .B(new_n879), .C1(new_n887), .C2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n894), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n871), .A2(new_n249), .A3(new_n579), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n889), .A2(new_n579), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n249), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n871), .B2(new_n624), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n625), .A2(new_n227), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n889), .B2(new_n900), .ZN(G1347gat));
  AND2_X1   g700(.A1(new_n692), .A2(new_n663), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n881), .A2(new_n657), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n554), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n358), .A2(KEYINPUT119), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n358), .A2(KEYINPUT119), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n904), .B2(new_n905), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n363), .A2(new_n364), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n903), .A2(new_n909), .A3(new_n655), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n903), .A2(new_n655), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(KEYINPUT120), .A3(new_n359), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT120), .B1(new_n913), .B2(new_n359), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n911), .A2(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n916), .B(new_n917), .ZN(G1349gat));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n377), .A3(new_n579), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(G183gat), .B1(new_n903), .B2(new_n579), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n658), .B1(new_n838), .B2(new_n839), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n902), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n926), .A2(new_n809), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n920), .B(KEYINPUT123), .C1(G183gat), .C2(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT60), .A4(new_n928), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n923), .A2(KEYINPUT60), .A3(new_n928), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n921), .A2(new_n922), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT124), .B1(new_n931), .B2(KEYINPUT60), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(G1350gat));
  NOR2_X1   g733(.A1(new_n926), .A2(new_n625), .ZN(new_n935));
  NAND2_X1  g734(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g736(.A(KEYINPUT61), .B(G190gat), .Z(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n935), .B2(new_n938), .ZN(G1351gat));
  XOR2_X1   g738(.A(KEYINPUT125), .B(G197gat), .Z(new_n940));
  NOR3_X1   g739(.A1(new_n449), .A2(new_n658), .A3(new_n662), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n883), .A2(new_n885), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n940), .B1(new_n942), .B2(new_n555), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n449), .A2(new_n297), .A3(new_n662), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n925), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n555), .A2(new_n940), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(G1352gat));
  NOR3_X1   g746(.A1(new_n945), .A2(G204gat), .A3(new_n720), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT62), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n883), .A2(new_n655), .A3(new_n885), .A4(new_n941), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G204gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT126), .ZN(G1353gat));
  INV_X1    g752(.A(G211gat), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(KEYINPUT127), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n956), .B1(new_n942), .B2(new_n809), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n955), .A2(KEYINPUT127), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  INV_X1    g759(.A(new_n945), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n954), .A3(new_n579), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(G218gat), .B1(new_n942), .B2(new_n625), .ZN(new_n964));
  OR3_X1    g763(.A1(new_n945), .A2(G218gat), .A3(new_n625), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1355gat));
endmodule


