//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n906, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1046, new_n1047;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT22), .ZN(new_n207));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT22), .ZN(new_n212));
  NAND2_X1  g011(.A1(G211gat), .A2(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(G197gat), .ZN(new_n214));
  INV_X1    g013(.A(G204gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G197gat), .A2(G204gat), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n212), .A2(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n209), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  OR2_X1    g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G141gat), .B(G148gat), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n221), .B(new_n222), .C1(new_n223), .C2(KEYINPUT2), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  INV_X1    g024(.A(G141gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G148gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT71), .B(G148gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(G141gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231));
  INV_X1    g030(.A(G155gat), .ZN(new_n232));
  INV_X1    g031(.A(G162gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n234), .A2(new_n221), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n224), .B(new_n225), .C1(new_n230), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n220), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G228gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(KEYINPUT71), .A2(G148gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT71), .A2(G148gat), .ZN(new_n243));
  OAI21_X1  g042(.A(G141gat), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n244), .A2(new_n227), .B1(new_n221), .B2(new_n234), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n221), .ZN(new_n246));
  INV_X1    g045(.A(G148gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G141gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n227), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n231), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n220), .B2(new_n237), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n239), .B(new_n241), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n209), .A2(new_n219), .A3(KEYINPUT77), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT77), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(new_n218), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT78), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT78), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n259), .B(new_n256), .C1(new_n220), .C2(new_n255), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n225), .A3(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n224), .B1(new_n230), .B2(new_n235), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n238), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n263), .B2(new_n241), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n205), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT79), .B(new_n253), .C1(new_n263), .C2(new_n241), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G22gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n260), .A2(new_n225), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n218), .B1(new_n207), .B2(new_n208), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT77), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n259), .B1(new_n271), .B2(new_n256), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n262), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n239), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n240), .ZN(new_n275));
  INV_X1    g074(.A(G22gat), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n275), .A2(KEYINPUT79), .A3(new_n276), .A4(new_n253), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n266), .A2(new_n268), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n264), .A2(new_n265), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n268), .A2(new_n277), .B1(new_n279), .B2(new_n204), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G183gat), .B2(G190gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT25), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT65), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n286), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n292), .B1(new_n295), .B2(new_n287), .ZN(new_n296));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT24), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n299), .A2(new_n302), .A3(new_n282), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n296), .A2(new_n303), .A3(new_n304), .A4(KEYINPUT25), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n291), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n299), .A2(KEYINPUT64), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n307), .A2(new_n302), .A3(new_n282), .A4(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT25), .B1(new_n310), .B2(new_n296), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT66), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n296), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT25), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n315), .A2(new_n316), .A3(new_n291), .A4(new_n305), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT27), .B(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n301), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(KEYINPUT28), .A3(new_n301), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n292), .B1(new_n325), .B2(new_n293), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n325), .B2(new_n293), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n297), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n318), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(G113gat), .A2(G120gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n331));
  NAND2_X1  g130(.A1(G113gat), .A2(G120gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT67), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n329), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G227gat), .ZN(new_n342));
  INV_X1    g141(.A(G233gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n328), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n312), .B2(new_n317), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n336), .B1(new_n333), .B2(new_n334), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n341), .A2(new_n344), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G15gat), .B(G43gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(G71gat), .B(G99gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n346), .A2(new_n349), .ZN(new_n358));
  AOI211_X1 g157(.A(new_n340), .B(new_n345), .C1(new_n312), .C2(new_n317), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT34), .B1(new_n360), .B2(new_n344), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(KEYINPUT32), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT34), .ZN(new_n363));
  INV_X1    g162(.A(new_n344), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n363), .B(new_n364), .C1(new_n358), .C2(new_n359), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n361), .B2(new_n365), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n357), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n350), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n369), .B2(new_n364), .ZN(new_n370));
  INV_X1    g169(.A(new_n365), .ZN(new_n371));
  OAI211_X1 g170(.A(KEYINPUT32), .B(new_n351), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n357), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(KEYINPUT80), .B(KEYINPUT35), .Z(new_n376));
  AND4_X1   g175(.A1(new_n281), .A2(new_n368), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n329), .B2(new_n237), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n328), .B1(new_n306), .B2(new_n311), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n379), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT68), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n381), .A2(KEYINPUT68), .A3(new_n379), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n270), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n318), .A2(new_n379), .A3(new_n328), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n378), .A2(new_n237), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n315), .A2(new_n291), .A3(new_n305), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n328), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT69), .A3(new_n220), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n391), .B1(new_n346), .B2(new_n379), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n270), .ZN(new_n397));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398));
  INV_X1    g197(.A(G64gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G92gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n387), .A2(new_n394), .A3(new_n397), .A4(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT69), .B1(new_n393), .B2(new_n220), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n396), .A2(new_n395), .A3(new_n270), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n403), .B1(new_n409), .B2(new_n387), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n409), .A2(KEYINPUT70), .A3(new_n387), .A4(new_n403), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT70), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n404), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n414), .A3(new_n405), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT0), .B(G57gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G85gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(G1gat), .B(G29gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT3), .B1(new_n245), .B2(new_n250), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n349), .A3(new_n236), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n423), .B(KEYINPUT72), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n340), .A2(new_n251), .A3(KEYINPUT4), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT73), .B1(new_n349), .B2(new_n262), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT73), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n340), .A2(new_n251), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n427), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT74), .ZN(new_n434));
  XOR2_X1   g233(.A(KEYINPUT75), .B(KEYINPUT5), .Z(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n428), .B(new_n430), .C1(new_n340), .C2(new_n251), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n424), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT74), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n426), .A2(new_n432), .A3(new_n439), .A4(new_n427), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n434), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n349), .A2(new_n262), .A3(KEYINPUT73), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n429), .B1(new_n340), .B2(new_n251), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT4), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n431), .B1(new_n349), .B2(new_n262), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n424), .A2(new_n435), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n422), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT76), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n422), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n430), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(KEYINPUT4), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n452), .A2(KEYINPUT76), .A3(new_n445), .A4(new_n446), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n420), .B1(new_n441), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n438), .A3(new_n440), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(new_n419), .A3(new_n449), .A4(new_n453), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n449), .A3(new_n453), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(KEYINPUT6), .A3(new_n420), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n411), .A2(new_n415), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n377), .A2(new_n463), .A3(KEYINPUT81), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n411), .A2(new_n415), .A3(new_n462), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n368), .A2(new_n281), .A3(new_n375), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT35), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT81), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n368), .A2(new_n281), .A3(new_n375), .A4(new_n376), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n468), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n445), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n424), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n419), .B1(new_n473), .B2(KEYINPUT39), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n437), .A2(new_n424), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(KEYINPUT39), .B2(new_n476), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n477), .A2(KEYINPUT40), .B1(new_n420), .B2(new_n460), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(KEYINPUT40), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n412), .A2(new_n414), .A3(new_n405), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n394), .A2(new_n397), .ZN(new_n481));
  INV_X1    g280(.A(new_n386), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n378), .B1(new_n346), .B2(KEYINPUT29), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n220), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n402), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n405), .B2(new_n404), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n478), .B(new_n479), .C1(new_n480), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n387), .A2(new_n488), .A3(new_n394), .A4(new_n397), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n220), .B1(new_n380), .B2(new_n386), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n393), .A2(new_n270), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT37), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n402), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT37), .B1(new_n481), .B2(new_n484), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n496), .A2(KEYINPUT38), .A3(new_n402), .A4(new_n489), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n462), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n412), .A2(new_n414), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n487), .A2(new_n501), .A3(new_n281), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n368), .A2(KEYINPUT36), .A3(new_n375), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504));
  NOR3_X1   g303(.A1(new_n366), .A2(new_n367), .A3(new_n357), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n373), .B1(new_n372), .B2(new_n374), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n281), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n503), .A2(new_n507), .B1(new_n465), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n502), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n471), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n471), .A2(new_n510), .A3(KEYINPUT82), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G15gat), .A2(G22gat), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(G15gat), .A2(G22gat), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT85), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n520));
  INV_X1    g319(.A(G15gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n276), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  OAI22_X1  g323(.A1(new_n519), .A2(new_n523), .B1(new_n524), .B2(G1gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT85), .B1(new_n517), .B2(new_n518), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n520), .A3(new_n516), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(KEYINPUT86), .A3(new_n529), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(G8gat), .C1(KEYINPUT86), .C2(new_n529), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n532), .B1(new_n525), .B2(new_n529), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n526), .A2(new_n527), .B1(KEYINPUT16), .B2(new_n528), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(KEYINPUT87), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT88), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n533), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT87), .B1(new_n539), .B2(new_n535), .ZN(new_n540));
  AOI21_X1  g339(.A(G8gat), .B1(new_n525), .B2(new_n532), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT88), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n531), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G50gat), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(G43gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(G43gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(KEYINPUT15), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(KEYINPUT83), .A2(G43gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(KEYINPUT83), .A2(G43gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT15), .B1(new_n550), .B2(new_n545), .ZN(new_n551));
  INV_X1    g350(.A(G29gat), .ZN(new_n552));
  INV_X1    g351(.A(G36gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT14), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT14), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n554), .B(new_n556), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n547), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n547), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT84), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n558), .A2(KEYINPUT84), .A3(KEYINPUT17), .A4(new_n559), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n537), .B1(new_n533), .B2(new_n536), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n540), .A2(new_n541), .A3(KEYINPUT88), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n570), .A3(new_n531), .ZN(new_n571));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n562), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n572), .B(KEYINPUT13), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n543), .A2(new_n561), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n560), .B1(new_n570), .B2(new_n531), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n562), .A2(new_n571), .A3(KEYINPUT18), .A4(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT11), .B(G169gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(G197gat), .ZN(new_n584));
  XOR2_X1   g383(.A(G113gat), .B(G141gat), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT12), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n575), .A2(new_n587), .A3(new_n580), .A4(new_n581), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n515), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT94), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT91), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n594), .A2(G85gat), .A3(G92gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT7), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n594), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(new_n401), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT92), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT92), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(G99gat), .A3(G106gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT8), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n599), .A2(new_n601), .A3(new_n603), .A4(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n608), .A2(new_n603), .A3(new_n597), .A4(new_n598), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n600), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n611), .A3(KEYINPUT93), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n613), .A3(new_n600), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n593), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(new_n593), .A3(new_n614), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n567), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n612), .A2(new_n593), .A3(new_n614), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n561), .B1(new_n619), .B2(new_n615), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT89), .Z(new_n623));
  INV_X1    g422(.A(KEYINPUT41), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n618), .A2(new_n620), .A3(new_n621), .A4(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G134gat), .B(G162gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT90), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n624), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n625), .A3(new_n620), .ZN(new_n634));
  INV_X1    g433(.A(new_n621), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n626), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n633), .A2(new_n637), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G230gat), .A2(G233gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(G71gat), .A2(G78gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(G71gat), .A2(G78gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G57gat), .B(G64gat), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G57gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G64gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n399), .A2(G57gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(G71gat), .B(G78gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n648), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT10), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n619), .B2(new_n615), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n609), .A2(new_n611), .A3(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT96), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT96), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n609), .A2(new_n611), .A3(new_n657), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n612), .A2(new_n614), .A3(new_n658), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n659), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n643), .B1(new_n661), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n643), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  INV_X1    g473(.A(G176gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(new_n215), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n677), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n670), .A2(new_n672), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n543), .B1(KEYINPUT21), .B2(new_n657), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(G183gat), .ZN(new_n684));
  AND2_X1   g483(.A1(G231gat), .A2(G233gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n684), .A2(new_n685), .ZN(new_n688));
  XNOR2_X1  g487(.A(G127gat), .B(G155gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(new_n210), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n690), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n684), .A2(new_n685), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n693), .B2(new_n686), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n657), .A2(KEYINPUT21), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n691), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n690), .B1(new_n687), .B2(new_n688), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n693), .A2(new_n686), .A3(new_n692), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n641), .B(new_n682), .C1(new_n699), .C2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n592), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(new_n462), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT97), .B(G1gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1324gat));
  NOR2_X1   g507(.A1(new_n480), .A2(new_n486), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n592), .A2(new_n710), .A3(new_n704), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT98), .B(G8gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(new_n524), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n711), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n711), .B2(G8gat), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n711), .A2(new_n714), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(G1325gat));
  INV_X1    g518(.A(new_n507), .ZN(new_n720));
  INV_X1    g519(.A(new_n503), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n705), .A2(new_n521), .A3(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n505), .A2(new_n506), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n592), .A2(new_n725), .A3(new_n704), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n521), .B2(new_n726), .ZN(G1326gat));
  NOR2_X1   g526(.A1(new_n705), .A2(new_n281), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT43), .B(G22gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  OAI21_X1  g529(.A(new_n698), .B1(new_n691), .B2(new_n694), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n700), .A2(new_n701), .A3(new_n697), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n589), .A2(KEYINPUT99), .A3(new_n590), .ZN(new_n735));
  AOI21_X1  g534(.A(KEYINPUT99), .B1(new_n589), .B2(new_n590), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n734), .A2(new_n682), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT100), .ZN(new_n740));
  INV_X1    g539(.A(new_n641), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n513), .A2(new_n514), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT44), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n471), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n464), .A2(new_n470), .A3(KEYINPUT101), .A4(new_n467), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n510), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT102), .B1(new_n639), .B2(new_n640), .ZN(new_n750));
  INV_X1    g549(.A(new_n640), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n752), .A3(new_n638), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n748), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n740), .B1(new_n743), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT103), .B1(new_n758), .B2(new_n462), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n760), .A3(new_n499), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n759), .A2(G29gat), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n589), .A2(new_n590), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n733), .A2(new_n763), .A3(new_n681), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n515), .A2(new_n741), .A3(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n552), .A3(new_n499), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT45), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n762), .A2(new_n767), .ZN(G1328gat));
  AOI21_X1  g567(.A(new_n553), .B1(new_n757), .B2(new_n710), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n515), .A2(new_n553), .A3(new_n741), .A4(new_n764), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT46), .B1(new_n772), .B2(new_n709), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n765), .A2(new_n774), .A3(new_n553), .A4(new_n710), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n770), .A2(new_n771), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n773), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT104), .B1(new_n777), .B2(new_n769), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1329gat));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n723), .B(new_n740), .C1(new_n743), .C2(new_n756), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n548), .A2(new_n549), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n725), .A3(new_n782), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT47), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OAI221_X1 g586(.A(new_n784), .B1(new_n780), .B2(KEYINPUT47), .C1(new_n781), .C2(new_n782), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1330gat));
  AOI21_X1  g588(.A(new_n544), .B1(new_n757), .B2(new_n508), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n281), .A2(G50gat), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT106), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n765), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT48), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n790), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n790), .B2(new_n793), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1331gat));
  AOI21_X1  g596(.A(new_n741), .B1(new_n731), .B2(new_n732), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n798), .A2(new_n681), .A3(new_n737), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT107), .ZN(new_n800));
  INV_X1    g599(.A(new_n510), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n745), .B2(new_n746), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n499), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g604(.A1(new_n800), .A2(new_n802), .A3(new_n709), .ZN(new_n806));
  NOR2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  AND2_X1   g606(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n806), .B2(new_n807), .ZN(G1333gat));
  NAND2_X1  g609(.A1(new_n803), .A2(new_n725), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT108), .ZN(new_n812));
  INV_X1    g611(.A(G71gat), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n803), .A2(new_n814), .A3(new_n725), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n803), .A2(G71gat), .A3(new_n722), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT50), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1334gat));
  NAND2_X1  g621(.A1(new_n803), .A2(new_n508), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g623(.A1(new_n733), .A2(new_n738), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n741), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n829), .B1(new_n802), .B2(new_n826), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n682), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(G85gat), .B1(new_n831), .B2(new_n499), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT44), .B1(new_n747), .B2(new_n510), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n755), .A2(new_n833), .B1(new_n742), .B2(KEYINPUT44), .ZN(new_n834));
  INV_X1    g633(.A(new_n825), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n682), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n462), .A2(new_n602), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(G1336gat));
  NAND2_X1  g637(.A1(new_n743), .A2(new_n756), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(new_n710), .A3(new_n681), .A4(new_n825), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G92gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n828), .A2(new_n830), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n709), .A2(G92gat), .A3(new_n682), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT52), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n843), .A2(KEYINPUT109), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n843), .A2(KEYINPUT109), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n847), .B(new_n848), .C1(new_n828), .C2(new_n830), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n840), .B2(G92gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n845), .B1(new_n846), .B2(new_n850), .ZN(G1337gat));
  AOI21_X1  g650(.A(G99gat), .B1(new_n831), .B2(new_n725), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n836), .A2(G99gat), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n722), .ZN(G1338gat));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n855));
  INV_X1    g654(.A(G106gat), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n281), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  NOR4_X1   g657(.A1(new_n834), .A2(new_n682), .A3(new_n835), .A4(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(G106gat), .B1(new_n831), .B2(new_n508), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n855), .B(KEYINPUT53), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n508), .A3(new_n681), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n856), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n855), .A2(KEYINPUT53), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n855), .A2(KEYINPUT53), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n839), .A2(new_n681), .A3(new_n825), .A4(new_n857), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n861), .A2(new_n867), .ZN(G1339gat));
  INV_X1    g667(.A(G113gat), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n661), .A2(new_n668), .A3(new_n643), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT54), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n669), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n661), .A2(new_n668), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n642), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n677), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n870), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n679), .B1(new_n669), .B2(new_n875), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n879), .B(KEYINPUT55), .C1(new_n669), .C2(new_n872), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n680), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT111), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n878), .A2(KEYINPUT111), .A3(new_n880), .A4(new_n680), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n883), .B(new_n884), .C1(new_n736), .C2(new_n735), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n578), .A2(new_n579), .A3(new_n577), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n572), .B1(new_n562), .B2(new_n571), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n586), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n590), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n681), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n755), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n750), .A2(new_n753), .A3(new_n889), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n883), .A2(new_n884), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n734), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n798), .A2(new_n682), .A3(new_n737), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n462), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n466), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n897), .A2(new_n709), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n869), .B1(new_n899), .B2(new_n591), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT112), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n869), .A3(new_n738), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1340gat));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n681), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g704(.A1(new_n899), .A2(new_n733), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g706(.A1(new_n899), .A2(new_n741), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n908), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n909));
  XOR2_X1   g708(.A(KEYINPUT56), .B(G134gat), .Z(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n908), .B2(new_n910), .ZN(G1343gat));
  NAND2_X1  g710(.A1(new_n709), .A2(new_n499), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n722), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n890), .B1(new_n763), .B2(new_n881), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT113), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT113), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n890), .B(new_n916), .C1(new_n763), .C2(new_n881), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n741), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n734), .B1(new_n918), .B2(new_n894), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n281), .B1(new_n919), .B2(new_n896), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT57), .B(new_n281), .C1(new_n895), .C2(new_n896), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT114), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n913), .ZN(new_n925));
  INV_X1    g724(.A(new_n917), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n591), .A2(new_n680), .A3(new_n880), .A4(new_n878), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n916), .B1(new_n927), .B2(new_n890), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n641), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n894), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n733), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n703), .A2(new_n738), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n508), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n925), .B1(new_n933), .B2(KEYINPUT57), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT114), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n895), .A2(new_n896), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n921), .A3(new_n508), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n924), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n226), .B1(new_n939), .B2(new_n738), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT115), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n723), .B(new_n508), .C1(new_n897), .C2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n890), .B1(new_n893), .B2(new_n737), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n754), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n733), .B1(new_n944), .B2(new_n930), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n941), .B(new_n499), .C1(new_n945), .C2(new_n932), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n709), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n942), .A2(new_n947), .A3(G141gat), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(new_n591), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT58), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT58), .B1(new_n948), .B2(new_n591), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n933), .A2(KEYINPUT57), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n952), .A2(new_n591), .A3(new_n937), .A4(new_n913), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT116), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n934), .A2(KEYINPUT116), .A3(new_n591), .A4(new_n937), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(G141gat), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT117), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n951), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n951), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n950), .B1(new_n959), .B2(new_n960), .ZN(G1344gat));
  NOR2_X1   g760(.A1(new_n942), .A2(new_n947), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(new_n229), .A3(new_n681), .ZN(new_n963));
  AOI211_X1 g762(.A(KEYINPUT59), .B(new_n229), .C1(new_n939), .C2(new_n681), .ZN(new_n964));
  XNOR2_X1  g763(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT119), .ZN(new_n966));
  OR3_X1    g765(.A1(new_n641), .A2(new_n881), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n641), .B2(new_n881), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n889), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n929), .A2(new_n969), .ZN(new_n970));
  OAI22_X1  g769(.A1(new_n970), .A2(new_n733), .B1(new_n591), .B2(new_n703), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT120), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI221_X1 g772(.A(KEYINPUT120), .B1(new_n591), .B2(new_n703), .C1(new_n970), .C2(new_n733), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n973), .A2(new_n921), .A3(new_n974), .A4(new_n508), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n936), .A2(new_n508), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT57), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n975), .A2(new_n681), .A3(new_n977), .A4(new_n913), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n965), .B1(new_n978), .B2(G148gat), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n979), .ZN(G1345gat));
  AOI21_X1  g779(.A(G155gat), .B1(new_n962), .B2(new_n733), .ZN(new_n981));
  INV_X1    g780(.A(new_n939), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n982), .A2(new_n734), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n981), .B1(new_n983), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g783(.A(G162gat), .B1(new_n982), .B2(new_n754), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n962), .A2(new_n233), .A3(new_n741), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1347gat));
  NOR2_X1   g786(.A1(new_n709), .A2(new_n499), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n936), .A2(new_n898), .A3(new_n988), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n989), .A2(G169gat), .A3(new_n737), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT121), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n988), .A2(new_n725), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n993), .A2(KEYINPUT122), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n994), .A2(new_n508), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(KEYINPUT122), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n936), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(new_n591), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n992), .B1(new_n999), .B2(G169gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n991), .B1(new_n1000), .B2(new_n990), .ZN(G1348gat));
  NOR3_X1   g800(.A1(new_n997), .A2(new_n675), .A3(new_n682), .ZN(new_n1002));
  INV_X1    g801(.A(new_n989), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(new_n681), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1002), .B1(new_n675), .B2(new_n1004), .ZN(G1349gat));
  OAI21_X1  g804(.A(G183gat), .B1(new_n997), .B2(new_n734), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n733), .A2(new_n319), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1006), .B1(new_n989), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g808(.A1(new_n1003), .A2(new_n301), .A3(new_n755), .ZN(new_n1010));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n998), .A2(new_n741), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1011), .B1(new_n1012), .B2(G190gat), .ZN(new_n1013));
  AOI211_X1 g812(.A(KEYINPUT61), .B(new_n301), .C1(new_n998), .C2(new_n741), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT123), .ZN(new_n1016));
  XNOR2_X1  g815(.A(new_n1015), .B(new_n1016), .ZN(G1351gat));
  AND2_X1   g816(.A1(new_n975), .A2(new_n977), .ZN(new_n1018));
  INV_X1    g817(.A(new_n988), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n1019), .A2(new_n722), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g820(.A(G197gat), .B1(new_n1021), .B2(new_n763), .ZN(new_n1022));
  NOR3_X1   g821(.A1(new_n976), .A2(new_n722), .A3(new_n1019), .ZN(new_n1023));
  NAND3_X1  g822(.A1(new_n1023), .A2(new_n214), .A3(new_n738), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1022), .A2(new_n1024), .ZN(G1352gat));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1026));
  NAND4_X1  g825(.A1(new_n1018), .A2(new_n1026), .A3(new_n681), .A4(new_n1020), .ZN(new_n1027));
  NAND4_X1  g826(.A1(new_n975), .A2(new_n681), .A3(new_n977), .A4(new_n1020), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1028), .A2(KEYINPUT126), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n1027), .A2(G204gat), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g829(.A1(new_n1023), .A2(new_n215), .A3(new_n681), .ZN(new_n1031));
  INV_X1    g830(.A(KEYINPUT124), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g832(.A1(new_n1023), .A2(KEYINPUT124), .A3(new_n215), .A4(new_n681), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g834(.A(KEYINPUT62), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n1035), .B1(KEYINPUT125), .B2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g836(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n1038));
  NAND3_X1  g837(.A1(new_n1033), .A2(new_n1034), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g838(.A1(new_n1030), .A2(new_n1037), .A3(new_n1039), .ZN(G1353gat));
  NAND3_X1  g839(.A1(new_n1023), .A2(new_n210), .A3(new_n733), .ZN(new_n1041));
  NAND4_X1  g840(.A1(new_n975), .A2(new_n733), .A3(new_n977), .A4(new_n1020), .ZN(new_n1042));
  AND3_X1   g841(.A1(new_n1042), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1043));
  AOI21_X1  g842(.A(KEYINPUT63), .B1(new_n1042), .B2(G211gat), .ZN(new_n1044));
  OAI21_X1  g843(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(G1354gat));
  OAI21_X1  g844(.A(G218gat), .B1(new_n1021), .B2(new_n641), .ZN(new_n1046));
  NAND3_X1  g845(.A1(new_n1023), .A2(new_n211), .A3(new_n755), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1046), .A2(new_n1047), .ZN(G1355gat));
endmodule


