

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n368, n369, n370, n371, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806;

  XNOR2_X1 U377 ( .A(n774), .B(n775), .ZN(n359) );
  AND2_X1 U378 ( .A1(n492), .A2(n730), .ZN(n711) );
  XNOR2_X1 U379 ( .A(n503), .B(n502), .ZN(n721) );
  INV_X1 U380 ( .A(n642), .ZN(n647) );
  INV_X1 U381 ( .A(G953), .ZN(n782) );
  BUF_X1 U382 ( .A(G143), .Z(n355) );
  XNOR2_X1 U383 ( .A(n356), .B(n371), .ZN(n600) );
  NAND2_X1 U384 ( .A1(n678), .A2(G234), .ZN(n356) );
  XNOR2_X2 U385 ( .A(n675), .B(KEYINPUT55), .ZN(n676) );
  XNOR2_X2 U386 ( .A(n764), .B(KEYINPUT59), .ZN(n765) );
  NAND2_X2 U387 ( .A1(n741), .A2(n745), .ZN(n486) );
  XNOR2_X1 U388 ( .A(n434), .B(G469), .ZN(n649) );
  XNOR2_X2 U389 ( .A(n358), .B(KEYINPUT34), .ZN(n526) );
  XNOR2_X2 U390 ( .A(n790), .B(n576), .ZN(n775) );
  AND2_X2 U391 ( .A1(n640), .A2(n522), .ZN(n731) );
  AND2_X1 U392 ( .A1(n357), .A2(n422), .ZN(n362) );
  NAND2_X1 U393 ( .A1(n717), .A2(n427), .ZN(n357) );
  NOR2_X2 U394 ( .A1(n617), .A2(n721), .ZN(n358) );
  NAND2_X2 U395 ( .A1(n666), .A2(n742), .ZN(n385) );
  NOR2_X1 U396 ( .A1(n359), .A2(n777), .ZN(G66) );
  NOR2_X1 U397 ( .A1(n428), .A2(n398), .ZN(n390) );
  NOR2_X1 U398 ( .A1(n647), .A2(n648), .ZN(n485) );
  NOR2_X1 U399 ( .A1(n775), .A2(G902), .ZN(n581) );
  XNOR2_X1 U400 ( .A(n510), .B(n509), .ZN(n402) );
  XNOR2_X1 U401 ( .A(n581), .B(n580), .ZN(n640) );
  XOR2_X1 U402 ( .A(n411), .B(KEYINPUT43), .Z(n360) );
  XNOR2_X1 U403 ( .A(KEYINPUT85), .B(n673), .ZN(n361) );
  XNOR2_X1 U404 ( .A(n510), .B(n509), .ZN(n410) );
  NAND2_X2 U405 ( .A1(n391), .A2(n389), .ZN(n388) );
  AND2_X2 U406 ( .A1(n362), .A2(n392), .ZN(n391) );
  NAND2_X2 U407 ( .A1(n536), .A2(n537), .ZN(n539) );
  AND2_X1 U408 ( .A1(n368), .A2(n363), .ZN(G54) );
  INV_X1 U409 ( .A(n720), .ZN(n386) );
  AND2_X1 U410 ( .A1(n781), .A2(n387), .ZN(n720) );
  AND2_X1 U411 ( .A1(n672), .A2(n361), .ZN(n387) );
  NOR2_X1 U412 ( .A1(n480), .A2(n648), .ZN(n464) );
  INV_X1 U413 ( .A(n511), .ZN(n398) );
  INV_X1 U414 ( .A(n795), .ZN(n678) );
  INV_X1 U415 ( .A(KEYINPUT66), .ZN(n509) );
  INV_X1 U416 ( .A(KEYINPUT8), .ZN(n371) );
  INV_X1 U417 ( .A(KEYINPUT79), .ZN(n399) );
  XNOR2_X1 U418 ( .A(n762), .B(n763), .ZN(n368) );
  NAND2_X1 U419 ( .A1(n390), .A2(n429), .ZN(n389) );
  AND2_X1 U420 ( .A1(n667), .A2(n714), .ZN(n516) );
  AND2_X1 U421 ( .A1(n504), .A2(n499), .ZN(n498) );
  NAND2_X1 U422 ( .A1(n451), .A2(n448), .ZN(n804) );
  BUF_X1 U423 ( .A(n709), .Z(n366) );
  NAND2_X1 U424 ( .A1(n450), .A2(n449), .ZN(n448) );
  AND2_X1 U425 ( .A1(n453), .A2(n452), .ZN(n451) );
  XNOR2_X1 U426 ( .A(n505), .B(KEYINPUT31), .ZN(n709) );
  XNOR2_X1 U427 ( .A(n460), .B(n459), .ZN(n645) );
  NOR2_X1 U428 ( .A1(n487), .A2(n730), .ZN(n376) );
  AND2_X1 U429 ( .A1(n471), .A2(n730), .ZN(n736) );
  AND2_X1 U430 ( .A1(n512), .A2(n416), .ZN(n436) );
  XNOR2_X1 U431 ( .A(n439), .B(n683), .ZN(n685) );
  NOR2_X1 U432 ( .A1(n759), .A2(G902), .ZN(n434) );
  INV_X1 U433 ( .A(n640), .ZN(n726) );
  XNOR2_X1 U434 ( .A(n393), .B(n587), .ZN(n430) );
  INV_X1 U435 ( .A(n777), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n523), .B(n560), .ZN(n393) );
  XNOR2_X1 U437 ( .A(n543), .B(n540), .ZN(n395) );
  XNOR2_X1 U438 ( .A(n496), .B(n532), .ZN(n560) );
  INV_X1 U439 ( .A(n397), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n533), .B(n607), .ZN(n523) );
  XNOR2_X1 U441 ( .A(n610), .B(KEYINPUT81), .ZN(n418) );
  XNOR2_X1 U442 ( .A(n497), .B(G119), .ZN(n496) );
  XNOR2_X1 U443 ( .A(n558), .B(G146), .ZN(n397) );
  XNOR2_X1 U444 ( .A(n531), .B(n530), .ZN(n587) );
  XNOR2_X1 U445 ( .A(G116), .B(G122), .ZN(n607) );
  XNOR2_X2 U446 ( .A(G953), .B(KEYINPUT64), .ZN(n795) );
  XOR2_X1 U447 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n533) );
  XOR2_X1 U448 ( .A(KEYINPUT71), .B(G101), .Z(n558) );
  INV_X1 U449 ( .A(G128), .ZN(n535) );
  INV_X1 U450 ( .A(G113), .ZN(n497) );
  INV_X2 U451 ( .A(G143), .ZN(n534) );
  INV_X1 U452 ( .A(KEYINPUT110), .ZN(n459) );
  XNOR2_X1 U453 ( .A(KEYINPUT3), .B(KEYINPUT75), .ZN(n532) );
  NOR2_X2 U454 ( .A1(n611), .A2(n613), .ZN(n745) );
  NOR2_X1 U455 ( .A1(n364), .A2(n709), .ZN(n618) );
  NOR2_X1 U456 ( .A1(n407), .A2(n506), .ZN(n364) );
  NAND2_X1 U457 ( .A1(n365), .A2(n498), .ZN(n369) );
  NAND2_X1 U458 ( .A1(n481), .A2(KEYINPUT44), .ZN(n365) );
  NAND2_X1 U459 ( .A1(n400), .A2(n736), .ZN(n505) );
  XNOR2_X2 U460 ( .A(n375), .B(n554), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n369), .B(KEYINPUT91), .ZN(n627) );
  NAND2_X1 U462 ( .A1(n370), .A2(n379), .ZN(n515) );
  NAND2_X1 U463 ( .A1(n381), .A2(n382), .ZN(n370) );
  NAND2_X1 U464 ( .A1(n600), .A2(G221), .ZN(n574) );
  NAND2_X1 U465 ( .A1(n373), .A2(G137), .ZN(n444) );
  INV_X1 U466 ( .A(n442), .ZN(n373) );
  XNOR2_X2 U467 ( .A(n442), .B(n374), .ZN(n396) );
  XNOR2_X2 U468 ( .A(n489), .B(KEYINPUT4), .ZN(n442) );
  NAND2_X1 U469 ( .A1(n650), .A2(n553), .ZN(n375) );
  NAND2_X1 U470 ( .A1(n431), .A2(n638), .ZN(n377) );
  AND2_X1 U471 ( .A1(n431), .A2(n376), .ZN(n690) );
  NOR2_X1 U472 ( .A1(n377), .A2(n642), .ZN(n620) );
  NAND2_X1 U473 ( .A1(n378), .A2(n463), .ZN(n382) );
  NOR2_X1 U474 ( .A1(n711), .A2(n518), .ZN(n378) );
  INV_X1 U475 ( .A(n380), .ZN(n381) );
  NAND2_X1 U476 ( .A1(n470), .A2(n415), .ZN(n380) );
  NAND2_X1 U477 ( .A1(n380), .A2(KEYINPUT48), .ZN(n379) );
  NAND2_X1 U478 ( .A1(n383), .A2(G210), .ZN(n677) );
  NAND2_X1 U479 ( .A1(n383), .A2(G475), .ZN(n766) );
  XNOR2_X2 U480 ( .A(n510), .B(n509), .ZN(n383) );
  XNOR2_X1 U481 ( .A(n791), .B(n437), .ZN(n684) );
  XNOR2_X2 U482 ( .A(n557), .B(n556), .ZN(n791) );
  XNOR2_X2 U483 ( .A(n384), .B(G472), .ZN(n616) );
  NOR2_X2 U484 ( .A1(n684), .A2(G902), .ZN(n384) );
  XNOR2_X2 U485 ( .A(n385), .B(KEYINPUT19), .ZN(n650) );
  XNOR2_X2 U486 ( .A(n546), .B(n545), .ZN(n666) );
  NAND2_X2 U487 ( .A1(n388), .A2(n386), .ZN(n510) );
  NAND2_X1 U488 ( .A1(n428), .A2(n427), .ZN(n392) );
  XNOR2_X2 U489 ( .A(n394), .B(n430), .ZN(n674) );
  XNOR2_X2 U490 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X2 U491 ( .A(n716), .B(n399), .ZN(n428) );
  BUF_X1 U492 ( .A(n674), .Z(n401) );
  NOR2_X1 U493 ( .A1(n407), .A2(n506), .ZN(n403) );
  BUF_X1 U494 ( .A(n526), .Z(n404) );
  NAND2_X1 U495 ( .A1(n404), .A2(n644), .ZN(n405) );
  NAND2_X1 U496 ( .A1(n526), .A2(n644), .ZN(n500) );
  BUF_X1 U497 ( .A(n650), .Z(n406) );
  XNOR2_X1 U498 ( .A(n400), .B(KEYINPUT99), .ZN(n407) );
  INV_X1 U499 ( .A(n781), .ZN(n408) );
  BUF_X1 U500 ( .A(n400), .Z(n409) );
  XNOR2_X1 U501 ( .A(n400), .B(KEYINPUT99), .ZN(n617) );
  NOR2_X1 U502 ( .A1(G953), .A2(G237), .ZN(n588) );
  INV_X1 U503 ( .A(G137), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n525), .B(n524), .ZN(n625) );
  XNOR2_X1 U505 ( .A(KEYINPUT44), .B(KEYINPUT92), .ZN(n524) );
  OR2_X1 U506 ( .A1(G237), .A2(G902), .ZN(n547) );
  NAND2_X1 U507 ( .A1(G214), .A2(n547), .ZN(n742) );
  XOR2_X1 U508 ( .A(G116), .B(KEYINPUT5), .Z(n562) );
  XOR2_X1 U509 ( .A(G140), .B(KEYINPUT80), .Z(n585) );
  XNOR2_X1 U510 ( .A(G125), .B(G140), .ZN(n565) );
  XOR2_X1 U511 ( .A(KEYINPUT10), .B(KEYINPUT72), .Z(n566) );
  NAND2_X1 U512 ( .A1(n456), .A2(n454), .ZN(n462) );
  NAND2_X1 U513 ( .A1(n455), .A2(n469), .ZN(n454) );
  AND2_X1 U514 ( .A1(n457), .A2(n467), .ZN(n456) );
  INV_X1 U515 ( .A(KEYINPUT1), .ZN(n527) );
  INV_X1 U516 ( .A(n731), .ZN(n472) );
  XNOR2_X1 U517 ( .A(n564), .B(KEYINPUT104), .ZN(n528) );
  INV_X1 U518 ( .A(KEYINPUT46), .ZN(n482) );
  AND2_X1 U519 ( .A1(n646), .A2(n479), .ZN(n477) );
  NOR2_X1 U520 ( .A1(n474), .A2(n473), .ZN(n478) );
  AND2_X1 U521 ( .A1(n645), .A2(n412), .ZN(n473) );
  INV_X1 U522 ( .A(n690), .ZN(n499) );
  NOR2_X1 U523 ( .A1(n423), .A2(n421), .ZN(n422) );
  NOR2_X1 U524 ( .A1(n425), .A2(n669), .ZN(n423) );
  INV_X1 U525 ( .A(n671), .ZN(n426) );
  XOR2_X1 U526 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n590) );
  XOR2_X1 U527 ( .A(G122), .B(G104), .Z(n592) );
  XOR2_X1 U528 ( .A(G902), .B(KEYINPUT15), .Z(n544) );
  XOR2_X1 U529 ( .A(G125), .B(KEYINPUT18), .Z(n542) );
  XNOR2_X1 U530 ( .A(KEYINPUT17), .B(KEYINPUT94), .ZN(n541) );
  INV_X1 U531 ( .A(KEYINPUT45), .ZN(n628) );
  INV_X1 U532 ( .A(KEYINPUT112), .ZN(n662) );
  AND2_X1 U533 ( .A1(n745), .A2(n522), .ZN(n521) );
  XNOR2_X1 U534 ( .A(n529), .B(n559), .ZN(n437) );
  XNOR2_X1 U535 ( .A(G128), .B(KEYINPUT100), .ZN(n569) );
  XNOR2_X1 U536 ( .A(G119), .B(G137), .ZN(n567) );
  XNOR2_X1 U537 ( .A(n488), .B(n603), .ZN(n604) );
  XNOR2_X1 U538 ( .A(G107), .B(KEYINPUT9), .ZN(n601) );
  XNOR2_X1 U539 ( .A(n413), .B(n559), .ZN(n435) );
  XNOR2_X1 U540 ( .A(n485), .B(KEYINPUT28), .ZN(n484) );
  INV_X1 U541 ( .A(KEYINPUT33), .ZN(n502) );
  NOR2_X1 U542 ( .A1(n647), .A2(n472), .ZN(n471) );
  XNOR2_X1 U543 ( .A(n579), .B(KEYINPUT25), .ZN(n580) );
  XOR2_X1 U544 ( .A(KEYINPUT95), .B(n679), .Z(n777) );
  NAND2_X1 U545 ( .A1(n360), .A2(n491), .ZN(n667) );
  XNOR2_X1 U546 ( .A(n432), .B(KEYINPUT32), .ZN(n803) );
  XNOR2_X1 U547 ( .A(n622), .B(KEYINPUT82), .ZN(n433) );
  INV_X1 U548 ( .A(KEYINPUT106), .ZN(n466) );
  NAND2_X1 U549 ( .A1(n731), .A2(n507), .ZN(n506) );
  AND2_X1 U550 ( .A1(n493), .A2(n638), .ZN(n411) );
  AND2_X1 U551 ( .A1(n644), .A2(KEYINPUT86), .ZN(n412) );
  INV_X1 U552 ( .A(n725), .ZN(n522) );
  XOR2_X1 U553 ( .A(n587), .B(n586), .Z(n413) );
  AND2_X1 U554 ( .A1(n641), .A2(n640), .ZN(n414) );
  NAND2_X1 U555 ( .A1(n703), .A2(n656), .ZN(n415) );
  AND2_X1 U556 ( .A1(n508), .A2(n414), .ZN(n416) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT111), .Z(n417) );
  XOR2_X1 U558 ( .A(KEYINPUT22), .B(n612), .Z(n419) );
  XOR2_X1 U559 ( .A(n405), .B(n418), .Z(n420) );
  INV_X1 U560 ( .A(n742), .ZN(n494) );
  AND2_X1 U561 ( .A1(n671), .A2(KEYINPUT67), .ZN(n427) );
  AND2_X1 U562 ( .A1(n426), .A2(n511), .ZN(n421) );
  INV_X1 U563 ( .A(KEYINPUT108), .ZN(n490) );
  INV_X1 U564 ( .A(KEYINPUT67), .ZN(n511) );
  NOR2_X1 U565 ( .A1(n717), .A2(n577), .ZN(n429) );
  INV_X1 U566 ( .A(n427), .ZN(n425) );
  XNOR2_X1 U567 ( .A(n430), .B(G101), .ZN(n778) );
  NAND2_X1 U568 ( .A1(n433), .A2(n431), .ZN(n432) );
  XNOR2_X2 U569 ( .A(n520), .B(n419), .ZN(n431) );
  NAND2_X1 U570 ( .A1(n697), .A2(n803), .ZN(n525) );
  XNOR2_X1 U571 ( .A(n791), .B(n435), .ZN(n759) );
  NAND2_X1 U572 ( .A1(n436), .A2(n438), .ZN(n660) );
  NAND2_X1 U573 ( .A1(n436), .A2(n461), .ZN(n460) );
  INV_X1 U574 ( .A(n667), .ZN(n715) );
  BUF_X1 U575 ( .A(n743), .Z(n438) );
  XNOR2_X1 U576 ( .A(n657), .B(KEYINPUT38), .ZN(n743) );
  XNOR2_X1 U577 ( .A(G113), .B(n355), .ZN(n591) );
  AND2_X1 U578 ( .A1(n706), .A2(n490), .ZN(n469) );
  OR2_X2 U579 ( .A1(n772), .A2(G902), .ZN(n465) );
  INV_X1 U580 ( .A(n461), .ZN(n491) );
  NAND2_X1 U581 ( .A1(n743), .A2(n742), .ZN(n663) );
  BUF_X1 U582 ( .A(n684), .Z(n439) );
  BUF_X1 U583 ( .A(n791), .Z(n440) );
  BUF_X1 U584 ( .A(n716), .Z(n793) );
  INV_X1 U585 ( .A(n657), .ZN(n461) );
  INV_X1 U586 ( .A(n666), .ZN(n657) );
  BUF_X1 U587 ( .A(n711), .Z(n441) );
  NAND2_X1 U588 ( .A1(n442), .A2(n443), .ZN(n445) );
  NAND2_X1 U589 ( .A1(n445), .A2(n444), .ZN(n557) );
  XNOR2_X1 U590 ( .A(n560), .B(n563), .ZN(n529) );
  XNOR2_X1 U591 ( .A(n616), .B(n528), .ZN(n480) );
  INV_X1 U592 ( .A(n450), .ZN(n446) );
  XNOR2_X1 U593 ( .A(n660), .B(n659), .ZN(n668) );
  XNOR2_X1 U594 ( .A(n405), .B(n418), .ZN(n447) );
  XNOR2_X1 U595 ( .A(n500), .B(n418), .ZN(n481) );
  NOR2_X2 U596 ( .A1(n674), .A2(n669), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n519), .A2(n518), .ZN(n514) );
  NAND2_X1 U598 ( .A1(n458), .A2(KEYINPUT108), .ZN(n457) );
  XNOR2_X1 U599 ( .A(n464), .B(KEYINPUT107), .ZN(n458) );
  INV_X1 U600 ( .A(n730), .ZN(n638) );
  INV_X1 U601 ( .A(n616), .ZN(n642) );
  OR2_X1 U602 ( .A1(n616), .A2(n494), .ZN(n643) );
  NAND2_X1 U603 ( .A1(n806), .A2(n804), .ZN(n483) );
  NOR2_X1 U604 ( .A1(n661), .A2(n417), .ZN(n449) );
  INV_X1 U605 ( .A(n668), .ZN(n450) );
  NAND2_X1 U606 ( .A1(n661), .A2(n417), .ZN(n452) );
  NAND2_X1 U607 ( .A1(n668), .A2(n417), .ZN(n453) );
  INV_X1 U608 ( .A(n458), .ZN(n455) );
  NAND2_X1 U609 ( .A1(n645), .A2(n644), .ZN(n702) );
  NOR2_X1 U610 ( .A1(n462), .A2(n491), .ZN(n637) );
  XNOR2_X1 U611 ( .A(n462), .B(KEYINPUT109), .ZN(n493) );
  OR2_X1 U612 ( .A1(n495), .A2(n711), .ZN(n519) );
  INV_X1 U613 ( .A(n495), .ZN(n463) );
  NAND2_X1 U614 ( .A1(n702), .A2(n477), .ZN(n476) );
  XNOR2_X2 U615 ( .A(n465), .B(G478), .ZN(n613) );
  XNOR2_X2 U616 ( .A(n661), .B(n466), .ZN(n706) );
  NAND2_X1 U617 ( .A1(n501), .A2(n730), .ZN(n503) );
  XNOR2_X2 U618 ( .A(n649), .B(n527), .ZN(n730) );
  NOR2_X1 U619 ( .A1(n468), .A2(n494), .ZN(n467) );
  NOR2_X1 U620 ( .A1(n706), .A2(n490), .ZN(n468) );
  XNOR2_X1 U621 ( .A(n483), .B(n482), .ZN(n470) );
  NAND2_X1 U622 ( .A1(n409), .A2(n521), .ZN(n520) );
  NAND2_X1 U623 ( .A1(n651), .A2(n475), .ZN(n474) );
  OR2_X1 U624 ( .A1(n646), .A2(n479), .ZN(n475) );
  NAND2_X1 U625 ( .A1(n478), .A2(n476), .ZN(n653) );
  INV_X1 U626 ( .A(KEYINPUT86), .ZN(n479) );
  NOR2_X1 U627 ( .A1(n480), .A2(n472), .ZN(n501) );
  NAND2_X1 U628 ( .A1(n480), .A2(n726), .ZN(n621) );
  NAND2_X1 U629 ( .A1(n480), .A2(n640), .ZN(n487) );
  NAND2_X1 U630 ( .A1(n447), .A2(n623), .ZN(n624) );
  XNOR2_X1 U631 ( .A(n420), .B(G122), .ZN(G24) );
  NAND2_X1 U632 ( .A1(n738), .A2(n664), .ZN(n665) );
  AND2_X1 U633 ( .A1(n484), .A2(n508), .ZN(n664) );
  XNOR2_X2 U634 ( .A(n486), .B(KEYINPUT41), .ZN(n738) );
  XNOR2_X2 U635 ( .A(n663), .B(n662), .ZN(n741) );
  INV_X1 U636 ( .A(n489), .ZN(n488) );
  XNOR2_X2 U637 ( .A(n539), .B(n538), .ZN(n489) );
  XNOR2_X2 U638 ( .A(n665), .B(KEYINPUT42), .ZN(n806) );
  NAND2_X2 U639 ( .A1(n517), .A2(n516), .ZN(n716) );
  XNOR2_X1 U640 ( .A(n637), .B(KEYINPUT36), .ZN(n492) );
  XNOR2_X1 U641 ( .A(n653), .B(n652), .ZN(n495) );
  NAND2_X1 U642 ( .A1(n515), .A2(n514), .ZN(n517) );
  XNOR2_X1 U643 ( .A(n605), .B(n606), .ZN(n608) );
  XNOR2_X1 U644 ( .A(n619), .B(KEYINPUT103), .ZN(n504) );
  AND2_X1 U645 ( .A1(n647), .A2(n508), .ZN(n507) );
  INV_X1 U646 ( .A(n649), .ZN(n508) );
  XNOR2_X1 U647 ( .A(n643), .B(n513), .ZN(n512) );
  INV_X1 U648 ( .A(KEYINPUT30), .ZN(n513) );
  AND2_X1 U649 ( .A1(n517), .A2(n667), .ZN(n672) );
  INV_X1 U650 ( .A(KEYINPUT48), .ZN(n518) );
  OR2_X2 U651 ( .A1(n614), .A2(n613), .ZN(n661) );
  INV_X1 U652 ( .A(KEYINPUT87), .ZN(n652) );
  INV_X1 U653 ( .A(n558), .ZN(n559) );
  INV_X1 U654 ( .A(n721), .ZN(n749) );
  INV_X1 U655 ( .A(KEYINPUT0), .ZN(n554) );
  INV_X1 U656 ( .A(KEYINPUT62), .ZN(n683) );
  XNOR2_X1 U657 ( .A(n604), .B(G134), .ZN(n605) );
  XNOR2_X1 U658 ( .A(n686), .B(n685), .ZN(n687) );
  XOR2_X1 U659 ( .A(G104), .B(G107), .Z(n531) );
  XNOR2_X1 U660 ( .A(KEYINPUT97), .B(G110), .ZN(n530) );
  NAND2_X1 U661 ( .A1(n534), .A2(G128), .ZN(n537) );
  NAND2_X1 U662 ( .A1(n535), .A2(G143), .ZN(n536) );
  XNOR2_X2 U663 ( .A(KEYINPUT65), .B(KEYINPUT83), .ZN(n538) );
  NAND2_X1 U664 ( .A1(G224), .A2(n678), .ZN(n540) );
  XNOR2_X1 U665 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U666 ( .A(KEYINPUT96), .B(n544), .Z(n577) );
  INV_X1 U667 ( .A(n577), .ZN(n669) );
  NAND2_X1 U668 ( .A1(G210), .A2(n547), .ZN(n545) );
  NOR2_X1 U669 ( .A1(G898), .A2(n782), .ZN(n779) );
  NAND2_X1 U670 ( .A1(G234), .A2(G237), .ZN(n548) );
  XNOR2_X1 U671 ( .A(n548), .B(KEYINPUT14), .ZN(n549) );
  AND2_X1 U672 ( .A1(G902), .A2(n549), .ZN(n630) );
  NAND2_X1 U673 ( .A1(n779), .A2(n630), .ZN(n552) );
  NAND2_X1 U674 ( .A1(G952), .A2(n549), .ZN(n550) );
  XNOR2_X1 U675 ( .A(KEYINPUT98), .B(n550), .ZN(n755) );
  NOR2_X1 U676 ( .A1(G953), .A2(n755), .ZN(n633) );
  INV_X1 U677 ( .A(n633), .ZN(n551) );
  NAND2_X1 U678 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U679 ( .A(G146), .B(KEYINPUT73), .ZN(n555) );
  XNOR2_X1 U680 ( .A(n555), .B(G131), .ZN(n595) );
  XOR2_X1 U681 ( .A(G134), .B(n595), .Z(n556) );
  NAND2_X1 U682 ( .A1(n588), .A2(G210), .ZN(n561) );
  XNOR2_X1 U683 ( .A(n562), .B(n561), .ZN(n563) );
  INV_X1 U684 ( .A(KEYINPUT6), .ZN(n564) );
  XNOR2_X1 U685 ( .A(n566), .B(n565), .ZN(n790) );
  XOR2_X1 U686 ( .A(G110), .B(G146), .Z(n568) );
  XNOR2_X1 U687 ( .A(n568), .B(n567), .ZN(n572) );
  XOR2_X1 U688 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n570) );
  XNOR2_X1 U689 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U690 ( .A(n572), .B(n571), .Z(n575) );
  XNOR2_X1 U691 ( .A(n575), .B(n574), .ZN(n576) );
  NAND2_X1 U692 ( .A1(G234), .A2(n577), .ZN(n578) );
  XNOR2_X1 U693 ( .A(n578), .B(KEYINPUT20), .ZN(n582) );
  NAND2_X1 U694 ( .A1(G217), .A2(n582), .ZN(n579) );
  NAND2_X1 U695 ( .A1(n582), .A2(G221), .ZN(n583) );
  XNOR2_X1 U696 ( .A(n583), .B(KEYINPUT21), .ZN(n725) );
  NAND2_X1 U697 ( .A1(G227), .A2(n678), .ZN(n584) );
  XNOR2_X1 U698 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U699 ( .A(KEYINPUT13), .B(G475), .ZN(n599) );
  NAND2_X1 U700 ( .A1(G214), .A2(n588), .ZN(n589) );
  XNOR2_X1 U701 ( .A(n590), .B(n589), .ZN(n594) );
  XNOR2_X1 U702 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U703 ( .A(n594), .B(n593), .Z(n597) );
  XNOR2_X1 U704 ( .A(n595), .B(n790), .ZN(n596) );
  XNOR2_X1 U705 ( .A(n597), .B(n596), .ZN(n764) );
  NOR2_X1 U706 ( .A1(G902), .A2(n764), .ZN(n598) );
  XOR2_X1 U707 ( .A(n599), .B(n598), .Z(n614) );
  INV_X1 U708 ( .A(n614), .ZN(n611) );
  NAND2_X1 U709 ( .A1(G217), .A2(n600), .ZN(n606) );
  XOR2_X1 U710 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n602) );
  XNOR2_X1 U711 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U712 ( .A(n608), .B(n607), .ZN(n772) );
  NAND2_X1 U713 ( .A1(n611), .A2(n613), .ZN(n609) );
  XNOR2_X1 U714 ( .A(KEYINPUT105), .B(n609), .ZN(n644) );
  XNOR2_X1 U715 ( .A(KEYINPUT89), .B(KEYINPUT35), .ZN(n610) );
  XOR2_X1 U716 ( .A(KEYINPUT77), .B(KEYINPUT68), .Z(n612) );
  NAND2_X1 U717 ( .A1(n613), .A2(n614), .ZN(n693) );
  NAND2_X1 U718 ( .A1(n693), .A2(n661), .ZN(n615) );
  XNOR2_X1 U719 ( .A(KEYINPUT102), .B(n615), .ZN(n740) );
  XOR2_X1 U720 ( .A(KEYINPUT88), .B(n740), .Z(n655) );
  NOR2_X1 U721 ( .A1(n618), .A2(n655), .ZN(n619) );
  NAND2_X1 U722 ( .A1(n620), .A2(n726), .ZN(n697) );
  NOR2_X1 U723 ( .A1(n638), .A2(n621), .ZN(n622) );
  INV_X1 U724 ( .A(KEYINPUT44), .ZN(n623) );
  NAND2_X1 U725 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U726 ( .A1(n627), .A2(n626), .ZN(n629) );
  XNOR2_X2 U727 ( .A(n629), .B(n628), .ZN(n717) );
  NAND2_X1 U728 ( .A1(n795), .A2(n630), .ZN(n631) );
  NOR2_X1 U729 ( .A1(G900), .A2(n631), .ZN(n632) );
  NOR2_X1 U730 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U731 ( .A(n634), .B(KEYINPUT84), .ZN(n635) );
  NOR2_X1 U732 ( .A1(n725), .A2(n635), .ZN(n641) );
  XNOR2_X1 U733 ( .A(KEYINPUT74), .B(n641), .ZN(n636) );
  NAND2_X1 U734 ( .A1(n636), .A2(n726), .ZN(n648) );
  INV_X1 U735 ( .A(n740), .ZN(n639) );
  NAND2_X1 U736 ( .A1(KEYINPUT47), .A2(n639), .ZN(n646) );
  NAND2_X1 U737 ( .A1(n664), .A2(n406), .ZN(n654) );
  NAND2_X1 U738 ( .A1(KEYINPUT47), .A2(n654), .ZN(n651) );
  INV_X1 U739 ( .A(n654), .ZN(n703) );
  NOR2_X1 U740 ( .A1(KEYINPUT47), .A2(n655), .ZN(n656) );
  XOR2_X1 U741 ( .A(KEYINPUT76), .B(KEYINPUT90), .Z(n658) );
  XNOR2_X1 U742 ( .A(KEYINPUT39), .B(n658), .ZN(n659) );
  OR2_X1 U743 ( .A1(n693), .A2(n446), .ZN(n714) );
  NAND2_X1 U744 ( .A1(KEYINPUT2), .A2(n669), .ZN(n670) );
  XOR2_X1 U745 ( .A(n670), .B(KEYINPUT69), .Z(n671) );
  INV_X1 U746 ( .A(n717), .ZN(n781) );
  NAND2_X1 U747 ( .A1(KEYINPUT2), .A2(n714), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n401), .B(KEYINPUT54), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n677), .B(n676), .ZN(n680) );
  NOR2_X1 U750 ( .A1(n678), .A2(G952), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n680), .A2(n363), .ZN(n682) );
  INV_X1 U752 ( .A(KEYINPUT56), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(G51) );
  NAND2_X1 U754 ( .A1(n410), .A2(G472), .ZN(n686) );
  NAND2_X1 U755 ( .A1(n687), .A2(n363), .ZN(n689) );
  XOR2_X1 U756 ( .A(KEYINPUT63), .B(KEYINPUT93), .Z(n688) );
  XNOR2_X1 U757 ( .A(n689), .B(n688), .ZN(G57) );
  XOR2_X1 U758 ( .A(n690), .B(G101), .Z(G3) );
  XOR2_X1 U759 ( .A(G104), .B(KEYINPUT113), .Z(n692) );
  NAND2_X1 U760 ( .A1(n403), .A2(n706), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n692), .B(n691), .ZN(G6) );
  XOR2_X1 U762 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n695) );
  INV_X1 U763 ( .A(n693), .ZN(n708) );
  NAND2_X1 U764 ( .A1(n403), .A2(n708), .ZN(n694) );
  XNOR2_X1 U765 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U766 ( .A(G107), .B(n696), .ZN(G9) );
  XNOR2_X1 U767 ( .A(G110), .B(KEYINPUT114), .ZN(n698) );
  XNOR2_X1 U768 ( .A(n698), .B(n697), .ZN(G12) );
  XOR2_X1 U769 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n700) );
  NAND2_X1 U770 ( .A1(n708), .A2(n703), .ZN(n699) );
  XNOR2_X1 U771 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U772 ( .A(G128), .B(n701), .Z(G30) );
  XNOR2_X1 U773 ( .A(n355), .B(n702), .ZN(G45) );
  NAND2_X1 U774 ( .A1(n706), .A2(n703), .ZN(n704) );
  XNOR2_X1 U775 ( .A(n704), .B(KEYINPUT116), .ZN(n705) );
  XNOR2_X1 U776 ( .A(G146), .B(n705), .ZN(G48) );
  NAND2_X1 U777 ( .A1(n706), .A2(n366), .ZN(n707) );
  XNOR2_X1 U778 ( .A(n707), .B(G113), .ZN(G15) );
  NAND2_X1 U779 ( .A1(n366), .A2(n708), .ZN(n710) );
  XNOR2_X1 U780 ( .A(n710), .B(G116), .ZN(G18) );
  XOR2_X1 U781 ( .A(KEYINPUT37), .B(KEYINPUT117), .Z(n713) );
  XNOR2_X1 U782 ( .A(n441), .B(G125), .ZN(n712) );
  XNOR2_X1 U783 ( .A(n713), .B(n712), .ZN(G27) );
  XNOR2_X1 U784 ( .A(G134), .B(n714), .ZN(G36) );
  XOR2_X1 U785 ( .A(n715), .B(G140), .Z(G42) );
  NOR2_X1 U786 ( .A1(n793), .A2(n408), .ZN(n718) );
  NOR2_X1 U787 ( .A1(KEYINPUT2), .A2(n718), .ZN(n719) );
  NOR2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n723) );
  AND2_X1 U789 ( .A1(n738), .A2(n749), .ZN(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U791 ( .A1(n724), .A2(n782), .ZN(n757) );
  NAND2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U793 ( .A(KEYINPUT49), .B(n727), .ZN(n728) );
  NOR2_X1 U794 ( .A1(n642), .A2(n728), .ZN(n729) );
  XOR2_X1 U795 ( .A(KEYINPUT118), .B(n729), .Z(n734) );
  NOR2_X1 U796 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U797 ( .A(KEYINPUT50), .B(n732), .ZN(n733) );
  NOR2_X1 U798 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U799 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U800 ( .A(n737), .B(KEYINPUT51), .ZN(n739) );
  NAND2_X1 U801 ( .A1(n739), .A2(n738), .ZN(n752) );
  NAND2_X1 U802 ( .A1(n741), .A2(n740), .ZN(n748) );
  NOR2_X1 U803 ( .A1(n438), .A2(n742), .ZN(n744) );
  XNOR2_X1 U804 ( .A(KEYINPUT119), .B(n744), .ZN(n746) );
  NAND2_X1 U805 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U806 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U807 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U808 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U809 ( .A(KEYINPUT52), .B(n753), .Z(n754) );
  NOR2_X1 U810 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U811 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U812 ( .A(n758), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U813 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n761) );
  XNOR2_X1 U814 ( .A(n759), .B(KEYINPUT57), .ZN(n760) );
  XNOR2_X1 U815 ( .A(n761), .B(n760), .ZN(n763) );
  NAND2_X1 U816 ( .A1(G469), .A2(n402), .ZN(n762) );
  XNOR2_X1 U817 ( .A(n766), .B(n765), .ZN(n767) );
  NAND2_X1 U818 ( .A1(n767), .A2(n363), .ZN(n770) );
  XNOR2_X1 U819 ( .A(KEYINPUT60), .B(KEYINPUT70), .ZN(n768) );
  XNOR2_X1 U820 ( .A(n768), .B(KEYINPUT121), .ZN(n769) );
  XNOR2_X1 U821 ( .A(n770), .B(n769), .ZN(G60) );
  NAND2_X1 U822 ( .A1(G478), .A2(n402), .ZN(n771) );
  XNOR2_X1 U823 ( .A(n772), .B(n771), .ZN(n773) );
  NOR2_X1 U824 ( .A1(n773), .A2(n777), .ZN(G63) );
  NAND2_X1 U825 ( .A1(G217), .A2(n402), .ZN(n774) );
  XNOR2_X1 U826 ( .A(n778), .B(KEYINPUT123), .ZN(n780) );
  NOR2_X1 U827 ( .A1(n780), .A2(n779), .ZN(n789) );
  NAND2_X1 U828 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U829 ( .A1(G953), .A2(G224), .ZN(n783) );
  XNOR2_X1 U830 ( .A(KEYINPUT61), .B(n783), .ZN(n784) );
  NAND2_X1 U831 ( .A1(n784), .A2(G898), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U833 ( .A(n787), .B(KEYINPUT122), .ZN(n788) );
  XNOR2_X1 U834 ( .A(n789), .B(n788), .ZN(G69) );
  XNOR2_X1 U835 ( .A(n440), .B(n790), .ZN(n792) );
  XNOR2_X1 U836 ( .A(n792), .B(KEYINPUT124), .ZN(n797) );
  XOR2_X1 U837 ( .A(n797), .B(n793), .Z(n794) );
  NOR2_X1 U838 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U839 ( .A(KEYINPUT125), .B(n796), .ZN(n802) );
  XNOR2_X1 U840 ( .A(G227), .B(n797), .ZN(n798) );
  NAND2_X1 U841 ( .A1(n798), .A2(G900), .ZN(n799) );
  NAND2_X1 U842 ( .A1(n799), .A2(G953), .ZN(n800) );
  XNOR2_X1 U843 ( .A(KEYINPUT126), .B(n800), .ZN(n801) );
  NAND2_X1 U844 ( .A1(n802), .A2(n801), .ZN(G72) );
  XNOR2_X1 U845 ( .A(G119), .B(n803), .ZN(G21) );
  XOR2_X1 U846 ( .A(n804), .B(G131), .Z(n805) );
  XNOR2_X1 U847 ( .A(KEYINPUT127), .B(n805), .ZN(G33) );
  XNOR2_X1 U848 ( .A(n806), .B(G137), .ZN(G39) );
endmodule

