//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1313, new_n1314, new_n1315,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n210), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT65), .ZN(new_n221));
  AND2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n220), .A2(new_n221), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n227), .B1(new_n203), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT64), .B(G77), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n229), .B1(G244), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n225), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(new_n215), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n212), .B(new_n218), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n248), .B(new_n252), .ZN(G351));
  NAND2_X1  g0053(.A1(new_n213), .A2(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n254), .A2(new_n255), .A3(G50), .A4(new_n209), .ZN(new_n256));
  INV_X1    g0056(.A(G13), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(G50), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n204), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n210), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n210), .A2(G33), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  OAI221_X1 g0066(.A(new_n261), .B1(new_n262), .B2(new_n264), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n255), .A2(new_n209), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n260), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AND2_X1   g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(new_n272), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G226), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(new_n279), .B(KEYINPUT68), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OR2_X1    g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(KEYINPUT69), .A3(G1698), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n282), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(G222), .A3(new_n287), .ZN(new_n294));
  INV_X1    g0094(.A(new_n230), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n291), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n281), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n280), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n269), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(G179), .B2(new_n298), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT70), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n269), .B(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n280), .A2(G190), .A3(new_n297), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n280), .B2(new_n297), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n304), .B(new_n305), .C1(new_n307), .C2(KEYINPUT72), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(KEYINPUT72), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT10), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n304), .A2(new_n305), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n307), .A2(KEYINPUT72), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n309), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n230), .A2(G20), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT15), .B(G87), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n317), .B1(new_n265), .B2(new_n318), .C1(new_n264), .C2(new_n266), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n319), .A2(new_n268), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n255), .A2(new_n209), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n254), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n323), .B1(new_n230), .B2(new_n259), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n228), .B1(new_n288), .B2(new_n292), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n291), .A2(G232), .A3(new_n287), .ZN(new_n327));
  INV_X1    g0127(.A(G107), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n291), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n281), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n281), .A2(new_n270), .A3(new_n274), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n277), .A2(new_n274), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(G244), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n306), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT71), .B1(new_n325), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT71), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n320), .A2(new_n324), .ZN(new_n338));
  AND2_X1   g0138(.A1(new_n330), .A2(new_n334), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n306), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n330), .A2(new_n334), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n336), .B(new_n340), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(new_n299), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n325), .A3(new_n346), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n302), .A2(new_n316), .A3(new_n343), .A4(new_n347), .ZN(new_n348));
  NOR3_X1   g0148(.A1(new_n257), .A2(new_n210), .A3(G1), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n266), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n322), .B2(new_n266), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n289), .A2(new_n210), .A3(new_n290), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n290), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n355), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n355), .A2(KEYINPUT76), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(G68), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G20), .A2(G33), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n359), .B1(new_n360), .B2(G159), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n359), .A3(G159), .ZN(new_n363));
  XNOR2_X1  g0163(.A(G58), .B(G68), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n362), .A2(new_n363), .B1(G20), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT16), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(G20), .ZN(new_n369));
  INV_X1    g0169(.A(new_n363), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n361), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n354), .A2(new_n355), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(G68), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n321), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n351), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n282), .A2(new_n287), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n376), .B1(G226), .B2(new_n287), .C1(new_n284), .C2(new_n285), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n277), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n276), .B1(new_n332), .B2(new_n237), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n299), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(G179), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT18), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n351), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT16), .B1(new_n358), .B2(new_n365), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n286), .B2(new_n210), .ZN(new_n387));
  INV_X1    g0187(.A(new_n355), .ZN(new_n388));
  OAI21_X1  g0188(.A(G68), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(KEYINPUT16), .A3(new_n365), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n268), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n385), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n381), .A2(G179), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n299), .B2(new_n381), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n384), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n331), .B1(G232), .B2(new_n333), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n377), .A2(new_n378), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n281), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n341), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n306), .B1(new_n379), .B2(new_n380), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n403), .B(new_n385), .C1(new_n386), .C2(new_n391), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT17), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n322), .A2(new_n203), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT73), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n360), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n323), .B2(new_n265), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n412), .A2(new_n268), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n349), .A2(new_n203), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n415), .B(KEYINPUT12), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(KEYINPUT11), .ZN(new_n417));
  AND4_X1   g0217(.A1(new_n410), .A2(new_n414), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n291), .A2(G232), .A3(G1698), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G97), .ZN(new_n424));
  OAI211_X1 g0224(.A(G226), .B(new_n287), .C1(new_n284), .C2(new_n285), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n281), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n331), .B1(G238), .B2(new_n333), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n427), .B2(new_n428), .ZN(new_n431));
  OAI211_X1 g0231(.A(G169), .B(new_n422), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n428), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(G179), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n435), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n422), .B1(new_n438), .B2(G169), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n419), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(G200), .B1(new_n430), .B2(new_n431), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(G190), .A3(new_n435), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n418), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n397), .A2(new_n408), .A3(new_n440), .A4(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n348), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(G20), .B1(new_n263), .B2(G97), .ZN(new_n447));
  AND3_X1   g0247(.A1(KEYINPUT77), .A2(G33), .A3(G283), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n255), .A2(new_n209), .B1(G20), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(KEYINPUT20), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT83), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n450), .A2(new_n455), .A3(KEYINPUT20), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n450), .A2(new_n452), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT20), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n259), .A2(new_n451), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n321), .B(new_n259), .C1(G1), .C2(new_n263), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(new_n451), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G303), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n289), .A2(new_n466), .A3(new_n290), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n281), .ZN(new_n468));
  OR2_X1    g0268(.A1(G257), .A2(G1698), .ZN(new_n469));
  INV_X1    g0269(.A(G264), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G1698), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n469), .A2(new_n471), .B1(new_n289), .B2(new_n290), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT82), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n471), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n291), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT82), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n281), .A4(new_n467), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(G1), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(G270), .A3(new_n277), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT81), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n486), .A3(G270), .A4(new_n277), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n273), .A2(new_n480), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n478), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n465), .A2(new_n491), .A3(G169), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT21), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(G200), .ZN(new_n495));
  INV_X1    g0295(.A(new_n465), .ZN(new_n496));
  INV_X1    g0296(.A(new_n490), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n497), .B1(new_n473), .B2(new_n477), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(G190), .A3(new_n488), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(KEYINPUT21), .A2(G169), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n478), .A2(new_n488), .A3(new_n344), .A4(new_n490), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n465), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n494), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n503), .A2(new_n465), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n507), .A2(new_n502), .B1(new_n492), .B2(new_n493), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT84), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n509), .A3(new_n500), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n356), .A2(G107), .A3(new_n357), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n328), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  INV_X1    g0313(.A(G97), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n514), .A2(new_n328), .ZN(new_n515));
  NOR2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n513), .B1(new_n517), .B2(KEYINPUT6), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G20), .B1(G77), .B2(new_n360), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n268), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n259), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n463), .B2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G250), .A2(G1698), .ZN(new_n524));
  NAND2_X1  g0324(.A1(KEYINPUT4), .A2(G244), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G1698), .ZN(new_n526));
  INV_X1    g0326(.A(new_n449), .ZN(new_n527));
  NAND3_X1  g0327(.A1(KEYINPUT77), .A2(G33), .A3(G283), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n291), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G244), .B(new_n287), .C1(new_n284), .C2(new_n285), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n277), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n483), .A2(G257), .A3(new_n277), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n490), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n341), .B1(new_n306), .B2(KEYINPUT78), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(KEYINPUT78), .B(G200), .C1(new_n533), .C2(new_n535), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n521), .A2(new_n523), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n321), .B1(new_n512), .B2(new_n519), .ZN(new_n541));
  INV_X1    g0341(.A(new_n523), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n529), .A2(new_n532), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n281), .ZN(new_n544));
  INV_X1    g0344(.A(new_n535), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n299), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n533), .A2(new_n535), .A3(new_n344), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n541), .A2(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G250), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(G1698), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n284), .B2(new_n285), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT86), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n291), .A2(G257), .A3(G1698), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G294), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT86), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n551), .B(new_n556), .C1(new_n285), .C2(new_n284), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n281), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n281), .B1(new_n480), .B2(new_n489), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G264), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n559), .A2(new_n341), .A3(new_n490), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT87), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n490), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n306), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n558), .A2(new_n281), .B1(G264), .B2(new_n560), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT87), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n341), .A4(new_n490), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n210), .B(G87), .C1(new_n284), .C2(new_n285), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT22), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT22), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n291), .A2(new_n572), .A3(new_n210), .A4(G87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n328), .A2(G20), .ZN(new_n575));
  OAI22_X1  g0375(.A1(KEYINPUT23), .A2(new_n575), .B1(new_n265), .B2(new_n451), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT85), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(KEYINPUT23), .C1(new_n210), .C2(G107), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n577), .B1(new_n575), .B2(KEYINPUT23), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n576), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n574), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n321), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n259), .A2(G107), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT25), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n588), .B1(new_n328), .B2(new_n462), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n569), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n549), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n550), .B1(new_n213), .B2(G45), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n273), .A2(new_n480), .B1(new_n277), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(G238), .A2(G1698), .ZN(new_n595));
  INV_X1    g0395(.A(G244), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(G1698), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n291), .B1(G33), .B2(G116), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n598), .B2(new_n277), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(G179), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n299), .B2(new_n599), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(new_n210), .A3(G33), .A4(G97), .ZN(new_n603));
  INV_X1    g0403(.A(G87), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n516), .A2(new_n604), .B1(new_n424), .B2(new_n210), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n605), .B2(new_n602), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT79), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n291), .A2(new_n607), .A3(new_n210), .A4(G68), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n210), .B(G68), .C1(new_n284), .C2(new_n285), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT79), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n606), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n268), .ZN(new_n612));
  INV_X1    g0412(.A(new_n318), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n463), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n318), .A2(new_n349), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT80), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n611), .A2(new_n268), .B1(new_n349), .B2(new_n318), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT80), .B1(new_n619), .B2(new_n614), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n601), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n564), .A2(new_n299), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n566), .A2(new_n344), .A3(new_n490), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n622), .B(new_n623), .C1(new_n586), .C2(new_n589), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n463), .A2(G87), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n599), .A2(G200), .ZN(new_n627));
  OAI211_X1 g0427(.A(G190), .B(new_n594), .C1(new_n598), .C2(new_n277), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n592), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n446), .A2(new_n511), .A3(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n302), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n316), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n311), .A2(new_n315), .A3(KEYINPUT90), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n408), .A2(new_n444), .ZN(new_n638));
  INV_X1    g0438(.A(new_n347), .ZN(new_n639));
  OAI21_X1  g0439(.A(G169), .B1(new_n430), .B2(new_n431), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n421), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n436), .A3(new_n432), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n419), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n397), .B1(new_n638), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n633), .B1(new_n637), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n446), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n616), .A2(new_n617), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n619), .A2(KEYINPUT80), .A3(new_n614), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n228), .A2(new_n287), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n596), .A2(G1698), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n650), .B(new_n651), .C1(new_n284), .C2(new_n285), .ZN(new_n652));
  NAND2_X1  g0452(.A1(G33), .A2(G116), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n277), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI211_X1 g0456(.A(KEYINPUT88), .B(new_n277), .C1(new_n652), .C2(new_n653), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n594), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n600), .B1(new_n658), .B2(new_n299), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n612), .A2(new_n625), .A3(new_n628), .A4(new_n615), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n661), .B1(G200), .B2(new_n658), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  INV_X1    g0464(.A(new_n548), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n660), .A2(new_n663), .A3(new_n664), .A4(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n621), .A2(new_n629), .A3(new_n665), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n660), .B(new_n666), .C1(new_n667), .C2(new_n664), .ZN(new_n668));
  INV_X1    g0468(.A(new_n624), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n494), .A2(new_n504), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n662), .B1(new_n649), .B2(new_n659), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n549), .A3(new_n591), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n673), .B2(KEYINPUT89), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT89), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n672), .A2(new_n549), .A3(new_n591), .A4(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n668), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n645), .B1(new_n646), .B2(new_n677), .ZN(G369));
  OR2_X1    g0478(.A1(new_n586), .A2(new_n589), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n622), .A2(new_n623), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n258), .A2(new_n210), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n258), .A2(new_n683), .A3(new_n210), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(G213), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT91), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n682), .A2(new_n687), .A3(G213), .A4(new_n684), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(G343), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n679), .B1(new_n680), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n591), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n669), .A2(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n509), .B1(new_n508), .B2(new_n500), .ZN(new_n695));
  AND4_X1   g0495(.A1(new_n509), .A2(new_n494), .A3(new_n500), .A4(new_n504), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT92), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n496), .A2(new_n689), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT92), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n506), .A2(new_n510), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n670), .A2(new_n698), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n706));
  OAI211_X1 g0506(.A(G330), .B(new_n694), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n690), .B1(new_n494), .B2(new_n504), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n691), .A2(new_n591), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n689), .B(KEYINPUT94), .Z(new_n710));
  NAND2_X1  g0510(.A1(new_n669), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n707), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(G41), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n216), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n516), .A2(new_n604), .A3(new_n451), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n715), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n207), .B2(new_n715), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n273), .A2(new_n480), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n277), .A2(new_n593), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n723), .A2(new_n654), .A3(new_n344), .ZN(new_n724));
  AND4_X1   g0524(.A1(new_n488), .A2(new_n566), .A3(new_n498), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT30), .B1(new_n725), .B2(new_n536), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n564), .A2(new_n491), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n544), .A2(new_n545), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n658), .A2(new_n728), .A3(new_n344), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n566), .A2(new_n488), .A3(new_n498), .A4(new_n724), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n536), .A2(KEYINPUT30), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n727), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n689), .B(KEYINPUT94), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT31), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT95), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n726), .B2(new_n732), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n730), .A2(new_n731), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n730), .B2(new_n728), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n536), .A2(G179), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n491), .A3(new_n564), .A4(new_n658), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n739), .A2(new_n741), .A3(KEYINPUT95), .A4(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n738), .A2(new_n690), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n736), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n631), .A2(new_n511), .A3(new_n710), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT96), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(new_n673), .B2(new_n671), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n540), .A2(new_n548), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n590), .B2(new_n569), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n508), .A2(new_n624), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(KEYINPUT96), .A3(new_n672), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n621), .A2(new_n665), .A3(new_n664), .A4(new_n629), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n660), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n664), .B1(new_n672), .B2(new_n665), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n751), .B(new_n690), .C1(new_n758), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n676), .A3(new_n756), .ZN(new_n765));
  INV_X1    g0565(.A(new_n668), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT29), .B1(new_n767), .B2(new_n710), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n750), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n720), .B1(new_n770), .B2(G1), .ZN(G364));
  NAND2_X1  g0571(.A1(new_n702), .A2(new_n704), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(KEYINPUT93), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G330), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(G330), .B1(new_n705), .B2(new_n706), .ZN(new_n779));
  INV_X1    g0579(.A(new_n715), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n257), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n213), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n778), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n210), .B1(KEYINPUT98), .B2(new_n299), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(KEYINPUT98), .B2(new_n299), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n271), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G13), .A2(G33), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT99), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n216), .A2(new_n291), .ZN(new_n797));
  INV_X1    g0597(.A(G355), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n798), .B1(G116), .B2(new_n216), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n252), .A2(G45), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n216), .A2(new_n286), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n479), .B2(new_n208), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n799), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n210), .A2(G179), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n286), .B1(new_n805), .B2(new_n466), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT100), .Z(new_n807));
  NOR2_X1   g0607(.A1(new_n210), .A2(new_n344), .ZN(new_n808));
  NOR2_X1   g0608(.A1(G190), .A2(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n804), .A2(new_n809), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G311), .A2(new_n811), .B1(new_n813), .B2(G329), .ZN(new_n814));
  INV_X1    g0614(.A(G322), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n808), .A2(G190), .A3(new_n306), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n808), .A2(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G190), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(KEYINPUT33), .B(G317), .Z(new_n821));
  NAND3_X1  g0621(.A1(new_n804), .A2(new_n341), .A3(G200), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n818), .A2(new_n341), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G326), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n341), .A2(G179), .A3(G200), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n210), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n826), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n817), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n813), .A2(G159), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT32), .ZN(new_n833));
  INV_X1    g0633(.A(new_n825), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n201), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G68), .B2(new_n819), .ZN(new_n836));
  INV_X1    g0636(.A(new_n805), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G87), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n514), .B2(new_n829), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n832), .A2(KEYINPUT32), .B1(new_n328), .B2(new_n822), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n291), .B1(new_n816), .B2(new_n202), .C1(new_n295), .C2(new_n810), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n807), .A2(new_n831), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n784), .B1(new_n796), .B2(new_n803), .C1(new_n843), .C2(new_n790), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n776), .B2(new_n794), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n787), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G396));
  OAI21_X1  g0647(.A(new_n286), .B1(new_n805), .B2(new_n328), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT101), .ZN(new_n849));
  INV_X1    g0649(.A(G311), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n810), .A2(new_n451), .B1(new_n812), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n816), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(G294), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n829), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G97), .A2(new_n854), .B1(new_n819), .B2(G283), .ZN(new_n855));
  INV_X1    g0655(.A(new_n822), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n825), .A2(G303), .B1(new_n856), .B2(G87), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n849), .A2(new_n853), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n852), .A2(G143), .B1(new_n811), .B2(G159), .ZN(new_n859));
  INV_X1    g0659(.A(G137), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n834), .B2(new_n860), .C1(new_n262), .C2(new_n820), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT102), .Z(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT34), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n856), .A2(G68), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n286), .B1(new_n813), .B2(G132), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n854), .A2(G58), .B1(new_n837), .B2(G50), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n864), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n862), .A2(KEYINPUT34), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n858), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n791), .A2(new_n792), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n869), .A2(new_n791), .B1(new_n323), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n347), .A2(new_n690), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n338), .A2(new_n689), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n343), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n875), .B2(new_n347), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n871), .B1(new_n876), .B2(new_n793), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n784), .ZN(new_n878));
  INV_X1    g0678(.A(new_n872), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n342), .A2(new_n341), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n338), .B1(new_n339), .B2(new_n306), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(KEYINPUT71), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n873), .B1(new_n882), .B2(new_n340), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n879), .B1(new_n883), .B2(new_n639), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n677), .B2(new_n734), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n767), .A2(new_n710), .A3(new_n876), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n750), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n785), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n750), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(G384));
  NOR2_X1   g0694(.A1(new_n781), .A2(new_n213), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT40), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n419), .A2(new_n690), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n440), .A2(new_n444), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n419), .B(new_n690), .C1(new_n642), .C2(new_n443), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n876), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n745), .A2(new_n746), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n690), .A4(new_n744), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n748), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n392), .A2(new_n395), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n686), .A2(new_n688), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n392), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n906), .A2(new_n909), .A3(new_n910), .A4(new_n405), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(new_n909), .A3(new_n405), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n384), .A2(new_n404), .A3(new_n407), .A4(new_n396), .ZN(new_n914));
  INV_X1    g0714(.A(new_n909), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n911), .A2(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT105), .B1(new_n916), .B2(KEYINPUT38), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n911), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT105), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT38), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n390), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n268), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n925), .B2(KEYINPUT104), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(new_n268), .C1(new_n373), .C2(KEYINPUT16), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n351), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n907), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n914), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT16), .B1(new_n389), .B2(new_n365), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT104), .B1(new_n932), .B2(new_n321), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n390), .A3(new_n928), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n385), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n935), .A2(new_n395), .B1(new_n375), .B2(new_n403), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n908), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n910), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n911), .ZN(new_n939));
  OAI211_X1 g0739(.A(KEYINPUT38), .B(new_n931), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n917), .A2(new_n923), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n896), .B1(new_n905), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n405), .B1(new_n929), .B2(new_n383), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT37), .B1(new_n943), .B2(new_n930), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n911), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n945), .B2(new_n931), .ZN(new_n946));
  INV_X1    g0746(.A(new_n940), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n901), .A2(new_n904), .A3(new_n896), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(G330), .B1(new_n942), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n446), .A2(G330), .A3(new_n904), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT106), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n938), .A2(new_n939), .ZN(new_n955));
  INV_X1    g0755(.A(new_n931), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n922), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n940), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n905), .A2(new_n958), .A3(new_n896), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n901), .A2(new_n904), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n944), .A2(new_n911), .B1(new_n914), .B2(new_n930), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT38), .B1(new_n918), .B2(new_n919), .ZN(new_n962));
  AOI22_X1  g0762(.A1(KEYINPUT38), .A2(new_n961), .B1(new_n962), .B2(new_n921), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n963), .B2(new_n917), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(new_n964), .B2(new_n896), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n965), .A2(new_n446), .A3(new_n904), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n953), .A2(KEYINPUT106), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n954), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n886), .A2(new_n879), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n958), .A3(new_n900), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT39), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n941), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n957), .A2(KEYINPUT39), .A3(new_n940), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n642), .A2(new_n419), .A3(new_n689), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n970), .B1(new_n397), .B2(new_n908), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n758), .A2(new_n762), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(KEYINPUT29), .A3(new_n689), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n751), .B1(new_n677), .B2(new_n734), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n978), .A2(new_n979), .A3(new_n446), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n645), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n976), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n895), .B1(new_n968), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n982), .B2(new_n968), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n518), .A2(KEYINPUT35), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n985), .A2(G116), .A3(new_n211), .A4(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT36), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n208), .B1(new_n202), .B2(new_n203), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n989), .A2(new_n295), .B1(G50), .B2(new_n203), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(G1), .A3(new_n257), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n984), .A2(new_n988), .A3(new_n991), .ZN(G367));
  OAI21_X1  g0792(.A(new_n795), .B1(new_n216), .B2(new_n318), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n243), .A2(new_n801), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n784), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n816), .A2(new_n262), .B1(new_n810), .B2(new_n201), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n286), .B(new_n996), .C1(G137), .C2(new_n813), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n837), .A2(G58), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n819), .A2(G159), .B1(new_n856), .B2(new_n230), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G68), .A2(new_n854), .B1(new_n825), .B2(G143), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(G317), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n286), .B1(new_n812), .B2(new_n1002), .C1(new_n823), .C2(new_n810), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n834), .A2(new_n850), .B1(new_n466), .B2(new_n816), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT111), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n829), .A2(new_n328), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n820), .A2(new_n827), .B1(new_n822), .B2(new_n514), .ZN(new_n1007));
  OR4_X1    g0807(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT112), .B1(new_n805), .B2(new_n451), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT46), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1001), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n995), .B1(new_n1012), .B2(new_n791), .ZN(new_n1013));
  OR3_X1    g0813(.A1(new_n660), .A2(new_n626), .A3(new_n689), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n672), .B1(new_n626), .B2(new_n689), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n794), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n709), .B1(new_n694), .B2(new_n708), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n775), .B2(G330), .ZN(new_n1021));
  OAI211_X1 g0821(.A(G330), .B(new_n1020), .C1(new_n705), .C2(new_n706), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n770), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT109), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1020), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n779), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n769), .B1(new_n1027), .B2(new_n1022), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT109), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT44), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT107), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n710), .B2(new_n548), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n665), .A2(KEYINPUT107), .A3(new_n734), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n734), .B1(new_n541), .B2(new_n542), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1033), .A2(new_n1034), .B1(new_n549), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1031), .B1(new_n712), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n709), .A2(new_n711), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1039), .A2(KEYINPUT44), .A3(new_n1036), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT45), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1039), .B2(new_n1036), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n707), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n775), .A2(new_n1048), .A3(G330), .A4(new_n694), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AND4_X1   g0850(.A1(KEYINPUT110), .A2(new_n1025), .A3(new_n1030), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1024), .B2(KEYINPUT109), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT110), .B1(new_n1053), .B2(new_n1030), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n770), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n715), .B(KEYINPUT41), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n783), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1036), .A2(new_n709), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT108), .Z(new_n1060));
  OR2_X1    g0860(.A1(new_n1060), .A2(KEYINPUT42), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n548), .B1(new_n1036), .B2(new_n624), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1060), .A2(KEYINPUT42), .B1(new_n710), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT43), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1017), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1016), .A2(KEYINPUT43), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .A4(new_n1017), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n707), .A2(new_n1036), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1070), .B(new_n1071), .Z(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1019), .B1(new_n1058), .B2(new_n1073), .ZN(G387));
  NAND3_X1  g0874(.A1(new_n692), .A2(new_n693), .A3(new_n794), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n797), .A2(new_n717), .B1(G107), .B2(new_n216), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n240), .A2(new_n479), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n266), .A2(G50), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT50), .ZN(new_n1080));
  AOI211_X1 g0880(.A(G45), .B(new_n716), .C1(G68), .C2(G77), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n801), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1077), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n784), .B1(new_n1083), .B2(new_n796), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n820), .A2(new_n266), .B1(new_n295), .B2(new_n805), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n613), .B2(new_n854), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n286), .B1(new_n852), .B2(G50), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT113), .B(G150), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n813), .A2(new_n1089), .B1(new_n811), .B2(G68), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n825), .A2(G159), .B1(new_n856), .B2(G97), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1086), .A2(new_n1087), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n291), .B1(new_n813), .B2(G326), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n816), .A2(new_n1002), .B1(new_n810), .B2(new_n466), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n819), .A2(G311), .B1(new_n825), .B2(G322), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT48), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n854), .A2(G283), .B1(new_n837), .B2(G294), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT49), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1093), .B1(new_n451), .B2(new_n822), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1092), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT115), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1076), .B(new_n1084), .C1(new_n1109), .C2(new_n791), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT116), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1027), .A2(new_n1022), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1111), .B1(new_n783), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1028), .A2(new_n715), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n770), .B2(new_n1112), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT117), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(G393));
  NAND2_X1  g0921(.A1(new_n1050), .A2(new_n783), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n795), .B1(new_n514), .B2(new_n216), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n247), .A2(new_n801), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n784), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G159), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n834), .A2(new_n262), .B1(new_n1126), .B2(new_n816), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT51), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n837), .A2(G68), .B1(new_n813), .B2(G143), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT118), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n829), .A2(new_n323), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n291), .B1(new_n810), .B2(new_n266), .C1(new_n604), .C2(new_n822), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(G50), .C2(new_n819), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1128), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT119), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G317), .A2(new_n825), .B1(new_n852), .B2(G311), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT52), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n286), .B1(new_n812), .B2(new_n815), .C1(new_n827), .C2(new_n810), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n820), .A2(new_n466), .B1(new_n822), .B2(new_n328), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n829), .A2(new_n451), .B1(new_n805), .B2(new_n823), .ZN(new_n1141));
  OR4_X1    g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1125), .B1(new_n1144), .B2(new_n791), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n794), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n1037), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1122), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT110), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1050), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n1024), .A2(KEYINPUT109), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1053), .A2(KEYINPUT110), .A3(new_n1030), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n715), .B1(new_n1024), .B2(new_n1052), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(G390));
  OAI211_X1 g0957(.A(G330), .B(new_n879), .C1(new_n883), .C2(new_n639), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n904), .A2(new_n900), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n677), .A2(new_n734), .A3(new_n884), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n900), .B1(new_n1162), .B2(new_n872), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n975), .B1(new_n972), .B2(new_n973), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n941), .A2(new_n975), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n690), .B1(new_n758), .B2(new_n762), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n875), .A2(new_n347), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n879), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1165), .B1(new_n1169), .B2(new_n900), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1161), .B1(new_n1164), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n872), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n900), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n975), .B(new_n941), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n749), .A2(new_n900), .A3(new_n1159), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n972), .A2(new_n973), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n975), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n969), .B2(new_n900), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1174), .B(new_n1176), .C1(new_n1177), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1171), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n980), .A2(new_n645), .A3(new_n952), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1158), .B1(new_n747), .B2(new_n748), .ZN(new_n1183));
  OAI21_X1  g0983(.A(KEYINPUT120), .B1(new_n1183), .B2(new_n900), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1160), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1183), .A2(KEYINPUT120), .A3(new_n900), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n969), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n900), .B1(new_n904), .B2(new_n1159), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1175), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1172), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1182), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1181), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1171), .A2(new_n1191), .A3(new_n1180), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n780), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1171), .A2(new_n783), .A3(new_n1180), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n820), .A2(new_n328), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1131), .B(new_n1197), .C1(G283), .C2(new_n825), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n810), .A2(new_n514), .B1(new_n812), .B2(new_n827), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n291), .B(new_n1199), .C1(G116), .C2(new_n852), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1198), .A2(new_n838), .A3(new_n864), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(G132), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT54), .B(G143), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n816), .A2(new_n1202), .B1(new_n810), .B2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n286), .B(new_n1204), .C1(G125), .C2(new_n813), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1088), .A2(new_n805), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT53), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n819), .A2(G137), .B1(new_n856), .B2(G50), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n829), .A2(new_n1126), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G128), .B2(new_n825), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1205), .A2(new_n1207), .A3(new_n1208), .A4(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n790), .B1(new_n1201), .B2(new_n1211), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n785), .B(new_n1212), .C1(new_n266), .C2(new_n870), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n1177), .B2(new_n793), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1195), .A2(new_n1196), .A3(new_n1214), .ZN(G378));
  XOR2_X1   g1015(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n907), .A2(new_n269), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT55), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n637), .B2(new_n301), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n311), .A2(new_n315), .A3(KEYINPUT90), .ZN(new_n1221));
  AOI21_X1  g1021(.A(KEYINPUT90), .B1(new_n311), .B2(new_n315), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n301), .B(new_n1219), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1217), .B1(new_n1220), .B2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n301), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1219), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1228), .A2(new_n1216), .A3(new_n1223), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n965), .B2(G330), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(G330), .C1(new_n942), .C2(new_n950), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n976), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n974), .A2(new_n975), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n1163), .A2(new_n948), .B1(new_n397), .B2(new_n908), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n951), .A2(new_n1229), .A3(new_n1225), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1232), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1234), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1225), .A2(new_n792), .A3(new_n1229), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n820), .A2(new_n514), .B1(new_n822), .B2(new_n202), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G116), .B2(new_n825), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n286), .A2(new_n714), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G283), .B2(new_n813), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n852), .A2(G107), .B1(new_n811), .B2(new_n613), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n854), .A2(G68), .B1(new_n837), .B2(new_n230), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1243), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1244), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1251));
  AND2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n825), .A2(G125), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n820), .B2(new_n1202), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n852), .A2(G128), .B1(new_n811), .B2(G137), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n805), .B2(new_n1203), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G150), .C2(new_n854), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT59), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n856), .A2(G159), .ZN(new_n1260));
  AOI211_X1 g1060(.A(G33), .B(G41), .C1(new_n813), .C2(G124), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1258), .A2(KEYINPUT59), .ZN(new_n1263));
  OAI221_X1 g1063(.A(new_n1252), .B1(new_n1249), .B2(new_n1248), .C1(new_n1262), .C2(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1264), .A2(new_n791), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n785), .B(new_n1265), .C1(new_n201), .C2(new_n870), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1240), .A2(new_n783), .B1(new_n1241), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1182), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1194), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1240), .A2(new_n1269), .A3(KEYINPUT57), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n780), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1269), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1267), .B1(new_n1271), .B2(new_n1272), .ZN(G375));
  NAND3_X1  g1073(.A1(new_n1187), .A2(new_n1182), .A3(new_n1190), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(KEYINPUT123), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n749), .A2(new_n1159), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT120), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1173), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(new_n1160), .A3(new_n1184), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1279), .A2(new_n969), .B1(new_n1189), .B2(new_n1172), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT123), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1280), .A2(new_n1281), .A3(new_n1182), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1275), .A2(new_n1282), .A3(new_n1192), .A4(new_n1057), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1173), .A2(new_n792), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n834), .A2(new_n827), .B1(new_n822), .B2(new_n323), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(G97), .B2(new_n837), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n816), .A2(new_n823), .B1(new_n812), .B2(new_n466), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n291), .B(new_n1287), .C1(G107), .C2(new_n811), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n613), .A2(new_n854), .B1(new_n819), .B2(G116), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n829), .A2(new_n201), .B1(new_n805), .B2(new_n1126), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1291), .B1(G132), .B2(new_n825), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n286), .B1(new_n813), .B2(G128), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n852), .A2(G137), .B1(new_n811), .B2(G150), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1203), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n819), .A2(new_n1295), .B1(new_n856), .B2(G58), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n790), .B1(new_n1290), .B2(new_n1297), .ZN(new_n1298));
  AOI211_X1 g1098(.A(new_n785), .B(new_n1298), .C1(new_n203), .C2(new_n870), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1284), .A2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1280), .B2(new_n782), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1283), .A2(new_n1302), .ZN(G381));
  INV_X1    g1103(.A(new_n1119), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n846), .A3(new_n1117), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1305), .A2(G384), .ZN(new_n1306));
  XOR2_X1   g1106(.A(new_n1306), .B(KEYINPUT124), .Z(new_n1307));
  AOI22_X1  g1107(.A1(new_n1239), .A2(new_n1234), .B1(new_n1194), .B2(new_n1268), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1270), .B(new_n780), .C1(KEYINPUT57), .C2(new_n1308), .ZN(new_n1309));
  NOR3_X1   g1109(.A1(G390), .A2(G378), .A3(G381), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1307), .A2(new_n1309), .A3(new_n1267), .A4(new_n1310), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1311), .A2(G387), .ZN(G407));
  INV_X1    g1112(.A(G378), .ZN(new_n1313));
  INV_X1    g1113(.A(G343), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  OAI221_X1 g1115(.A(G213), .B1(G375), .B2(new_n1315), .C1(new_n1311), .C2(G387), .ZN(G409));
  XOR2_X1   g1116(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1317));
  INV_X1    g1117(.A(KEYINPUT125), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n893), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT125), .B1(new_n891), .B2(new_n892), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT60), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1275), .B(new_n1282), .C1(new_n1323), .C2(new_n1191), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1274), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n715), .B1(new_n1325), .B2(KEYINPUT60), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1324), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1320), .B(new_n1322), .C1(new_n1327), .C2(new_n1301), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1301), .B1(new_n1324), .B2(new_n1326), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(new_n1318), .A3(new_n893), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1314), .A2(G213), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(G2897), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1328), .A2(new_n1330), .A3(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1333), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1309), .A2(G378), .A3(new_n1267), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1308), .A2(new_n1057), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1267), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1313), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1332), .B1(new_n1337), .B2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1317), .B1(new_n1336), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1341), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1343), .B1(new_n1341), .B2(new_n1344), .ZN(new_n1346));
  NOR3_X1   g1146(.A1(new_n1342), .A2(new_n1345), .A3(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(G396), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1305), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n769), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n782), .B1(new_n1350), .B2(new_n1056), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1072), .ZN(new_n1352));
  AOI21_X1  g1152(.A(G390), .B1(new_n1352), .B2(new_n1019), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1019), .ZN(new_n1354));
  AOI211_X1 g1154(.A(new_n1354), .B(new_n1156), .C1(new_n1351), .C2(new_n1072), .ZN(new_n1355));
  OAI21_X1  g1155(.A(new_n1349), .B1(new_n1353), .B2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G387), .A2(new_n1156), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1349), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1352), .A2(new_n1019), .A3(G390), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1357), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1356), .A2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  AND2_X1   g1162(.A1(new_n1337), .A2(new_n1340), .ZN(new_n1363));
  OAI22_X1  g1163(.A1(new_n1363), .A2(new_n1332), .B1(new_n1335), .B2(new_n1334), .ZN(new_n1364));
  AOI22_X1  g1164(.A1(new_n1364), .A2(KEYINPUT63), .B1(new_n1341), .B2(new_n1344), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1341), .A2(KEYINPUT63), .A3(new_n1344), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT61), .ZN(new_n1367));
  NAND4_X1  g1167(.A1(new_n1366), .A2(new_n1356), .A3(new_n1367), .A4(new_n1360), .ZN(new_n1368));
  OAI22_X1  g1168(.A1(new_n1347), .A2(new_n1362), .B1(new_n1365), .B2(new_n1368), .ZN(G405));
  AND3_X1   g1169(.A1(new_n1309), .A2(G378), .A3(new_n1267), .ZN(new_n1370));
  AOI21_X1  g1170(.A(G378), .B1(new_n1309), .B2(new_n1267), .ZN(new_n1371));
  NOR3_X1   g1171(.A1(new_n1370), .A2(new_n1371), .A3(new_n1344), .ZN(new_n1372));
  AND3_X1   g1172(.A1(new_n1329), .A2(new_n1318), .A3(new_n893), .ZN(new_n1373));
  NOR3_X1   g1173(.A1(new_n1329), .A2(new_n1319), .A3(new_n1321), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(G375), .A2(new_n1313), .ZN(new_n1376));
  AOI21_X1  g1176(.A(new_n1375), .B1(new_n1376), .B2(new_n1337), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1372), .A2(new_n1377), .ZN(new_n1378));
  INV_X1    g1178(.A(KEYINPUT127), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1378), .B1(new_n1361), .B2(new_n1379), .ZN(new_n1380));
  NOR3_X1   g1180(.A1(new_n1353), .A2(new_n1355), .A3(new_n1349), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1358), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1382));
  OAI21_X1  g1182(.A(new_n1379), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1356), .A2(new_n1360), .A3(KEYINPUT127), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1383), .A2(new_n1384), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1380), .B1(new_n1385), .B2(new_n1378), .ZN(G402));
endmodule


