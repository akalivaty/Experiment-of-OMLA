//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n598, new_n599, new_n600, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  XOR2_X1   g029(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(new_n457), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(KEYINPUT71), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(KEYINPUT70), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n467), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n472), .A2(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI211_X1 g053(.A(new_n466), .B(new_n469), .C1(new_n478), .C2(G137), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n472), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n477), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(G137), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(KEYINPUT71), .B1(new_n482), .B2(new_n468), .ZN(new_n483));
  OR2_X1    g058(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n481), .ZN(new_n485));
  XOR2_X1   g060(.A(KEYINPUT3), .B(G2104), .Z(new_n486));
  INV_X1    g061(.A(G125), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(G113), .A2(G2104), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n484), .A2(new_n490), .ZN(G160));
  NAND2_X1  g066(.A1(new_n485), .A2(new_n480), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT72), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  OR2_X1    g069(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n480), .A2(new_n467), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n495), .A2(new_n496), .B1(G136), .B2(new_n498), .ZN(new_n499));
  OAI221_X1 g074(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n481), .C2(G112), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  AND3_X1   g077(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT3), .B1(new_n473), .B2(G2104), .ZN(new_n504));
  OAI21_X1  g079(.A(G126), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT74), .A2(G114), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT74), .A2(G114), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G2104), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n467), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n467), .A2(G102), .A3(G2104), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT75), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n516));
  OAI21_X1  g091(.A(G138), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n514), .B1(new_n486), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n480), .A2(KEYINPUT4), .A3(G138), .A4(new_n481), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G126), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n472), .B2(new_n474), .ZN(new_n522));
  NOR3_X1   g097(.A1(new_n506), .A2(new_n507), .A3(new_n471), .ZN(new_n523));
  OAI21_X1  g098(.A(G2105), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT75), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(new_n525), .A3(new_n511), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n513), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(G164));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT5), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT5), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(G62), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n529), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G651), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT76), .B1(new_n538), .B2(KEYINPUT6), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT76), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT6), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(new_n541), .A3(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n538), .A2(KEYINPUT6), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n543), .A2(G50), .A3(G543), .A4(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT5), .B(G543), .ZN(new_n546));
  NAND4_X1  g121(.A1(new_n543), .A2(G88), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n537), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(G166));
  NAND3_X1  g124(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n551), .A2(G89), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n543), .A2(new_n544), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n530), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G51), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n534), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n546), .A2(KEYINPUT77), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n562), .A2(G63), .A3(G651), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n555), .A2(new_n558), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n555), .A2(new_n566), .A3(new_n558), .A4(new_n563), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G168));
  NAND2_X1  g143(.A1(new_n557), .A2(G52), .ZN(new_n569));
  INV_X1    g144(.A(G90), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n570), .B2(new_n550), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n562), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n538), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n571), .A2(new_n573), .ZN(G301));
  INV_X1    g149(.A(G301), .ZN(G171));
  AOI22_X1  g150(.A1(new_n562), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n538), .ZN(new_n577));
  AOI22_X1  g152(.A1(G43), .A2(new_n557), .B1(new_n551), .B2(G81), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G860), .ZN(G153));
  AND3_X1   g156(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G36), .ZN(G176));
  NAND2_X1  g158(.A1(G1), .A2(G3), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT8), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(G188));
  INV_X1    g161(.A(KEYINPUT9), .ZN(new_n587));
  INV_X1    g162(.A(new_n557), .ZN(new_n588));
  INV_X1    g163(.A(G53), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G78), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G65), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n534), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n551), .A2(G91), .B1(G651), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n557), .A2(KEYINPUT9), .A3(G53), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(G299));
  INV_X1    g171(.A(G168), .ZN(G286));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n548), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n537), .A2(KEYINPUT79), .A3(new_n545), .A4(new_n547), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(G303));
  NAND2_X1  g176(.A1(new_n557), .A2(G49), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n562), .B2(G74), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n551), .A2(G87), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G288));
  NAND2_X1  g180(.A1(G73), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G61), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n534), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n543), .A2(G48), .A3(G543), .A4(new_n544), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n543), .A2(G86), .A3(new_n544), .A4(new_n546), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(G47), .A2(new_n557), .B1(new_n551), .B2(G85), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n562), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n538), .B2(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT80), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(new_n534), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n557), .A2(G54), .B1(new_n620), .B2(G651), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  OAI21_X1  g197(.A(KEYINPUT10), .B1(new_n550), .B2(new_n622), .ZN(new_n623));
  OR3_X1    g198(.A1(new_n550), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT81), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n616), .B1(new_n626), .B2(G868), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT82), .Z(G284));
  XOR2_X1   g203(.A(new_n627), .B(KEYINPUT83), .Z(G321));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NAND2_X1  g205(.A1(G299), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(G168), .B2(new_n630), .ZN(G297));
  OAI21_X1  g207(.A(new_n631), .B1(G168), .B2(new_n630), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(G860), .ZN(G148));
  NAND2_X1  g210(.A1(new_n579), .A2(new_n630), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n626), .A2(new_n634), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n636), .B1(new_n638), .B2(new_n630), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g215(.A1(new_n493), .A2(G123), .B1(G135), .B2(new_n498), .ZN(new_n641));
  OAI221_X1 g216(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n481), .C2(G111), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT85), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT13), .B(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n650), .ZN(G156));
  XOR2_X1   g226(.A(G2427), .B(G2430), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT87), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT86), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2443), .B(G2446), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1341), .B(G1348), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT88), .Z(new_n666));
  OR2_X1    g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n667), .A2(G14), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  XOR2_X1   g245(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT89), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT92), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n670), .ZN(new_n678));
  INV_X1    g253(.A(new_n675), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n679), .C1(new_n674), .C2(new_n672), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n674), .A2(new_n670), .A3(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT94), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n690), .A2(KEYINPUT94), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT20), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n687), .A2(new_n688), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  OR3_X1    g274(.A1(new_n694), .A2(new_n698), .A3(new_n690), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  INV_X1    g279(.A(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n703), .B(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G5), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G171), .B2(new_n709), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1961), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT30), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT103), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n715), .A2(new_n714), .A3(G28), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n714), .B2(G28), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n713), .B1(new_n714), .B2(G28), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n709), .A2(G19), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n580), .B2(new_n709), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G1341), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n493), .A2(G129), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n498), .A2(G141), .ZN(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT100), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT26), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n722), .A2(new_n723), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G29), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G29), .B2(G32), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n718), .B(new_n721), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT31), .B(G11), .Z(new_n734));
  NOR2_X1   g309(.A1(new_n720), .A2(G1341), .ZN(new_n735));
  OR4_X1    g310(.A1(new_n712), .A2(new_n733), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n709), .A2(G4), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n626), .B2(new_n709), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G1348), .ZN(new_n739));
  NAND2_X1  g314(.A1(G299), .A2(G16), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n709), .A2(KEYINPUT23), .A3(G20), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT23), .ZN(new_n742));
  INV_X1    g317(.A(G20), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G16), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT25), .Z(new_n749));
  INV_X1    g324(.A(G139), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n497), .A2(KEYINPUT97), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(KEYINPUT97), .B1(new_n497), .B2(new_n750), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT98), .Z(new_n754));
  INV_X1    g329(.A(G127), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n486), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G115), .B2(G2104), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(new_n481), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G29), .B2(G33), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n747), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n736), .A2(new_n739), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n644), .A2(new_n713), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT102), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n713), .A2(G26), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n493), .A2(G128), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n498), .A2(G140), .ZN(new_n769));
  OAI221_X1 g344(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n481), .C2(G116), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(new_n713), .ZN(new_n773));
  MUX2_X1   g348(.A(new_n767), .B(new_n773), .S(KEYINPUT28), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  NAND2_X1  g352(.A1(G160), .A2(G29), .ZN(new_n778));
  NOR2_X1   g353(.A1(KEYINPUT24), .A2(G34), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT24), .A2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(G29), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n778), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n731), .A2(new_n732), .B1(new_n777), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G164), .A2(new_n713), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G27), .B2(new_n713), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n761), .B2(new_n762), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n776), .A2(new_n786), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n764), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n713), .A2(G35), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G162), .B2(new_n713), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n797));
  INV_X1    g372(.A(G2090), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n796), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n709), .A2(G23), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n709), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT33), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1976), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT32), .B(G1981), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G16), .A2(G22), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G166), .B2(G16), .ZN(new_n810));
  INV_X1    g385(.A(G1971), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n805), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n709), .A2(G24), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G290), .B2(G16), .ZN(new_n816));
  MUX2_X1   g391(.A(new_n815), .B(new_n816), .S(KEYINPUT96), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1986), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n713), .A2(G25), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n493), .A2(G119), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT95), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n493), .A2(KEYINPUT95), .A3(G119), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI221_X1 g400(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n481), .C2(G107), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n498), .A2(G131), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n820), .B1(new_n829), .B2(new_n713), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT35), .B(G1991), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n830), .B(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n814), .A2(new_n818), .A3(new_n819), .A4(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT36), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n794), .B(new_n800), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n709), .A2(G21), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G168), .B2(new_n709), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT101), .B(G1966), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n785), .A2(new_n777), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n837), .A2(new_n841), .A3(new_n842), .ZN(G311));
  INV_X1    g418(.A(G311), .ZN(G150));
  XOR2_X1   g419(.A(KEYINPUT106), .B(G55), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n557), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n551), .A2(G93), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n562), .A2(G67), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT105), .B1(new_n850), .B2(G651), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(G651), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n846), .B(new_n847), .C1(new_n851), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n626), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT39), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n580), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n855), .A2(new_n580), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n861), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n857), .B1(new_n866), .B2(G860), .ZN(G145));
  XOR2_X1   g442(.A(new_n771), .B(new_n648), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n501), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n828), .A2(new_n729), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n498), .A2(G142), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT109), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n493), .A2(G130), .ZN(new_n874));
  OAI221_X1 g449(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n481), .C2(G118), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n828), .A2(new_n729), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n829), .A2(new_n728), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n870), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n759), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n524), .A2(new_n518), .A3(new_n519), .A4(new_n511), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n876), .B1(new_n871), .B2(new_n877), .ZN(new_n885));
  INV_X1    g460(.A(new_n759), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n880), .A2(new_n879), .A3(new_n870), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n882), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n884), .B1(new_n882), .B2(new_n888), .ZN(new_n891));
  XOR2_X1   g466(.A(G160), .B(KEYINPUT108), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n644), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n890), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n882), .A2(new_n888), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n883), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n893), .B1(new_n897), .B2(new_n889), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n869), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n894), .B1(new_n890), .B2(new_n891), .ZN(new_n901));
  INV_X1    g476(.A(new_n869), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(new_n889), .A3(new_n893), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g481(.A(G299), .B(new_n625), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n855), .A2(new_n580), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n862), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n911), .A2(new_n912), .A3(new_n637), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n638), .B1(new_n914), .B2(new_n910), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n907), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n637), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  INV_X1    g492(.A(new_n907), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT111), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n907), .B(new_n920), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n919), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n914), .A2(new_n910), .A3(new_n638), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n917), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(KEYINPUT112), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(KEYINPUT112), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n916), .A2(new_n930), .A3(new_n926), .ZN(new_n931));
  XNOR2_X1  g506(.A(G288), .B(new_n548), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(G305), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(G290), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(KEYINPUT112), .B2(new_n928), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n929), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n929), .B2(new_n931), .ZN(new_n938));
  OAI21_X1  g513(.A(G868), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n855), .A2(new_n630), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(G295));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n940), .ZN(G331));
  NOR2_X1   g517(.A1(new_n934), .A2(KEYINPUT114), .ZN(new_n943));
  NOR2_X1   g518(.A1(G168), .A2(KEYINPUT113), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n908), .B2(new_n862), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G301), .B1(G168), .B2(KEYINPUT113), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n908), .A2(new_n862), .A3(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n948), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n863), .A2(new_n864), .A3(new_n944), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n946), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n950), .A2(new_n923), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n907), .B1(new_n950), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n953), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n918), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n950), .A2(new_n923), .A3(new_n953), .ZN(new_n959));
  INV_X1    g534(.A(new_n943), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n961), .A3(new_n900), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n957), .A2(new_n922), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n935), .B1(new_n964), .B2(new_n955), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n958), .A2(new_n934), .A3(new_n959), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n900), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n966), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n965), .A2(KEYINPUT43), .A3(new_n900), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  MUX2_X1   g547(.A(new_n969), .B(new_n972), .S(KEYINPUT44), .Z(G397));
  INV_X1    g548(.A(KEYINPUT119), .ZN(new_n974));
  OAI211_X1 g549(.A(G40), .B(new_n490), .C1(new_n479), .C2(new_n483), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n883), .A2(KEYINPUT116), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT116), .B1(new_n883), .B2(new_n977), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n802), .A2(G1976), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(G8), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT52), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n982), .B2(KEYINPUT52), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(G305), .A2(G1981), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n609), .A2(new_n705), .A3(new_n610), .A4(new_n611), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(KEYINPUT49), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT49), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n980), .A2(G8), .A3(new_n989), .A4(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1976), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT52), .B1(G288), .B2(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n980), .A2(G8), .A3(new_n981), .A4(new_n995), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n974), .B1(new_n986), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n982), .A2(KEYINPUT52), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT118), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n982), .A2(new_n983), .A3(KEYINPUT52), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n1000), .A2(new_n997), .A3(new_n974), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n883), .A2(new_n977), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n883), .A2(KEYINPUT116), .A3(new_n977), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n527), .A2(KEYINPUT45), .A3(new_n977), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n976), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1966), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n527), .A2(new_n977), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n975), .B1(new_n1016), .B2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n978), .B2(new_n979), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n777), .A3(new_n1019), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1005), .B(G286), .C1(new_n1015), .C2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1005), .B1(new_n599), .B2(new_n600), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT50), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1018), .B1(new_n527), .B2(new_n977), .ZN(new_n1027));
  NOR4_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(G2090), .A4(new_n975), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n975), .B1(new_n1016), .B2(new_n1009), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1971), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1025), .B(G8), .C1(new_n1028), .C2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1021), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1016), .A2(new_n1009), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n976), .A3(new_n1031), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n811), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1017), .A2(new_n798), .A3(new_n1019), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1005), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT63), .B1(new_n1039), .B2(new_n1025), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1034), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT122), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1004), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1000), .A2(new_n997), .A3(new_n1001), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT119), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1002), .ZN(new_n1046));
  OAI21_X1  g621(.A(G8), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1024), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1048), .A2(KEYINPUT63), .A3(new_n1033), .A4(new_n1021), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT122), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT63), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1008), .A2(KEYINPUT50), .A3(new_n1010), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n527), .A2(new_n1018), .A3(new_n977), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n798), .A3(new_n976), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n527), .B2(new_n977), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1055), .A2(new_n975), .A3(new_n1030), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1056), .B2(G1971), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n1024), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(new_n1033), .A3(new_n997), .A4(new_n986), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1021), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1051), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1043), .A2(new_n1050), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1033), .ZN(new_n1064));
  INV_X1    g639(.A(new_n980), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(new_n1005), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n993), .A2(new_n994), .A3(new_n802), .ZN(new_n1067));
  XOR2_X1   g642(.A(new_n988), .B(KEYINPUT120), .Z(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT121), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1004), .A2(new_n1064), .B1(new_n1066), .B2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1056), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1052), .A2(new_n976), .A3(new_n1053), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n746), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(G299), .B(KEYINPUT57), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  AOI21_X1  g654(.A(G1348), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n980), .A2(G2067), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G2067), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1065), .A2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1026), .A2(new_n1027), .A3(new_n975), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT123), .B(new_n1084), .C1(new_n1085), .C2(G1348), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1077), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1073), .A2(new_n1088), .A3(new_n1075), .ZN(new_n1089));
  INV_X1    g664(.A(new_n625), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1078), .B1(new_n1087), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n625), .B1(new_n1087), .B2(KEYINPUT60), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n1094));
  AOI211_X1 g669(.A(new_n1094), .B(new_n1090), .C1(new_n1082), .C2(new_n1086), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1093), .A2(new_n1095), .B1(KEYINPUT60), .B2(new_n1087), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1089), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1088), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT61), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT61), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1078), .A2(new_n1100), .A3(new_n1089), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1036), .A2(G1996), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT58), .B(G1341), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1065), .A2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n580), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT59), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1107), .B(new_n580), .C1(new_n1102), .C2(new_n1104), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1099), .A2(new_n1101), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1092), .B1(new_n1096), .B2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1035), .A2(new_n1031), .A3(new_n789), .A4(new_n976), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1112), .A2(G2078), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1011), .A2(new_n976), .A3(new_n1012), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n976), .A3(new_n1019), .ZN(new_n1117));
  INV_X1    g692(.A(G1961), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1113), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G301), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1112), .A2(new_n1111), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT45), .B1(new_n883), .B2(new_n977), .ZN(new_n1123));
  OR3_X1    g698(.A1(new_n1123), .A2(new_n975), .A3(KEYINPUT125), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT125), .B1(new_n1123), .B2(new_n975), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1124), .A2(new_n1031), .A3(new_n1114), .A4(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(G171), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1121), .A2(new_n1127), .A3(KEYINPUT54), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT126), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1120), .A2(G171), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1113), .A2(new_n1119), .A3(G301), .A4(new_n1126), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1129), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1128), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n565), .A2(G8), .A3(new_n567), .ZN(new_n1137));
  XNOR2_X1  g712(.A(new_n1137), .B(KEYINPUT124), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1085), .A2(new_n777), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT51), .B(new_n1138), .C1(new_n1139), .C2(new_n1005), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1137), .B(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1015), .A2(new_n1020), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(G8), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1140), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1025), .B1(new_n1057), .B2(G8), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1064), .A2(new_n1044), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1136), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1063), .B(new_n1071), .C1(new_n1110), .C2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1092), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1087), .A2(KEYINPUT60), .ZN(new_n1155));
  INV_X1    g730(.A(G1348), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1117), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT123), .B1(new_n1157), .B2(new_n1084), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1080), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT60), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1090), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1087), .A2(KEYINPUT60), .A3(new_n625), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1155), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1097), .A2(new_n1098), .A3(KEYINPUT61), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1100), .B1(new_n1078), .B2(new_n1089), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1154), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1149), .A2(new_n1147), .ZN(new_n1169));
  AOI21_X1  g744(.A(G301), .B1(new_n1122), .B2(new_n1115), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1131), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT126), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT54), .B1(new_n1131), .B2(new_n1129), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1169), .B1(new_n1128), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1176), .A2(KEYINPUT127), .A3(new_n1071), .A4(new_n1063), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1060), .B1(new_n1147), .B2(KEYINPUT62), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1178), .B(new_n1170), .C1(KEYINPUT62), .C2(new_n1147), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1153), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n771), .B(new_n1083), .ZN(new_n1181));
  INV_X1    g756(.A(G1996), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n729), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n976), .A2(new_n1123), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT115), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1184), .A2(G1996), .ZN(new_n1187));
  AOI22_X1  g762(.A1(new_n1183), .A2(new_n1186), .B1(new_n729), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n829), .A2(new_n832), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n828), .A2(new_n831), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1186), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1188), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1184), .ZN(new_n1193));
  XNOR2_X1  g768(.A(G290), .B(G1986), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1180), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n772), .A2(new_n1083), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1185), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1185), .B1(new_n729), .B2(new_n1181), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1187), .B(KEYINPUT46), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT47), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1192), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1184), .A2(G1986), .A3(G290), .ZN(new_n1205));
  XOR2_X1   g780(.A(new_n1205), .B(KEYINPUT48), .Z(new_n1206));
  AOI211_X1 g781(.A(new_n1199), .B(new_n1203), .C1(new_n1204), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1196), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g783(.A(G229), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n969), .A2(G319), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g785(.A(G227), .B1(new_n666), .B2(new_n668), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n905), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1213), .ZN(G308));
  AOI21_X1  g788(.A(new_n464), .B1(new_n963), .B2(new_n968), .ZN(new_n1215));
  NAND4_X1  g789(.A1(new_n1215), .A2(new_n1210), .A3(new_n905), .A4(new_n1212), .ZN(G225));
endmodule


