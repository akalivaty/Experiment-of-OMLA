//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1338, new_n1339,
    new_n1340, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400, new_n1401,
    new_n1402, new_n1403;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT65), .Z(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n204), .A2(G50), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT66), .Z(new_n216));
  AOI21_X1  g0016(.A(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n217), .B1(KEYINPUT1), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G169), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT74), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G33), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G1698), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT76), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT76), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n254), .A2(new_n261), .A3(new_n256), .A4(new_n258), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G87), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n254), .A2(G226), .A3(G1698), .A4(new_n256), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n260), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  INV_X1    g0070(.A(G45), .ZN(new_n271));
  AOI21_X1  g0071(.A(G1), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(new_n267), .A3(G274), .ZN(new_n273));
  INV_X1    g0073(.A(G232), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n249), .B1(new_n269), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  AOI211_X1 g0081(.A(new_n281), .B(new_n278), .C1(new_n265), .C2(new_n268), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n275), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n275), .A2(G20), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n212), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT70), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n287), .A2(new_n291), .A3(KEYINPUT70), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n288), .B1(new_n296), .B2(new_n285), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n290), .A2(new_n212), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n301));
  NOR2_X1   g0101(.A1(KEYINPUT74), .A2(KEYINPUT3), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n301), .A2(new_n302), .A3(new_n255), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n251), .A2(G33), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n300), .B(new_n213), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT7), .ZN(new_n306));
  AOI21_X1  g0106(.A(G20), .B1(new_n254), .B2(new_n256), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n305), .B(G68), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G58), .ZN(new_n309));
  INV_X1    g0109(.A(G68), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(G20), .B1(new_n311), .B2(new_n203), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G20), .A2(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G159), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT16), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n298), .B1(new_n308), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(G33), .B1(new_n252), .B2(new_n253), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n320));
  OAI211_X1 g0120(.A(KEYINPUT7), .B(new_n213), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n304), .A2(new_n320), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n300), .B1(new_n322), .B2(G20), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n310), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n316), .B1(new_n324), .B2(new_n315), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n297), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(KEYINPUT18), .B1(new_n283), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT17), .ZN(new_n328));
  AOI21_X1  g0128(.A(G200), .B1(new_n269), .B2(new_n279), .ZN(new_n329));
  AOI211_X1 g0129(.A(G190), .B(new_n278), .C1(new_n265), .C2(new_n268), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n318), .A2(new_n325), .ZN(new_n332));
  INV_X1    g0132(.A(new_n288), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n298), .A2(new_n286), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n292), .A2(new_n293), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n336), .B1(new_n275), .B2(G20), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n333), .B1(new_n337), .B2(new_n284), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n328), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n278), .B1(new_n265), .B2(new_n268), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G179), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n249), .B2(new_n341), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(new_n339), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n326), .B(KEYINPUT17), .C1(new_n330), .C2(new_n329), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n327), .A2(new_n340), .A3(new_n345), .A4(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n286), .A2(G68), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT12), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n349), .B(new_n350), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n313), .A2(G50), .B1(G20), .B2(new_n310), .ZN(new_n352));
  INV_X1    g0152(.A(G77), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n213), .A2(G33), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n292), .A2(G68), .A3(new_n289), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n351), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT11), .B1(new_n355), .B2(new_n291), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G226), .ZN(new_n362));
  INV_X1    g0162(.A(G1698), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n251), .A2(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n274), .A2(G1698), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n256), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(G33), .A2(G97), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n268), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n267), .A2(G238), .A3(new_n276), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n273), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n267), .B1(new_n367), .B2(new_n368), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n273), .A2(new_n372), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT13), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(G169), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(G179), .A3(new_n377), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n379), .B1(new_n378), .B2(G169), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n361), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n371), .B1(new_n370), .B2(new_n373), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT13), .ZN(new_n386));
  OAI21_X1  g0186(.A(G200), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n374), .A2(G190), .A3(new_n377), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n387), .A2(new_n360), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT73), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(KEYINPUT73), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n348), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT72), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n213), .B1(new_n201), .B2(new_n203), .ZN(new_n395));
  INV_X1    g0195(.A(G150), .ZN(new_n396));
  INV_X1    g0196(.A(new_n313), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n284), .A2(new_n354), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n291), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G50), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n287), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n337), .A2(G50), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n273), .B1(new_n362), .B2(new_n277), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n322), .A2(G222), .A3(new_n363), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n256), .A2(new_n365), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G77), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n322), .A2(G1698), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(new_n408), .C1(new_n409), .C2(new_n257), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n405), .B1(new_n410), .B2(new_n268), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n281), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n404), .B(new_n412), .C1(G169), .C2(new_n411), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(G190), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n411), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT9), .B1(new_n402), .B2(new_n403), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n402), .A2(new_n403), .A3(KEYINPUT9), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT71), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT71), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n402), .A2(new_n403), .A3(new_n421), .A4(KEYINPUT9), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT10), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n418), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(new_n418), .B2(new_n423), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n413), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n285), .A2(new_n313), .B1(G20), .B2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n429), .A2(new_n354), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n298), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n292), .A2(G77), .A3(new_n289), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G77), .B2(new_n286), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G238), .ZN(new_n436));
  INV_X1    g0236(.A(G107), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n409), .A2(new_n436), .B1(new_n437), .B2(new_n322), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n407), .A2(new_n274), .A3(G1698), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n268), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n273), .ZN(new_n441));
  INV_X1    g0241(.A(new_n277), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(G244), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n435), .B1(new_n445), .B2(G190), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(G200), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n281), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n434), .B1(new_n444), .B2(new_n249), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n394), .B1(new_n427), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n420), .A2(new_n422), .ZN(new_n454));
  INV_X1    g0254(.A(new_n417), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n411), .A2(new_n415), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n414), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT10), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n418), .A2(new_n423), .A3(new_n424), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n452), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(KEYINPUT72), .A3(new_n413), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n393), .B1(new_n453), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n271), .A2(G1), .ZN(new_n464));
  NAND2_X1  g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G264), .A3(new_n267), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n275), .A2(G45), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(new_n465), .ZN(new_n472));
  INV_X1    g0272(.A(G274), .ZN(new_n473));
  AND2_X1   g0273(.A1(G1), .A2(G13), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n266), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(G250), .A2(G1698), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n222), .B2(G1698), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(new_n254), .A3(new_n256), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G294), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n267), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n477), .B1(new_n482), .B2(KEYINPUT84), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n301), .A2(new_n302), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n304), .B1(new_n485), .B2(G33), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(new_n479), .B1(G33), .B2(G294), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n484), .B1(new_n487), .B2(new_n267), .ZN(new_n488));
  INV_X1    g0288(.A(G190), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n469), .B(new_n476), .C1(new_n487), .C2(new_n267), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n415), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n254), .A2(new_n213), .A3(G87), .A4(new_n256), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT22), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n219), .A2(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(new_n256), .A3(new_n365), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n213), .B2(G107), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n437), .A2(KEYINPUT23), .A3(G20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G116), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(G20), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n494), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n500), .B1(new_n495), .B2(KEYINPUT22), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n511), .A2(KEYINPUT24), .A3(new_n508), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n291), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  XOR2_X1   g0313(.A(KEYINPUT83), .B(KEYINPUT25), .Z(new_n514));
  NOR2_X1   g0314(.A1(new_n286), .A2(G107), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n275), .A2(G33), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n298), .A2(new_n286), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n437), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n493), .A2(new_n513), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n502), .A2(new_n494), .A3(new_n509), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT24), .B1(new_n511), .B2(new_n508), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n298), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n520), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n249), .B1(new_n483), .B2(new_n488), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n491), .A2(new_n281), .ZN(new_n527));
  OAI22_X1  g0327(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  MUX2_X1   g0329(.A(G257), .B(G264), .S(G1698), .Z(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n254), .A3(new_n256), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n407), .A2(G303), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n267), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n468), .A2(new_n267), .ZN(new_n534));
  INV_X1    g0334(.A(G270), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n476), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR2_X1    g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G116), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n287), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n290), .A2(new_n212), .B1(G20), .B2(new_n538), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G33), .A2(G283), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n541), .B(new_n213), .C1(G33), .C2(new_n221), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(KEYINPUT20), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT20), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI221_X1 g0344(.A(new_n539), .B1(new_n518), .B2(new_n538), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n537), .A2(KEYINPUT21), .A3(G169), .A4(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  OAI21_X1  g0347(.A(G169), .B1(new_n533), .B2(new_n536), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n543), .A2(new_n544), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n539), .B1(new_n518), .B2(new_n538), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n547), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n533), .A2(new_n536), .A3(new_n281), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n545), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n546), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n533), .A2(new_n536), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n545), .B1(G190), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n415), .B2(new_n556), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT81), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n555), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(G97), .A2(G107), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(new_n219), .B1(new_n368), .B2(new_n213), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G97), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n564), .A2(new_n565), .B1(new_n354), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n254), .A2(new_n213), .A3(G68), .A4(new_n256), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n291), .ZN(new_n570));
  INV_X1    g0370(.A(new_n429), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n286), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT79), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n298), .B1(new_n567), .B2(new_n568), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT79), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n575), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n574), .A2(new_n577), .B1(new_n429), .B2(new_n518), .ZN(new_n578));
  MUX2_X1   g0378(.A(G238), .B(G244), .S(G1698), .Z(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(new_n254), .A3(new_n256), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n507), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n268), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n267), .A2(G274), .A3(new_n464), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(KEYINPUT78), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT78), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n475), .A2(new_n585), .A3(new_n464), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n464), .A2(new_n220), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n584), .A2(new_n586), .B1(new_n267), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n582), .A2(new_n281), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n267), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n267), .B1(new_n580), .B2(new_n507), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n249), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n578), .A2(new_n589), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n476), .B1(new_n534), .B2(new_n222), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n256), .A2(new_n365), .A3(G250), .A4(G1698), .ZN(new_n598));
  AND2_X1   g0398(.A1(KEYINPUT4), .A2(G244), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n256), .A2(new_n365), .A3(new_n599), .A4(new_n363), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n600), .A3(new_n541), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n254), .A2(G244), .A3(new_n363), .A4(new_n256), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n281), .B(new_n597), .C1(new_n604), .C2(new_n267), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n597), .B1(new_n604), .B2(new_n267), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n249), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n313), .A2(G77), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT6), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n609), .A2(new_n221), .A3(G107), .ZN(new_n610));
  XNOR2_X1  g0410(.A(G97), .B(G107), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n608), .B1(new_n612), .B2(new_n213), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n213), .A2(KEYINPUT7), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n255), .B1(new_n301), .B2(new_n302), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n365), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n299), .B1(new_n213), .B2(new_n407), .ZN(new_n617));
  OAI21_X1  g0417(.A(G107), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT77), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n613), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(KEYINPUT77), .B(G107), .C1(new_n616), .C2(new_n617), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n298), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n287), .A2(new_n221), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n518), .B2(new_n221), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n605), .B(new_n607), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n619), .ZN(new_n626));
  INV_X1    g0426(.A(new_n613), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n628), .B2(new_n291), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n603), .A2(new_n602), .ZN(new_n630));
  INV_X1    g0430(.A(new_n601), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n267), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n415), .B1(new_n632), .B2(new_n596), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n489), .B(new_n597), .C1(new_n604), .C2(new_n267), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n629), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n518), .A2(new_n219), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n582), .A2(new_n588), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(G200), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n570), .A2(KEYINPUT79), .A3(new_n573), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n576), .B1(new_n575), .B2(new_n572), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n582), .A2(G190), .A3(new_n588), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT80), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n582), .A2(new_n588), .A3(KEYINPUT80), .A4(G190), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n639), .A2(new_n642), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  AND4_X1   g0447(.A1(new_n595), .A2(new_n625), .A3(new_n636), .A4(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n463), .A2(new_n529), .A3(new_n562), .A4(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n413), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n341), .A2(new_n489), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(G200), .B2(new_n341), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT17), .B1(new_n652), .B2(new_n326), .ZN(new_n653));
  INV_X1    g0453(.A(new_n346), .ZN(new_n654));
  INV_X1    g0454(.A(new_n451), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n389), .ZN(new_n656));
  AOI211_X1 g0456(.A(new_n653), .B(new_n654), .C1(new_n656), .C2(new_n384), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n327), .A2(KEYINPUT87), .A3(new_n345), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT87), .B1(new_n327), .B2(new_n345), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n650), .B1(new_n661), .B2(new_n460), .ZN(new_n662));
  INV_X1    g0462(.A(new_n463), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n521), .A2(new_n625), .A3(new_n636), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT85), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n480), .A2(new_n481), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(KEYINPUT84), .A3(new_n268), .ZN(new_n667));
  INV_X1    g0467(.A(new_n477), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n670));
  OAI21_X1  g0470(.A(G169), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n534), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n482), .B1(G264), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(G179), .A3(new_n476), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n513), .A2(new_n520), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n665), .B1(new_n675), .B2(new_n555), .ZN(new_n676));
  INV_X1    g0476(.A(new_n637), .ZN(new_n677));
  OAI21_X1  g0477(.A(G200), .B1(new_n592), .B2(new_n593), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n677), .B(new_n678), .C1(new_n574), .C2(new_n577), .ZN(new_n679));
  INV_X1    g0479(.A(new_n643), .ZN(new_n680));
  INV_X1    g0480(.A(new_n518), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n640), .A2(new_n641), .B1(new_n571), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n594), .A2(new_n589), .ZN(new_n683));
  OAI22_X1  g0483(.A1(new_n679), .A2(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n546), .A2(new_n552), .A3(new_n554), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n528), .A2(new_n686), .A3(KEYINPUT85), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n664), .A2(new_n676), .A3(new_n685), .A4(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT26), .ZN(new_n689));
  OAI211_X1 g0489(.A(KEYINPUT86), .B(new_n689), .C1(new_n684), .C2(new_n625), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n632), .A2(new_n596), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n605), .B1(new_n691), .B2(G169), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n629), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(new_n595), .A3(KEYINPUT26), .A4(new_n647), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n595), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT86), .B1(new_n697), .B2(new_n689), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n688), .B(new_n595), .C1(new_n695), .C2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n662), .B1(new_n663), .B2(new_n700), .ZN(G369));
  NAND3_X1  g0501(.A1(new_n275), .A2(new_n213), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n551), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n562), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n555), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT89), .ZN(new_n712));
  OR2_X1    g0512(.A1(new_n711), .A2(KEYINPUT89), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n714), .B(new_n715), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT91), .B(G330), .Z(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n706), .B1(new_n513), .B2(new_n520), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT92), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT92), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(new_n529), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n706), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n675), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n716), .A2(new_n718), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n528), .A2(new_n723), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n686), .A2(new_n723), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n722), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n726), .A2(new_n728), .A3(new_n731), .ZN(G399));
  NAND3_X1  g0532(.A1(new_n563), .A2(new_n219), .A3(new_n538), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n208), .A2(new_n270), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(G1), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n215), .B2(new_n735), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n528), .A2(new_n686), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n664), .A2(new_n685), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n645), .A2(new_n646), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n679), .A2(new_n741), .B1(new_n682), .B2(new_n683), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n689), .B1(new_n742), .B2(new_n625), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n693), .A2(new_n595), .A3(KEYINPUT26), .A4(new_n696), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n740), .A2(new_n745), .A3(new_n595), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT29), .A3(new_n706), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n699), .A2(new_n706), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n281), .B1(new_n592), .B2(new_n593), .ZN(new_n751));
  OAI21_X1  g0551(.A(KEYINPUT93), .B1(new_n751), .B2(new_n556), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT93), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n537), .A2(new_n638), .A3(new_n753), .A4(new_n281), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n752), .A2(new_n754), .A3(new_n491), .A4(new_n606), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n592), .A2(new_n593), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n691), .A2(new_n553), .A3(new_n673), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT30), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n756), .A2(new_n673), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n760), .A2(KEYINPUT30), .A3(new_n553), .A4(new_n691), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n755), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(new_n723), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT31), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n762), .A2(new_n765), .A3(new_n723), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n562), .A2(new_n648), .A3(new_n529), .A4(new_n706), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n717), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n750), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n738), .B1(new_n774), .B2(G1), .ZN(G364));
  NOR2_X1   g0575(.A1(G13), .A2(G33), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT95), .Z(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT96), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n716), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n213), .A2(G13), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n275), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n735), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n322), .A2(new_n208), .ZN(new_n786));
  INV_X1    g0586(.A(G355), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n786), .A2(new_n787), .B1(G116), .B2(new_n208), .ZN(new_n788));
  INV_X1    g0588(.A(new_n486), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n208), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(new_n216), .B2(new_n271), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n244), .A2(G45), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n788), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n212), .B1(G20), .B2(new_n249), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n778), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n785), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n489), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n213), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n221), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n213), .A2(new_n281), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G200), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n489), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n213), .A2(G179), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(new_n489), .A3(G200), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n804), .A2(new_n400), .B1(new_n806), .B2(new_n437), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n802), .A2(G190), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n800), .B(new_n807), .C1(G68), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G190), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G159), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n813), .A2(KEYINPUT32), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n805), .A2(G190), .A3(G200), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n813), .A2(KEYINPUT32), .B1(new_n816), .B2(G87), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n801), .A2(new_n810), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n322), .B1(new_n818), .B2(new_n353), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n801), .A2(G190), .A3(new_n415), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(G58), .B2(new_n821), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n809), .A2(new_n814), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G322), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n407), .B1(new_n818), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(G329), .C2(new_n812), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n803), .A2(G326), .ZN(new_n829));
  XNOR2_X1  g0629(.A(KEYINPUT33), .B(G317), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n808), .A2(new_n830), .B1(new_n816), .B2(G303), .ZN(new_n831));
  INV_X1    g0631(.A(new_n799), .ZN(new_n832));
  INV_X1    g0632(.A(new_n806), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n832), .A2(G294), .B1(new_n833), .B2(G283), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n828), .A2(new_n829), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n823), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n797), .B1(new_n836), .B2(new_n794), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n780), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(KEYINPUT97), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT97), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n780), .A2(new_n840), .A3(new_n837), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n714), .A2(new_n715), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n714), .A2(new_n715), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n842), .A2(new_n843), .A3(new_n717), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n717), .B1(new_n842), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n785), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n839), .A2(new_n841), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G396));
  NOR2_X1   g0648(.A1(new_n451), .A2(new_n723), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n446), .A2(new_n447), .B1(new_n435), .B2(new_n723), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n655), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n700), .B2(new_n723), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT99), .ZN(new_n854));
  INV_X1    g0654(.A(new_n852), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n699), .A2(new_n706), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(KEYINPUT99), .B(new_n852), .C1(new_n700), .C2(new_n723), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n771), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(new_n858), .A3(new_n772), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n860), .B(new_n861), .C1(new_n784), .C2(new_n783), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n794), .A2(new_n776), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n785), .B1(G77), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n818), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n821), .A2(G143), .B1(new_n865), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(new_n808), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n396), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G137), .B2(new_n803), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT34), .Z(new_n870));
  NAND2_X1  g0670(.A1(new_n833), .A2(G68), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n871), .B1(new_n400), .B2(new_n815), .C1(new_n309), .C2(new_n799), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n789), .B(new_n872), .C1(G132), .C2(new_n812), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT98), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n873), .A2(KEYINPUT98), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n870), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(G283), .ZN(new_n877));
  INV_X1    g0677(.A(G303), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n867), .A2(new_n877), .B1(new_n804), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(G107), .B2(new_n816), .ZN(new_n880));
  INV_X1    g0680(.A(G294), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n820), .A2(new_n881), .B1(new_n811), .B2(new_n826), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n322), .B(new_n882), .C1(G116), .C2(new_n865), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n800), .B1(G87), .B2(new_n833), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n876), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n864), .B1(new_n886), .B2(new_n794), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n855), .B2(new_n777), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n862), .A2(new_n888), .ZN(G384));
  INV_X1    g0689(.A(new_n612), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n890), .A2(KEYINPUT35), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(KEYINPUT35), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(G116), .A3(new_n214), .A4(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(KEYINPUT100), .B(KEYINPUT36), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  OR3_X1    g0695(.A1(new_n215), .A2(new_n353), .A3(new_n311), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n201), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n275), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n856), .A2(new_n850), .ZN(new_n900));
  OAI21_X1  g0700(.A(G68), .B1(new_n307), .B2(new_n306), .ZN(new_n901));
  INV_X1    g0701(.A(new_n305), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n317), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n291), .ZN(new_n904));
  INV_X1    g0704(.A(new_n315), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT16), .B1(new_n308), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n338), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n705), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n347), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(new_n280), .B2(new_n282), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n326), .B1(new_n330), .B2(new_n329), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n908), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n318), .A2(new_n325), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n915), .A2(new_n297), .B1(new_n280), .B2(new_n282), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n339), .A2(new_n705), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT37), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n916), .A2(new_n917), .A3(new_n912), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n910), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n910), .A2(new_n920), .A3(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT102), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n360), .A2(new_n706), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n384), .A2(new_n389), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(G169), .B1(new_n385), .B2(new_n386), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT14), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n389), .A2(new_n930), .A3(new_n381), .A4(new_n380), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(KEYINPUT101), .A3(new_n926), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT101), .B1(new_n931), .B2(new_n926), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n925), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n934), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n936), .A2(KEYINPUT102), .A3(new_n928), .A4(new_n932), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n900), .A2(new_n924), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n705), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n660), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n384), .A2(new_n723), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n910), .A2(new_n920), .A3(KEYINPUT38), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NOR3_X1   g0746(.A1(new_n945), .A2(new_n921), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n916), .A2(new_n917), .A3(new_n912), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT37), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(new_n919), .ZN(new_n950));
  OAI21_X1  g0750(.A(KEYINPUT103), .B1(new_n654), .B2(new_n653), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT103), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n340), .A2(new_n952), .A3(new_n346), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(new_n658), .C2(new_n659), .ZN(new_n954));
  INV_X1    g0754(.A(new_n917), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n923), .B1(new_n956), .B2(KEYINPUT38), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n947), .B1(new_n957), .B2(new_n946), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n942), .B1(new_n944), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n463), .B(new_n747), .C1(new_n748), .C2(new_n749), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n960), .A2(new_n662), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n852), .B1(new_n935), .B2(new_n937), .ZN(new_n963));
  AND3_X1   g0763(.A1(new_n963), .A2(KEYINPUT40), .A3(new_n769), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n963), .B(new_n769), .C1(new_n945), .C2(new_n921), .ZN(new_n966));
  XNOR2_X1  g0766(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n663), .B2(new_n770), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n957), .A2(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n463), .A3(new_n769), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n718), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n962), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n275), .B2(new_n781), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n962), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n899), .B1(new_n975), .B2(new_n976), .ZN(G367));
  NOR2_X1   g0777(.A1(new_n240), .A2(new_n790), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n795), .B1(new_n208), .B2(new_n429), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n785), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n815), .A2(new_n309), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n799), .A2(new_n310), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(G159), .C2(new_n808), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n407), .B1(new_n812), .B2(G137), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G150), .A2(new_n821), .B1(new_n202), .B2(new_n865), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n803), .A2(G143), .B1(new_n833), .B2(G77), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n983), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n804), .A2(new_n826), .B1(new_n437), .B2(new_n799), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(G294), .B2(new_n808), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n820), .A2(new_n878), .B1(new_n818), .B2(new_n877), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G317), .B2(new_n812), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n486), .B1(G97), .B2(new_n833), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n815), .A2(new_n538), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n987), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n980), .B1(new_n997), .B2(new_n794), .ZN(new_n998));
  INV_X1    g0798(.A(new_n642), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n723), .B1(new_n999), .B2(new_n637), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n595), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n685), .B2(new_n1000), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n998), .B1(new_n1003), .B2(new_n779), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n625), .B(new_n636), .C1(new_n629), .C2(new_n706), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n693), .A2(new_n723), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n731), .A2(new_n728), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n731), .A2(new_n728), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1007), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT44), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND3_X1   g0813(.A1(new_n1011), .A2(KEYINPUT44), .A3(new_n1012), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1010), .B(new_n726), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT107), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n726), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1014), .A2(new_n1013), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1008), .B(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1017), .B(KEYINPUT107), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n716), .A2(new_n718), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT108), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n722), .A2(new_n724), .A3(new_n730), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n731), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1026), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n845), .B2(KEYINPUT108), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1030), .A2(new_n773), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1021), .A2(new_n1022), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n774), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n735), .B(KEYINPUT41), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n783), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n625), .B1(new_n1005), .B2(new_n528), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1037), .A2(KEYINPUT105), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(KEYINPUT105), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n706), .A3(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n722), .A2(new_n730), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n1041), .A2(KEYINPUT42), .A3(new_n1007), .ZN(new_n1042));
  AOI21_X1  g0842(.A(KEYINPUT42), .B1(new_n1041), .B2(new_n1007), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT106), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n1002), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1044), .A2(new_n1045), .A3(new_n1003), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT43), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(KEYINPUT43), .A3(new_n1044), .A4(new_n1048), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n726), .B2(new_n1012), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1051), .A2(new_n1017), .A3(new_n1007), .A4(new_n1052), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1004), .B1(new_n1036), .B2(new_n1056), .ZN(G387));
  NAND3_X1  g0857(.A1(new_n1027), .A2(new_n1029), .A3(new_n783), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n786), .A2(new_n734), .B1(G107), .B2(new_n208), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n236), .A2(G45), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n284), .A2(G50), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT50), .ZN(new_n1062));
  AOI211_X1 g0862(.A(G45), .B(new_n733), .C1(G68), .C2(G77), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n790), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1059), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT109), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n795), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n785), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n789), .B1(G97), .B2(new_n833), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n820), .A2(new_n400), .B1(new_n818), .B2(new_n310), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G150), .B2(new_n812), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n571), .A2(new_n832), .B1(new_n803), .B2(G159), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n808), .A2(new_n285), .B1(new_n816), .B2(G77), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n799), .A2(new_n877), .B1(new_n815), .B2(new_n881), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n821), .A2(G317), .B1(new_n865), .B2(G303), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(KEYINPUT110), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(KEYINPUT110), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G311), .A2(new_n808), .B1(new_n803), .B2(G322), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT48), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1076), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT49), .Z(new_n1085));
  AOI21_X1  g0885(.A(new_n486), .B1(G326), .B2(new_n812), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n538), .B2(new_n806), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1075), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1069), .B1(new_n1088), .B2(new_n794), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n725), .B2(new_n779), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1058), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n735), .B1(new_n1092), .B2(new_n774), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1030), .A2(new_n773), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(G393));
  INV_X1    g0896(.A(KEYINPUT111), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1020), .A2(new_n1097), .A3(new_n1015), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(KEYINPUT111), .A3(new_n726), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(new_n773), .C2(new_n1030), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1101), .A2(new_n1032), .A3(new_n784), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1012), .A2(new_n778), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n795), .B1(new_n221), .B2(new_n208), .C1(new_n247), .C2(new_n790), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n785), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G150), .A2(new_n803), .B1(new_n821), .B2(G159), .ZN(new_n1107));
  XOR2_X1   g0907(.A(new_n1107), .B(KEYINPUT51), .Z(new_n1108));
  AOI22_X1  g0908(.A1(new_n285), .A2(new_n865), .B1(new_n812), .B2(G143), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n799), .A2(new_n353), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n806), .A2(new_n219), .B1(new_n815), .B2(new_n310), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n202), .C2(new_n808), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1108), .A2(new_n486), .A3(new_n1109), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G317), .A2(new_n803), .B1(new_n821), .B2(G311), .ZN(new_n1114));
  XOR2_X1   g0914(.A(new_n1114), .B(KEYINPUT52), .Z(new_n1115));
  AOI22_X1  g0915(.A1(new_n832), .A2(G116), .B1(new_n865), .B2(G294), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n878), .C2(new_n867), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n407), .B1(new_n811), .B2(new_n824), .C1(new_n437), .C2(new_n806), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G283), .B2(new_n816), .ZN(new_n1119));
  XOR2_X1   g0919(.A(new_n1119), .B(KEYINPUT112), .Z(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1106), .B1(new_n1121), .B2(new_n794), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n1103), .A2(new_n783), .B1(new_n1104), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1102), .A2(new_n1123), .ZN(G390));
  INV_X1    g0924(.A(KEYINPUT38), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n340), .A2(new_n952), .A3(new_n346), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n952), .B1(new_n340), .B2(new_n346), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT87), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n283), .A2(KEYINPUT18), .A3(new_n326), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n344), .B1(new_n343), .B2(new_n339), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n327), .A2(new_n345), .A3(KEYINPUT87), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n917), .B1(new_n1128), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1125), .B1(new_n1135), .B2(new_n950), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n1136), .B2(new_n923), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n938), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n856), .B2(new_n850), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1137), .A2(new_n947), .B1(new_n944), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n771), .A2(new_n855), .A3(new_n938), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT113), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n944), .B1(new_n1136), .B2(new_n923), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n851), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n451), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n746), .A2(new_n706), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n850), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n938), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1142), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  AND4_X1   g0949(.A1(new_n1142), .A2(new_n1148), .A3(new_n957), .A4(new_n943), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1140), .B(new_n1141), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n957), .A3(new_n943), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT113), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1143), .A2(new_n1142), .A3(new_n1148), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n947), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n951), .A2(new_n953), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n955), .B1(new_n660), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n950), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n945), .B1(new_n1159), .B2(new_n1125), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1155), .B1(new_n1160), .B2(KEYINPUT39), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n1139), .A2(new_n944), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1153), .A2(new_n1154), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(G330), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n767), .B2(new_n768), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1165), .A2(new_n963), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1151), .B(new_n783), .C1(new_n1163), .C2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n785), .B1(new_n285), .B2(new_n863), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n818), .A2(new_n221), .B1(new_n811), .B2(new_n881), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n322), .B(new_n1170), .C1(G116), .C2(new_n821), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n816), .A2(G87), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n871), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1110), .B1(G283), .B2(new_n803), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n437), .B2(new_n867), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n816), .A2(G150), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT53), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(G159), .A2(new_n832), .B1(new_n803), .B2(G128), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(G137), .A2(new_n808), .B1(new_n202), .B2(new_n833), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n407), .B1(new_n812), .B2(G125), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(KEYINPUT54), .B(G143), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n821), .A2(G132), .B1(new_n865), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .A4(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1173), .A2(new_n1175), .B1(new_n1177), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1169), .B1(new_n1185), .B2(new_n794), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n958), .B2(new_n777), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1168), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT114), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT114), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1168), .A2(new_n1190), .A3(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1151), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n463), .A2(new_n1165), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n960), .A2(new_n662), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n938), .B1(new_n771), .B2(new_n855), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n900), .B1(new_n1196), .B2(new_n1166), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1165), .A2(new_n855), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1138), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1141), .A2(new_n850), .A3(new_n1146), .A4(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1195), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1193), .A2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1151), .B(new_n1201), .C1(new_n1163), .C2(new_n1167), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n784), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1192), .A2(new_n1205), .ZN(G378));
  INV_X1    g1006(.A(KEYINPUT118), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n404), .A2(new_n705), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n427), .A2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n460), .A2(new_n413), .A3(new_n1208), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1207), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1212), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n427), .A2(new_n1209), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1208), .B1(new_n460), .B2(new_n413), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(KEYINPUT118), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1215), .A2(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1222), .A2(new_n777), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n785), .B1(new_n202), .B2(new_n863), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n803), .A2(G125), .ZN(new_n1225));
  INV_X1    g1025(.A(G132), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1225), .B1(new_n867), .B2(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n821), .A2(G128), .B1(new_n865), .B2(G137), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n815), .B2(new_n1181), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(G150), .C2(new_n832), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n833), .A2(G159), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n812), .C2(G124), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n820), .A2(new_n437), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT116), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1238), .A2(new_n1239), .B1(G116), .B2(new_n803), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n309), .B2(new_n806), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n818), .A2(new_n429), .B1(new_n811), .B2(new_n877), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n1238), .A2(new_n1239), .B1(new_n867), .B2(new_n221), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(new_n1241), .A2(new_n982), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n789), .A2(new_n270), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G77), .B2(new_n816), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT115), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1246), .A2(KEYINPUT115), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  XOR2_X1   g1049(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1250));
  OR2_X1    g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1245), .B(new_n400), .C1(G33), .C2(G41), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1236), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1224), .B1(new_n1254), .B2(new_n794), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1223), .A2(new_n1255), .ZN(new_n1256));
  AND4_X1   g1056(.A1(G330), .A2(new_n1222), .A3(new_n968), .A4(new_n965), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n971), .B2(G330), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n959), .B1(new_n1257), .B2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n969), .B2(new_n1164), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1139), .A2(new_n924), .B1(new_n660), .B2(new_n940), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1161), .B2(new_n943), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n971), .A2(G330), .A3(new_n1222), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1261), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1256), .B1(new_n1267), .B2(new_n782), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1195), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1204), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1267), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT57), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1261), .A2(KEYINPUT57), .A3(new_n1266), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n735), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  AOI211_X1 g1076(.A(KEYINPUT119), .B(new_n1268), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT119), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1270), .A2(new_n1275), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1267), .B1(new_n1269), .B2(new_n1204), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1279), .B(new_n784), .C1(new_n1280), .C2(KEYINPUT57), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1268), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1277), .A2(new_n1283), .ZN(G375));
  NAND2_X1  g1084(.A1(new_n1138), .A2(new_n776), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n785), .B1(G68), .B2(new_n863), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n867), .A2(new_n538), .B1(new_n804), .B2(new_n881), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(G97), .B2(new_n816), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n833), .A2(G77), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n832), .A2(new_n571), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n820), .A2(new_n877), .B1(new_n818), .B2(new_n437), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n322), .B(new_n1291), .C1(G303), .C2(new_n812), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .A4(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n789), .B1(G58), .B2(new_n833), .ZN(new_n1294));
  INV_X1    g1094(.A(G128), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n818), .A2(new_n396), .B1(new_n811), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G137), .B2(new_n821), .ZN(new_n1297));
  AOI22_X1  g1097(.A1(new_n803), .A2(G132), .B1(new_n816), .B2(G159), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(G50), .A2(new_n832), .B1(new_n808), .B2(new_n1182), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1294), .A2(new_n1297), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1286), .B1(new_n1301), .B2(new_n794), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1285), .A2(new_n1302), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n782), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1201), .A2(new_n1034), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1195), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(G381));
  INV_X1    g1110(.A(KEYINPUT121), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1277), .B2(new_n1283), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1279), .A2(new_n784), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT57), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1282), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT119), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1281), .A2(new_n1278), .A3(new_n1282), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(KEYINPUT121), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(G378), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1095), .A2(new_n862), .A3(new_n847), .A4(new_n888), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(G390), .A2(new_n1320), .A3(G381), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1034), .B1(new_n1032), .B2(new_n774), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1054), .B(new_n1055), .C1(new_n1322), .C2(new_n783), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1321), .A2(KEYINPUT120), .A3(new_n1004), .A4(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT120), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1091), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1094), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n784), .B1(new_n1030), .B2(new_n773), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n847), .B(new_n1326), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1329), .A2(G384), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1305), .B1(new_n1308), .B2(new_n1307), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1330), .A2(new_n1102), .A3(new_n1123), .A4(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1325), .B1(G387), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1324), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1312), .A2(new_n1318), .A3(new_n1319), .A4(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT122), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1335), .B(new_n1336), .ZN(G407));
  INV_X1    g1137(.A(G343), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1312), .A2(new_n1318), .A3(new_n1338), .A4(new_n1319), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1339), .A2(G213), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1340), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT123), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(G407), .A2(KEYINPUT123), .A3(new_n1340), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(G409));
  NAND2_X1  g1147(.A1(G393), .A2(G396), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1329), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1323), .A2(new_n1004), .A3(G390), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(G390), .B1(new_n1323), .B2(new_n1004), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1349), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(G390), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(G387), .A2(new_n1354), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1355), .A2(new_n1329), .A3(new_n1348), .A4(new_n1350), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1353), .A2(new_n1356), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(G378), .A2(new_n1282), .A3(new_n1281), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1282), .B1(new_n1272), .B2(new_n1034), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1359), .A2(new_n1192), .A3(new_n1205), .ZN(new_n1360));
  AOI22_X1  g1160(.A1(new_n1358), .A2(new_n1360), .B1(G213), .B2(new_n1338), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1304), .A2(KEYINPUT60), .A3(new_n1195), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(new_n784), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1202), .A2(KEYINPUT60), .ZN(new_n1365));
  AOI21_X1  g1165(.A(new_n1364), .B1(new_n1308), .B2(new_n1365), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n862), .B(new_n888), .C1(new_n1366), .C2(new_n1305), .ZN(new_n1367));
  AND2_X1   g1167(.A1(new_n1365), .A2(new_n1308), .ZN(new_n1368));
  OAI211_X1 g1168(.A(G384), .B(new_n1306), .C1(new_n1368), .C2(new_n1364), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1367), .A2(new_n1369), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1338), .A2(G213), .A3(G2897), .ZN(new_n1371));
  XNOR2_X1  g1171(.A(new_n1370), .B(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(KEYINPUT61), .B1(new_n1362), .B2(new_n1372), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n1370), .ZN(new_n1374));
  INV_X1    g1174(.A(KEYINPUT125), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(KEYINPUT62), .ZN(new_n1376));
  OR2_X1    g1176(.A1(new_n1375), .A2(KEYINPUT62), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1361), .A2(new_n1374), .A3(new_n1376), .A4(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1373), .A2(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1361), .A2(new_n1374), .ZN(new_n1380));
  AND3_X1   g1180(.A1(new_n1380), .A2(new_n1375), .A3(KEYINPUT62), .ZN(new_n1381));
  OAI21_X1  g1181(.A(new_n1357), .B1(new_n1379), .B2(new_n1381), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1362), .A2(new_n1372), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT61), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1361), .A2(KEYINPUT63), .A3(new_n1374), .ZN(new_n1385));
  AND3_X1   g1185(.A1(new_n1383), .A2(new_n1384), .A3(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT63), .ZN(new_n1387));
  AOI21_X1  g1187(.A(new_n1357), .B1(new_n1380), .B2(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(KEYINPUT124), .B1(new_n1386), .B2(new_n1388), .ZN(new_n1389));
  AND4_X1   g1189(.A1(KEYINPUT124), .A2(new_n1388), .A3(new_n1385), .A4(new_n1373), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1382), .B1(new_n1389), .B2(new_n1390), .ZN(G405));
  NAND3_X1  g1191(.A1(new_n1316), .A2(new_n1319), .A3(new_n1317), .ZN(new_n1392));
  AND3_X1   g1192(.A1(new_n1392), .A2(KEYINPUT126), .A3(new_n1358), .ZN(new_n1393));
  NOR2_X1   g1193(.A1(new_n1392), .A2(KEYINPUT126), .ZN(new_n1394));
  OAI21_X1  g1194(.A(new_n1370), .B1(new_n1393), .B2(new_n1394), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1392), .A2(KEYINPUT126), .A3(new_n1358), .ZN(new_n1396));
  OAI211_X1 g1196(.A(new_n1396), .B(new_n1374), .C1(KEYINPUT126), .C2(new_n1392), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1395), .A2(new_n1397), .ZN(new_n1398));
  INV_X1    g1198(.A(new_n1357), .ZN(new_n1399));
  OR2_X1    g1199(.A1(new_n1399), .A2(KEYINPUT127), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1399), .A2(KEYINPUT127), .ZN(new_n1401));
  NAND3_X1  g1201(.A1(new_n1398), .A2(new_n1400), .A3(new_n1401), .ZN(new_n1402));
  NAND4_X1  g1202(.A1(new_n1395), .A2(KEYINPUT127), .A3(new_n1397), .A4(new_n1399), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1402), .A2(new_n1403), .ZN(G402));
endmodule


