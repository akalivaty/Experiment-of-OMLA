

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797;

  XNOR2_X1 U381 ( .A(G113), .B(G143), .ZN(n533) );
  XNOR2_X1 U382 ( .A(KEYINPUT76), .B(G110), .ZN(n478) );
  XNOR2_X1 U383 ( .A(KEYINPUT101), .B(KEYINPUT23), .ZN(n503) );
  XNOR2_X1 U384 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n476) );
  NAND2_X1 U385 ( .A1(G234), .A2(G237), .ZN(n486) );
  NOR2_X2 U386 ( .A1(n691), .A2(n769), .ZN(n693) );
  NOR2_X2 U387 ( .A1(n685), .A2(n769), .ZN(n687) );
  BUF_X1 U388 ( .A(G116), .Z(n411) );
  XNOR2_X2 U389 ( .A(G902), .B(KEYINPUT15), .ZN(n667) );
  NAND2_X1 U390 ( .A1(n716), .A2(n719), .ZN(n624) );
  NOR2_X1 U391 ( .A1(n662), .A2(KEYINPUT67), .ZN(n663) );
  XNOR2_X1 U392 ( .A(G140), .B(G107), .ZN(n495) );
  XNOR2_X1 U393 ( .A(G119), .B(G128), .ZN(n501) );
  INV_X1 U394 ( .A(G953), .ZN(n600) );
  XNOR2_X2 U395 ( .A(G131), .B(KEYINPUT70), .ZN(n459) );
  XNOR2_X2 U396 ( .A(n454), .B(n532), .ZN(n757) );
  NOR2_X2 U397 ( .A1(n797), .A2(n707), .ZN(n573) );
  XNOR2_X2 U398 ( .A(n363), .B(n362), .ZN(n797) );
  XNOR2_X2 U399 ( .A(n623), .B(KEYINPUT112), .ZN(n694) );
  OR2_X1 U400 ( .A1(n581), .A2(n580), .ZN(n716) );
  INV_X1 U401 ( .A(n725), .ZN(n433) );
  NOR2_X1 U402 ( .A1(n775), .A2(n679), .ZN(n725) );
  NOR2_X1 U403 ( .A1(n658), .A2(n716), .ZN(n446) );
  NOR2_X2 U404 ( .A1(G953), .A2(G237), .ZN(n536) );
  XNOR2_X1 U405 ( .A(KEYINPUT96), .B(G113), .ZN(n423) );
  INV_X1 U406 ( .A(KEYINPUT34), .ZN(n451) );
  INV_X1 U407 ( .A(KEYINPUT32), .ZN(n362) );
  NAND2_X1 U408 ( .A1(n428), .A2(n365), .ZN(n764) );
  AND2_X1 U409 ( .A1(n433), .A2(G478), .ZN(n365) );
  NOR2_X1 U410 ( .A1(n725), .A2(n726), .ZN(n462) );
  AND2_X1 U411 ( .A1(n788), .A2(n664), .ZN(n457) );
  NOR2_X1 U412 ( .A1(n796), .A2(n689), .ZN(n620) );
  NAND2_X1 U413 ( .A1(n442), .A2(n439), .ZN(n796) );
  XNOR2_X1 U414 ( .A(n446), .B(KEYINPUT40), .ZN(n689) );
  AND2_X1 U415 ( .A1(n445), .A2(n443), .ZN(n442) );
  OR2_X1 U416 ( .A1(n756), .A2(n440), .ZN(n439) );
  XNOR2_X1 U417 ( .A(n415), .B(n598), .ZN(n756) );
  OR2_X1 U418 ( .A1(n567), .A2(n382), .ZN(n455) );
  XNOR2_X1 U419 ( .A(n562), .B(n561), .ZN(n579) );
  BUF_X2 U420 ( .A(n612), .Z(n730) );
  XNOR2_X1 U421 ( .A(n548), .B(n547), .ZN(n581) );
  NOR2_X1 U422 ( .A1(n766), .A2(G902), .ZN(n518) );
  XNOR2_X1 U423 ( .A(n785), .B(n477), .ZN(n524) );
  XNOR2_X1 U424 ( .A(n522), .B(n411), .ZN(n438) );
  XNOR2_X1 U425 ( .A(n512), .B(n511), .ZN(n784) );
  XNOR2_X1 U426 ( .A(n476), .B(n553), .ZN(n785) );
  XNOR2_X1 U427 ( .A(n410), .B(n409), .ZN(n460) );
  XNOR2_X1 U428 ( .A(n425), .B(G104), .ZN(n539) );
  XNOR2_X1 U429 ( .A(n453), .B(G119), .ZN(n452) );
  XNOR2_X1 U430 ( .A(n423), .B(n472), .ZN(n422) );
  INV_X1 U431 ( .A(n769), .ZN(n361) );
  XNOR2_X2 U432 ( .A(KEYINPUT71), .B(G137), .ZN(n410) );
  XNOR2_X2 U433 ( .A(KEYINPUT97), .B(KEYINPUT81), .ZN(n467) );
  XNOR2_X2 U434 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n466) );
  INV_X1 U435 ( .A(KEYINPUT73), .ZN(n472) );
  INV_X1 U436 ( .A(KEYINPUT88), .ZN(n662) );
  INV_X4 U437 ( .A(G122), .ZN(n425) );
  NAND2_X1 U438 ( .A1(n587), .A2(n569), .ZN(n363) );
  NAND2_X1 U439 ( .A1(n593), .A2(n594), .ZN(n379) );
  XNOR2_X2 U440 ( .A(n592), .B(KEYINPUT93), .ZN(n593) );
  XNOR2_X1 U441 ( .A(n364), .B(n366), .ZN(n428) );
  XNOR2_X2 U442 ( .A(n364), .B(KEYINPUT65), .ZN(n680) );
  NAND2_X2 U443 ( .A1(n673), .A2(n672), .ZN(n364) );
  INV_X1 U444 ( .A(KEYINPUT65), .ZN(n366) );
  XNOR2_X1 U445 ( .A(n368), .B(n367), .ZN(G51) );
  INV_X1 U446 ( .A(KEYINPUT56), .ZN(n367) );
  NAND2_X1 U447 ( .A1(n369), .A2(n361), .ZN(n368) );
  XNOR2_X1 U448 ( .A(n371), .B(n370), .ZN(n369) );
  INV_X1 U449 ( .A(n699), .ZN(n370) );
  NAND2_X1 U450 ( .A1(n430), .A2(n431), .ZN(n371) );
  XNOR2_X1 U451 ( .A(n373), .B(n372), .ZN(G60) );
  INV_X1 U452 ( .A(KEYINPUT60), .ZN(n372) );
  NAND2_X1 U453 ( .A1(n374), .A2(n361), .ZN(n373) );
  XNOR2_X1 U454 ( .A(n376), .B(n375), .ZN(n374) );
  INV_X1 U455 ( .A(n763), .ZN(n375) );
  NAND2_X1 U456 ( .A1(n427), .A2(n378), .ZN(n376) );
  NAND2_X1 U457 ( .A1(n428), .A2(n377), .ZN(n767) );
  AND2_X1 U458 ( .A1(n433), .A2(G217), .ZN(n377) );
  INV_X1 U459 ( .A(n680), .ZN(n378) );
  NAND2_X1 U460 ( .A1(n594), .A2(n593), .ZN(n380) );
  NOR2_X1 U461 ( .A1(n797), .A2(n707), .ZN(n381) );
  NAND2_X1 U462 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U463 ( .A(n484), .B(n483), .ZN(n596) );
  NAND2_X1 U464 ( .A1(n596), .A2(n741), .ZN(n391) );
  AND2_X2 U465 ( .A1(n671), .A2(n670), .ZN(n673) );
  XNOR2_X1 U466 ( .A(n408), .B(n451), .ZN(n450) );
  NOR2_X2 U467 ( .A1(n394), .A2(n563), .ZN(n592) );
  XNOR2_X1 U468 ( .A(KEYINPUT10), .B(G140), .ZN(n512) );
  AND2_X1 U469 ( .A1(n742), .A2(n413), .ZN(n415) );
  NOR2_X1 U470 ( .A1(n744), .A2(n414), .ZN(n413) );
  OR2_X1 U471 ( .A1(G237), .A2(G902), .ZN(n485) );
  XOR2_X1 U472 ( .A(KEYINPUT5), .B(KEYINPUT103), .Z(n523) );
  INV_X1 U473 ( .A(G101), .ZN(n477) );
  INV_X1 U474 ( .A(G134), .ZN(n409) );
  INV_X1 U475 ( .A(KEYINPUT3), .ZN(n453) );
  NAND2_X1 U476 ( .A1(G214), .A2(n485), .ZN(n741) );
  INV_X1 U477 ( .A(G902), .ZN(n528) );
  INV_X1 U478 ( .A(n433), .ZN(n429) );
  NOR2_X1 U479 ( .A1(n629), .A2(n388), .ZN(n441) );
  NAND2_X1 U480 ( .A1(n444), .A2(n388), .ZN(n443) );
  NAND2_X1 U481 ( .A1(n448), .A2(n447), .ZN(n444) );
  XNOR2_X1 U482 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U483 ( .A(n510), .B(n465), .ZN(n474) );
  XNOR2_X1 U484 ( .A(n467), .B(n466), .ZN(n465) );
  XNOR2_X1 U485 ( .A(n678), .B(n677), .ZN(n679) );
  INV_X1 U486 ( .A(n741), .ZN(n414) );
  XNOR2_X1 U487 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U488 ( .A(n611), .B(n500), .ZN(n567) );
  XNOR2_X1 U489 ( .A(n436), .B(n524), .ZN(n526) );
  XNOR2_X1 U490 ( .A(n525), .B(n437), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n438), .B(n523), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n618), .B(n617), .ZN(n658) );
  NOR2_X1 U493 ( .A1(n581), .A2(n579), .ZN(n469) );
  BUF_X1 U494 ( .A(n567), .Z(n727) );
  XNOR2_X1 U495 ( .A(n544), .B(n543), .ZN(n762) );
  XNOR2_X1 U496 ( .A(n542), .B(n541), .ZN(n543) );
  INV_X1 U497 ( .A(KEYINPUT12), .ZN(n541) );
  NOR2_X1 U498 ( .A1(n429), .A2(n481), .ZN(n430) );
  NAND2_X1 U499 ( .A1(n448), .A2(n441), .ZN(n440) );
  AND2_X1 U500 ( .A1(n383), .A2(n611), .ZN(n435) );
  XNOR2_X1 U501 ( .A(n764), .B(n765), .ZN(n412) );
  XNOR2_X1 U502 ( .A(n417), .B(n416), .ZN(G75) );
  INV_X1 U503 ( .A(KEYINPUT53), .ZN(n416) );
  NAND2_X1 U504 ( .A1(n419), .A2(n600), .ZN(n417) );
  XNOR2_X1 U505 ( .A(n420), .B(KEYINPUT123), .ZN(n419) );
  NAND2_X1 U506 ( .A1(n609), .A2(n731), .ZN(n382) );
  INV_X1 U507 ( .A(n629), .ZN(n447) );
  NOR2_X1 U508 ( .A1(n730), .A2(n382), .ZN(n383) );
  AND2_X1 U509 ( .A1(n611), .A2(n610), .ZN(n384) );
  XNOR2_X1 U510 ( .A(KEYINPUT122), .B(n761), .ZN(n385) );
  OR2_X1 U511 ( .A1(n744), .A2(n521), .ZN(n386) );
  AND2_X1 U512 ( .A1(n469), .A2(n622), .ZN(n387) );
  XOR2_X1 U513 ( .A(n607), .B(KEYINPUT42), .Z(n388) );
  XOR2_X1 U514 ( .A(KEYINPUT92), .B(KEYINPUT35), .Z(n389) );
  XNOR2_X1 U515 ( .A(KEYINPUT2), .B(KEYINPUT85), .ZN(n390) );
  INV_X1 U516 ( .A(G210), .ZN(n481) );
  XNOR2_X2 U517 ( .A(n641), .B(KEYINPUT19), .ZN(n628) );
  XNOR2_X2 U518 ( .A(n391), .B(KEYINPUT95), .ZN(n641) );
  BUF_X1 U519 ( .A(n641), .Z(n392) );
  BUF_X1 U520 ( .A(n394), .Z(n393) );
  NAND2_X2 U521 ( .A1(n660), .A2(n468), .ZN(n675) );
  XNOR2_X2 U522 ( .A(n518), .B(n517), .ZN(n609) );
  XNOR2_X1 U523 ( .A(n449), .B(n389), .ZN(n394) );
  NAND2_X1 U524 ( .A1(n424), .A2(n525), .ZN(n397) );
  NAND2_X1 U525 ( .A1(n395), .A2(n396), .ZN(n398) );
  NAND2_X1 U526 ( .A1(n397), .A2(n398), .ZN(n770) );
  INV_X1 U527 ( .A(n424), .ZN(n395) );
  INV_X1 U528 ( .A(n525), .ZN(n396) );
  NAND2_X1 U529 ( .A1(n450), .A2(n469), .ZN(n449) );
  XNOR2_X1 U530 ( .A(n449), .B(n389), .ZN(n564) );
  XNOR2_X1 U531 ( .A(n399), .B(n400), .ZN(n685) );
  NOR2_X1 U532 ( .A1(n680), .A2(n426), .ZN(n399) );
  XOR2_X1 U533 ( .A(n683), .B(n682), .Z(n400) );
  XNOR2_X1 U534 ( .A(n401), .B(n402), .ZN(n691) );
  NOR2_X1 U535 ( .A1(n680), .A2(n432), .ZN(n401) );
  XNOR2_X1 U536 ( .A(KEYINPUT62), .B(n690), .ZN(n402) );
  XNOR2_X1 U537 ( .A(n407), .B(n493), .ZN(n403) );
  XNOR2_X1 U538 ( .A(n379), .B(KEYINPUT45), .ZN(n404) );
  XNOR2_X1 U539 ( .A(n380), .B(KEYINPUT45), .ZN(n405) );
  XNOR2_X1 U540 ( .A(n407), .B(n493), .ZN(n406) );
  XNOR2_X1 U541 ( .A(n595), .B(KEYINPUT45), .ZN(n674) );
  NAND2_X1 U542 ( .A1(n406), .A2(n757), .ZN(n408) );
  NAND2_X1 U543 ( .A1(n403), .A2(n435), .ZN(n702) );
  NOR2_X1 U544 ( .A1(n407), .A2(n386), .ZN(n463) );
  NOR2_X1 U545 ( .A1(n407), .A2(n736), .ZN(n578) );
  XNOR2_X2 U546 ( .A(n492), .B(n491), .ZN(n407) );
  NAND2_X1 U547 ( .A1(n433), .A2(G472), .ZN(n432) );
  XNOR2_X2 U548 ( .A(n786), .B(G146), .ZN(n527) );
  XOR2_X1 U549 ( .A(KEYINPUT16), .B(KEYINPUT78), .Z(n471) );
  NAND2_X1 U550 ( .A1(n674), .A2(n457), .ZN(n671) );
  INV_X2 U551 ( .A(G116), .ZN(n470) );
  XNOR2_X1 U552 ( .A(n554), .B(n425), .ZN(n555) );
  NAND2_X1 U553 ( .A1(n756), .A2(n388), .ZN(n445) );
  AND2_X2 U554 ( .A1(n591), .A2(n590), .ZN(n594) );
  NOR2_X1 U555 ( .A1(n412), .A2(n769), .ZN(G63) );
  XNOR2_X1 U556 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U557 ( .A1(n621), .A2(n387), .ZN(n623) );
  NAND2_X1 U558 ( .A1(n742), .A2(n741), .ZN(n745) );
  INV_X1 U559 ( .A(G953), .ZN(n418) );
  NAND2_X1 U560 ( .A1(n461), .A2(n385), .ZN(n420) );
  XNOR2_X1 U561 ( .A(n558), .B(n471), .ZN(n421) );
  XNOR2_X2 U562 ( .A(n470), .B(G107), .ZN(n558) );
  XNOR2_X1 U563 ( .A(n421), .B(n539), .ZN(n424) );
  XNOR2_X2 U564 ( .A(n422), .B(n452), .ZN(n525) );
  INV_X1 U565 ( .A(n680), .ZN(n431) );
  NAND2_X1 U566 ( .A1(n433), .A2(G469), .ZN(n426) );
  NOR2_X1 U567 ( .A1(n429), .A2(n545), .ZN(n427) );
  XNOR2_X1 U568 ( .A(n434), .B(KEYINPUT104), .ZN(n583) );
  NAND2_X1 U569 ( .A1(n718), .A2(n702), .ZN(n434) );
  INV_X1 U570 ( .A(n627), .ZN(n448) );
  NAND2_X1 U571 ( .A1(n577), .A2(n639), .ZN(n454) );
  XNOR2_X2 U572 ( .A(n455), .B(KEYINPUT79), .ZN(n577) );
  XNOR2_X1 U573 ( .A(n456), .B(n498), .ZN(n683) );
  XNOR2_X1 U574 ( .A(n524), .B(n479), .ZN(n498) );
  XNOR2_X1 U575 ( .A(n527), .B(n497), .ZN(n456) );
  XNOR2_X2 U576 ( .A(n675), .B(n661), .ZN(n788) );
  NAND2_X1 U577 ( .A1(n615), .A2(n384), .ZN(n458) );
  XNOR2_X2 U578 ( .A(n458), .B(n616), .ZN(n621) );
  XNOR2_X2 U579 ( .A(n460), .B(n540), .ZN(n786) );
  XNOR2_X2 U580 ( .A(n459), .B(KEYINPUT69), .ZN(n540) );
  XNOR2_X1 U581 ( .A(n462), .B(KEYINPUT89), .ZN(n461) );
  XNOR2_X1 U582 ( .A(n463), .B(n565), .ZN(n587) );
  XNOR2_X1 U583 ( .A(n393), .B(G122), .ZN(G24) );
  NAND2_X1 U584 ( .A1(n404), .A2(n788), .ZN(n464) );
  NAND2_X1 U585 ( .A1(n464), .A2(n662), .ZN(n672) );
  AND2_X1 U586 ( .A1(n464), .A2(n390), .ZN(n726) );
  AND2_X1 U587 ( .A1(n659), .A2(n688), .ZN(n468) );
  INV_X1 U588 ( .A(KEYINPUT48), .ZN(n651) );
  INV_X1 U589 ( .A(KEYINPUT30), .ZN(n613) );
  INV_X1 U590 ( .A(KEYINPUT91), .ZN(n677) );
  XOR2_X1 U591 ( .A(G146), .B(G125), .Z(n510) );
  NAND2_X1 U592 ( .A1(G224), .A2(n600), .ZN(n473) );
  XNOR2_X1 U593 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U594 ( .A(n770), .B(n475), .ZN(n480) );
  XNOR2_X2 U595 ( .A(G143), .B(G128), .ZN(n553) );
  XNOR2_X1 U596 ( .A(n478), .B(KEYINPUT75), .ZN(n479) );
  XNOR2_X1 U597 ( .A(n480), .B(n498), .ZN(n695) );
  NAND2_X1 U598 ( .A1(n695), .A2(n667), .ZN(n484) );
  INV_X1 U599 ( .A(n485), .ZN(n482) );
  NOR2_X1 U600 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U601 ( .A(n486), .B(KEYINPUT98), .ZN(n487) );
  XNOR2_X1 U602 ( .A(KEYINPUT14), .B(n487), .ZN(n488) );
  NAND2_X1 U603 ( .A1(G952), .A2(n488), .ZN(n755) );
  NOR2_X1 U604 ( .A1(G953), .A2(n755), .ZN(n603) );
  XNOR2_X1 U605 ( .A(G898), .B(KEYINPUT99), .ZN(n778) );
  NAND2_X1 U606 ( .A1(G953), .A2(n778), .ZN(n774) );
  NAND2_X1 U607 ( .A1(G902), .A2(n488), .ZN(n599) );
  NOR2_X1 U608 ( .A1(n774), .A2(n599), .ZN(n489) );
  NOR2_X1 U609 ( .A1(n603), .A2(n489), .ZN(n490) );
  NOR2_X2 U610 ( .A1(n628), .A2(n490), .ZN(n492) );
  INV_X1 U611 ( .A(KEYINPUT0), .ZN(n491) );
  INV_X1 U612 ( .A(KEYINPUT100), .ZN(n493) );
  NAND2_X1 U613 ( .A1(n600), .A2(G227), .ZN(n494) );
  XNOR2_X1 U614 ( .A(n494), .B(G104), .ZN(n496) );
  XNOR2_X1 U615 ( .A(n496), .B(n495), .ZN(n497) );
  OR2_X2 U616 ( .A1(n683), .A2(G902), .ZN(n499) );
  XNOR2_X2 U617 ( .A(n499), .B(G469), .ZN(n611) );
  INV_X1 U618 ( .A(KEYINPUT1), .ZN(n500) );
  XOR2_X1 U619 ( .A(G110), .B(G137), .Z(n502) );
  XNOR2_X1 U620 ( .A(n502), .B(n501), .ZN(n506) );
  XOR2_X1 U621 ( .A(KEYINPUT24), .B(KEYINPUT74), .Z(n504) );
  XNOR2_X1 U622 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U623 ( .A(n506), .B(n505), .Z(n509) );
  NAND2_X1 U624 ( .A1(G234), .A2(n418), .ZN(n507) );
  XOR2_X1 U625 ( .A(KEYINPUT8), .B(n507), .Z(n550) );
  NAND2_X1 U626 ( .A1(G221), .A2(n550), .ZN(n508) );
  XNOR2_X1 U627 ( .A(n509), .B(n508), .ZN(n513) );
  INV_X1 U628 ( .A(n510), .ZN(n511) );
  XNOR2_X1 U629 ( .A(n513), .B(n784), .ZN(n766) );
  NAND2_X1 U630 ( .A1(n667), .A2(G234), .ZN(n514) );
  XNOR2_X1 U631 ( .A(n514), .B(KEYINPUT20), .ZN(n519) );
  NAND2_X1 U632 ( .A1(n519), .A2(G217), .ZN(n516) );
  XNOR2_X1 U633 ( .A(KEYINPUT102), .B(KEYINPUT25), .ZN(n515) );
  XNOR2_X1 U634 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U635 ( .A1(n519), .A2(G221), .ZN(n520) );
  XNOR2_X1 U636 ( .A(n520), .B(KEYINPUT21), .ZN(n521) );
  INV_X1 U637 ( .A(n521), .ZN(n731) );
  NAND2_X1 U638 ( .A1(n536), .A2(G210), .ZN(n522) );
  XNOR2_X1 U639 ( .A(n527), .B(n526), .ZN(n690) );
  NAND2_X1 U640 ( .A1(n690), .A2(n528), .ZN(n529) );
  XNOR2_X2 U641 ( .A(n529), .B(G472), .ZN(n612) );
  INV_X1 U642 ( .A(KEYINPUT6), .ZN(n530) );
  XNOR2_X1 U643 ( .A(n730), .B(n530), .ZN(n639) );
  INV_X1 U644 ( .A(KEYINPUT77), .ZN(n531) );
  XNOR2_X1 U645 ( .A(n531), .B(KEYINPUT33), .ZN(n532) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(KEYINPUT105), .Z(n534) );
  XNOR2_X1 U647 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U648 ( .A(n784), .B(n535), .ZN(n538) );
  NAND2_X1 U649 ( .A1(G214), .A2(n536), .ZN(n537) );
  XNOR2_X1 U650 ( .A(n538), .B(n537), .ZN(n544) );
  XNOR2_X1 U651 ( .A(n540), .B(n539), .ZN(n542) );
  NOR2_X1 U652 ( .A1(G902), .A2(n762), .ZN(n548) );
  XNOR2_X1 U653 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n546) );
  INV_X1 U654 ( .A(G475), .ZN(n545) );
  XOR2_X1 U655 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n549) );
  XNOR2_X1 U656 ( .A(G478), .B(n549), .ZN(n562) );
  XOR2_X1 U657 ( .A(KEYINPUT107), .B(KEYINPUT7), .Z(n552) );
  NAND2_X1 U658 ( .A1(G217), .A2(n550), .ZN(n551) );
  XNOR2_X1 U659 ( .A(n552), .B(n551), .ZN(n556) );
  XOR2_X1 U660 ( .A(n553), .B(G134), .Z(n554) );
  XNOR2_X1 U661 ( .A(KEYINPUT9), .B(n557), .ZN(n560) );
  INV_X1 U662 ( .A(n558), .ZN(n559) );
  XNOR2_X1 U663 ( .A(n560), .B(n559), .ZN(n765) );
  NOR2_X1 U664 ( .A1(G902), .A2(n765), .ZN(n561) );
  INV_X1 U665 ( .A(KEYINPUT44), .ZN(n563) );
  NAND2_X1 U666 ( .A1(n564), .A2(n563), .ZN(n572) );
  NAND2_X1 U667 ( .A1(n579), .A2(n581), .ZN(n744) );
  XNOR2_X1 U668 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n565) );
  XNOR2_X1 U669 ( .A(KEYINPUT110), .B(n609), .ZN(n732) );
  XNOR2_X1 U670 ( .A(n639), .B(KEYINPUT82), .ZN(n566) );
  NOR2_X1 U671 ( .A1(n732), .A2(n566), .ZN(n568) );
  INV_X1 U672 ( .A(n727), .ZN(n644) );
  AND2_X1 U673 ( .A1(n568), .A2(n644), .ZN(n569) );
  NOR2_X1 U674 ( .A1(n730), .A2(n609), .ZN(n570) );
  AND2_X1 U675 ( .A1(n727), .A2(n570), .ZN(n571) );
  AND2_X1 U676 ( .A1(n587), .A2(n571), .ZN(n707) );
  NAND2_X1 U677 ( .A1(n572), .A2(n381), .ZN(n576) );
  INV_X1 U678 ( .A(n573), .ZN(n574) );
  NAND2_X1 U679 ( .A1(n574), .A2(n563), .ZN(n575) );
  NAND2_X1 U680 ( .A1(n576), .A2(n575), .ZN(n591) );
  NAND2_X1 U681 ( .A1(n577), .A2(n730), .ZN(n736) );
  XNOR2_X1 U682 ( .A(n578), .B(KEYINPUT31), .ZN(n718) );
  INV_X1 U683 ( .A(n579), .ZN(n580) );
  NAND2_X1 U684 ( .A1(n581), .A2(n580), .ZN(n719) );
  INV_X1 U685 ( .A(KEYINPUT87), .ZN(n582) );
  XNOR2_X1 U686 ( .A(n624), .B(n582), .ZN(n636) );
  NAND2_X1 U687 ( .A1(n583), .A2(n636), .ZN(n588) );
  INV_X1 U688 ( .A(n732), .ZN(n584) );
  OR2_X1 U689 ( .A1(n584), .A2(n639), .ZN(n585) );
  NOR2_X1 U690 ( .A1(n585), .A2(n644), .ZN(n586) );
  NAND2_X1 U691 ( .A1(n587), .A2(n586), .ZN(n700) );
  NAND2_X1 U692 ( .A1(n588), .A2(n700), .ZN(n589) );
  XNOR2_X1 U693 ( .A(n589), .B(KEYINPUT111), .ZN(n590) );
  BUF_X1 U694 ( .A(n596), .Z(n622) );
  INV_X1 U695 ( .A(KEYINPUT38), .ZN(n597) );
  XNOR2_X1 U696 ( .A(n622), .B(n597), .ZN(n742) );
  XNOR2_X1 U697 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n598) );
  OR2_X1 U698 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U699 ( .A1(n601), .A2(G900), .ZN(n602) );
  OR2_X1 U700 ( .A1(n603), .A2(n602), .ZN(n604) );
  AND2_X1 U701 ( .A1(n604), .A2(n731), .ZN(n608) );
  XOR2_X1 U702 ( .A(n608), .B(KEYINPUT72), .Z(n605) );
  NOR2_X1 U703 ( .A1(n609), .A2(n605), .ZN(n638) );
  AND2_X1 U704 ( .A1(n730), .A2(n638), .ZN(n606) );
  XOR2_X1 U705 ( .A(KEYINPUT28), .B(n606), .Z(n627) );
  XNOR2_X1 U706 ( .A(n611), .B(KEYINPUT113), .ZN(n629) );
  INV_X1 U707 ( .A(KEYINPUT115), .ZN(n607) );
  AND2_X1 U708 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U709 ( .A1(n612), .A2(n741), .ZN(n614) );
  INV_X1 U710 ( .A(KEYINPUT80), .ZN(n616) );
  NAND2_X1 U711 ( .A1(n621), .A2(n742), .ZN(n618) );
  INV_X1 U712 ( .A(KEYINPUT39), .ZN(n617) );
  XNOR2_X1 U713 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n619) );
  XNOR2_X1 U714 ( .A(n620), .B(n619), .ZN(n650) );
  INV_X1 U715 ( .A(n624), .ZN(n746) );
  NAND2_X1 U716 ( .A1(n746), .A2(KEYINPUT47), .ZN(n625) );
  NAND2_X1 U717 ( .A1(n694), .A2(n625), .ZN(n626) );
  XNOR2_X1 U718 ( .A(n626), .B(KEYINPUT83), .ZN(n633) );
  NOR2_X1 U719 ( .A1(n627), .A2(n628), .ZN(n630) );
  AND2_X1 U720 ( .A1(n630), .A2(n447), .ZN(n713) );
  INV_X1 U721 ( .A(n713), .ZN(n631) );
  NAND2_X1 U722 ( .A1(n631), .A2(KEYINPUT47), .ZN(n632) );
  NAND2_X1 U723 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U724 ( .A(n634), .B(KEYINPUT86), .ZN(n648) );
  INV_X1 U725 ( .A(KEYINPUT47), .ZN(n635) );
  AND2_X1 U726 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n713), .A2(n637), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U729 ( .A1(n716), .A2(n640), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n653), .A2(n392), .ZN(n643) );
  XOR2_X1 U731 ( .A(KEYINPUT94), .B(KEYINPUT36), .Z(n642) );
  XNOR2_X1 U732 ( .A(n643), .B(n642), .ZN(n645) );
  NAND2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n722) );
  NAND2_X1 U734 ( .A1(n646), .A2(n722), .ZN(n647) );
  NOR2_X1 U735 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n652) );
  XNOR2_X1 U737 ( .A(n652), .B(n651), .ZN(n660) );
  AND2_X1 U738 ( .A1(n653), .A2(n741), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n654), .A2(n727), .ZN(n655) );
  XNOR2_X1 U740 ( .A(n655), .B(KEYINPUT43), .ZN(n657) );
  INV_X1 U741 ( .A(n622), .ZN(n656) );
  AND2_X1 U742 ( .A1(n657), .A2(n656), .ZN(n724) );
  INV_X1 U743 ( .A(n724), .ZN(n659) );
  OR2_X1 U744 ( .A1(n658), .A2(n719), .ZN(n688) );
  INV_X1 U745 ( .A(KEYINPUT90), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n667), .A2(n663), .ZN(n665) );
  AND2_X1 U747 ( .A1(KEYINPUT88), .A2(n665), .ZN(n664) );
  INV_X1 U748 ( .A(n665), .ZN(n669) );
  XOR2_X1 U749 ( .A(KEYINPUT2), .B(KEYINPUT67), .Z(n666) );
  NOR2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n668) );
  OR2_X1 U751 ( .A1(n669), .A2(n668), .ZN(n670) );
  INV_X1 U752 ( .A(n405), .ZN(n775) );
  INV_X1 U753 ( .A(n675), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n676), .A2(KEYINPUT2), .ZN(n678) );
  XOR2_X1 U755 ( .A(KEYINPUT124), .B(KEYINPUT57), .Z(n681) );
  XNOR2_X1 U756 ( .A(n681), .B(KEYINPUT58), .ZN(n682) );
  INV_X1 U757 ( .A(G952), .ZN(n684) );
  AND2_X1 U758 ( .A1(n684), .A2(G953), .ZN(n769) );
  INV_X1 U759 ( .A(KEYINPUT125), .ZN(n686) );
  XNOR2_X1 U760 ( .A(n687), .B(n686), .ZN(G54) );
  XNOR2_X1 U761 ( .A(n688), .B(G134), .ZN(G36) );
  XOR2_X1 U762 ( .A(G131), .B(n689), .Z(G33) );
  XOR2_X1 U763 ( .A(KEYINPUT116), .B(KEYINPUT63), .Z(n692) );
  XNOR2_X1 U764 ( .A(n693), .B(n692), .ZN(G57) );
  XNOR2_X1 U765 ( .A(n694), .B(G143), .ZN(G45) );
  BUF_X1 U766 ( .A(n695), .Z(n696) );
  XNOR2_X1 U767 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n697) );
  XNOR2_X1 U768 ( .A(n697), .B(KEYINPUT55), .ZN(n698) );
  XNOR2_X1 U769 ( .A(n696), .B(n698), .ZN(n699) );
  XNOR2_X1 U770 ( .A(G101), .B(n700), .ZN(G3) );
  NOR2_X1 U771 ( .A1(n716), .A2(n702), .ZN(n701) );
  XOR2_X1 U772 ( .A(G104), .B(n701), .Z(G6) );
  NOR2_X1 U773 ( .A1(n719), .A2(n702), .ZN(n706) );
  XOR2_X1 U774 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n704) );
  XNOR2_X1 U775 ( .A(G107), .B(KEYINPUT117), .ZN(n703) );
  XNOR2_X1 U776 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U777 ( .A(n706), .B(n705), .ZN(G9) );
  XOR2_X1 U778 ( .A(G110), .B(n707), .Z(n708) );
  XNOR2_X1 U779 ( .A(KEYINPUT118), .B(n708), .ZN(G12) );
  XOR2_X1 U780 ( .A(G128), .B(KEYINPUT29), .Z(n711) );
  INV_X1 U781 ( .A(n719), .ZN(n709) );
  NAND2_X1 U782 ( .A1(n713), .A2(n709), .ZN(n710) );
  XNOR2_X1 U783 ( .A(n711), .B(n710), .ZN(G30) );
  XOR2_X1 U784 ( .A(G146), .B(KEYINPUT119), .Z(n715) );
  INV_X1 U785 ( .A(n716), .ZN(n712) );
  NAND2_X1 U786 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U787 ( .A(n715), .B(n714), .ZN(G48) );
  NOR2_X1 U788 ( .A1(n716), .A2(n718), .ZN(n717) );
  XOR2_X1 U789 ( .A(G113), .B(n717), .Z(G15) );
  NOR2_X1 U790 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U791 ( .A(KEYINPUT120), .B(n720), .Z(n721) );
  XNOR2_X1 U792 ( .A(n411), .B(n721), .ZN(G18) );
  XOR2_X1 U793 ( .A(G125), .B(n722), .Z(n723) );
  XNOR2_X1 U794 ( .A(n723), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U795 ( .A(G140), .B(n724), .Z(G42) );
  NAND2_X1 U796 ( .A1(n727), .A2(n382), .ZN(n728) );
  XOR2_X1 U797 ( .A(KEYINPUT50), .B(n728), .Z(n729) );
  NOR2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n735) );
  NOR2_X1 U799 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U800 ( .A(n733), .B(KEYINPUT49), .ZN(n734) );
  NAND2_X1 U801 ( .A1(n735), .A2(n734), .ZN(n737) );
  NAND2_X1 U802 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U803 ( .A(KEYINPUT51), .B(n738), .ZN(n739) );
  NOR2_X1 U804 ( .A1(n756), .A2(n739), .ZN(n740) );
  XOR2_X1 U805 ( .A(KEYINPUT121), .B(n740), .Z(n752) );
  INV_X1 U806 ( .A(n757), .ZN(n750) );
  NOR2_X1 U807 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U808 ( .A1(n744), .A2(n743), .ZN(n748) );
  NOR2_X1 U809 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U810 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U811 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U812 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U813 ( .A(n753), .B(KEYINPUT52), .ZN(n754) );
  NOR2_X1 U814 ( .A1(n755), .A2(n754), .ZN(n760) );
  INV_X1 U815 ( .A(n756), .ZN(n758) );
  AND2_X1 U816 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U817 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U818 ( .A(n762), .B(KEYINPUT59), .Z(n763) );
  XNOR2_X1 U819 ( .A(n767), .B(n766), .ZN(n768) );
  NOR2_X1 U820 ( .A1(n769), .A2(n768), .ZN(G66) );
  BUF_X1 U821 ( .A(n770), .Z(n772) );
  XOR2_X1 U822 ( .A(G101), .B(G110), .Z(n771) );
  XNOR2_X1 U823 ( .A(n772), .B(n771), .ZN(n773) );
  NAND2_X1 U824 ( .A1(n774), .A2(n773), .ZN(n783) );
  NOR2_X1 U825 ( .A1(n775), .A2(G953), .ZN(n781) );
  XOR2_X1 U826 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n777) );
  NAND2_X1 U827 ( .A1(G224), .A2(G953), .ZN(n776) );
  XNOR2_X1 U828 ( .A(n777), .B(n776), .ZN(n779) );
  NOR2_X1 U829 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U830 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U831 ( .A(n783), .B(n782), .ZN(G69) );
  XNOR2_X1 U832 ( .A(n785), .B(n784), .ZN(n787) );
  XNOR2_X1 U833 ( .A(n787), .B(n786), .ZN(n791) );
  XNOR2_X1 U834 ( .A(n788), .B(n791), .ZN(n789) );
  NOR2_X1 U835 ( .A1(n789), .A2(G953), .ZN(n790) );
  XNOR2_X1 U836 ( .A(n790), .B(KEYINPUT127), .ZN(n795) );
  XNOR2_X1 U837 ( .A(G227), .B(n791), .ZN(n792) );
  NAND2_X1 U838 ( .A1(n792), .A2(G900), .ZN(n793) );
  NAND2_X1 U839 ( .A1(n793), .A2(G953), .ZN(n794) );
  NAND2_X1 U840 ( .A1(n795), .A2(n794), .ZN(G72) );
  XOR2_X1 U841 ( .A(n796), .B(G137), .Z(G39) );
  XOR2_X1 U842 ( .A(n797), .B(G119), .Z(G21) );
endmodule

