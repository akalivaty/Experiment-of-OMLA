

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770;

  BUF_X1 U369 ( .A(n654), .Z(n354) );
  NAND2_X1 U370 ( .A1(n350), .A2(n423), .ZN(n418) );
  NAND2_X1 U371 ( .A1(n425), .A2(n426), .ZN(n350) );
  XNOR2_X2 U372 ( .A(n499), .B(n449), .ZN(n514) );
  NOR2_X2 U373 ( .A1(n352), .A2(n351), .ZN(n568) );
  INV_X1 U374 ( .A(n417), .ZN(n351) );
  NAND2_X1 U375 ( .A1(n353), .A2(n371), .ZN(n352) );
  INV_X1 U376 ( .A(n760), .ZN(n353) );
  XNOR2_X1 U377 ( .A(n464), .B(n465), .ZN(n497) );
  XNOR2_X1 U378 ( .A(n621), .B(n380), .ZN(n678) );
  XNOR2_X2 U379 ( .A(n584), .B(KEYINPUT107), .ZN(n761) );
  NOR2_X2 U380 ( .A1(n608), .A2(n442), .ZN(n441) );
  XNOR2_X2 U381 ( .A(n593), .B(KEYINPUT41), .ZN(n676) );
  NAND2_X2 U382 ( .A1(n386), .A2(n385), .ZN(n593) );
  XNOR2_X1 U383 ( .A(n439), .B(n438), .ZN(n662) );
  XNOR2_X2 U384 ( .A(G113), .B(G119), .ZN(n463) );
  NOR2_X1 U385 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U386 ( .A1(n767), .A2(n766), .ZN(n602) );
  OR2_X1 U387 ( .A1(n759), .A2(KEYINPUT44), .ZN(n550) );
  XNOR2_X1 U388 ( .A(n548), .B(n370), .ZN(n759) );
  XNOR2_X1 U389 ( .A(n540), .B(KEYINPUT32), .ZN(n765) );
  XNOR2_X1 U390 ( .A(n591), .B(KEYINPUT40), .ZN(n767) );
  OR2_X1 U391 ( .A1(n553), .A2(n539), .ZN(n540) );
  XNOR2_X1 U392 ( .A(n363), .B(KEYINPUT22), .ZN(n553) );
  AND2_X1 U393 ( .A1(n651), .A2(n615), .ZN(n591) );
  XNOR2_X1 U394 ( .A(n546), .B(n454), .ZN(n687) );
  NAND2_X1 U395 ( .A1(n406), .A2(n402), .ZN(n608) );
  NOR2_X1 U396 ( .A1(n408), .A2(n407), .ZN(n406) );
  NAND2_X2 U397 ( .A1(n401), .A2(n405), .ZN(n621) );
  XNOR2_X1 U398 ( .A(n599), .B(n481), .ZN(n545) );
  NOR2_X1 U399 ( .A1(n663), .A2(n662), .ZN(n666) );
  OR2_X1 U400 ( .A1(n702), .A2(n400), .ZN(n397) );
  XNOR2_X1 U401 ( .A(n702), .B(n703), .ZN(n704) );
  XNOR2_X1 U402 ( .A(n379), .B(n504), .ZN(n702) );
  XNOR2_X1 U403 ( .A(n521), .B(n430), .ZN(n722) );
  XNOR2_X1 U404 ( .A(n503), .B(n355), .ZN(n504) );
  XNOR2_X1 U405 ( .A(n730), .B(n500), .ZN(n379) );
  XNOR2_X1 U406 ( .A(n497), .B(n496), .ZN(n730) );
  XNOR2_X1 U407 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U408 ( .A(n461), .B(KEYINPUT70), .ZN(n465) );
  AND2_X4 U409 ( .A1(n715), .A2(n713), .ZN(n711) );
  NAND2_X2 U410 ( .A1(n628), .A2(n627), .ZN(n715) );
  NOR2_X1 U411 ( .A1(G902), .A2(G237), .ZN(n506) );
  NAND2_X1 U412 ( .A1(n446), .A2(n505), .ZN(n416) );
  INV_X1 U413 ( .A(KEYINPUT76), .ZN(n509) );
  NOR2_X1 U414 ( .A1(n411), .A2(n510), .ZN(n410) );
  INV_X1 U415 ( .A(KEYINPUT38), .ZN(n380) );
  INV_X1 U416 ( .A(n545), .ZN(n665) );
  AND2_X1 U417 ( .A1(n768), .A2(n623), .ZN(n624) );
  XNOR2_X1 U418 ( .A(n441), .B(n440), .ZN(n558) );
  INV_X1 U419 ( .A(KEYINPUT0), .ZN(n440) );
  NAND2_X1 U420 ( .A1(n361), .A2(n693), .ZN(n442) );
  NAND2_X1 U421 ( .A1(n422), .A2(n421), .ZN(n420) );
  NAND2_X1 U422 ( .A1(n589), .A2(KEYINPUT91), .ZN(n421) );
  XOR2_X1 U423 ( .A(KEYINPUT69), .B(G131), .Z(n531) );
  NAND2_X1 U424 ( .A1(n414), .A2(n625), .ZN(n413) );
  XOR2_X1 U425 ( .A(G137), .B(G140), .Z(n482) );
  INV_X1 U426 ( .A(G134), .ZN(n449) );
  XNOR2_X1 U427 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n486) );
  INV_X1 U428 ( .A(n595), .ZN(n365) );
  NAND2_X1 U429 ( .A1(n398), .A2(n416), .ZN(n415) );
  NAND2_X1 U430 ( .A1(n702), .A2(n446), .ZN(n398) );
  NAND2_X1 U431 ( .A1(n411), .A2(n510), .ZN(n409) );
  NAND2_X1 U432 ( .A1(n358), .A2(n397), .ZN(n396) );
  AND2_X1 U433 ( .A1(n412), .A2(n410), .ZN(n407) );
  INV_X1 U434 ( .A(n412), .ZN(n405) );
  XNOR2_X1 U435 ( .A(KEYINPUT88), .B(n559), .ZN(n589) );
  XNOR2_X1 U436 ( .A(n558), .B(KEYINPUT87), .ZN(n561) );
  XNOR2_X1 U437 ( .A(G128), .B(G110), .ZN(n483) );
  XNOR2_X1 U438 ( .A(n501), .B(n433), .ZN(n745) );
  XNOR2_X1 U439 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n433) );
  XNOR2_X1 U440 ( .A(G116), .B(G107), .ZN(n522) );
  INV_X1 U441 ( .A(KEYINPUT96), .ZN(n432) );
  XNOR2_X1 U442 ( .A(G122), .B(KEYINPUT95), .ZN(n515) );
  XOR2_X1 U443 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n516) );
  XNOR2_X1 U444 ( .A(n743), .B(n459), .ZN(n708) );
  XNOR2_X1 U445 ( .A(n503), .B(n357), .ZN(n459) );
  XNOR2_X1 U446 ( .A(G146), .B(G125), .ZN(n501) );
  INV_X1 U447 ( .A(KEYINPUT33), .ZN(n454) );
  NOR2_X1 U448 ( .A1(n394), .A2(n448), .ZN(n659) );
  OR2_X1 U449 ( .A1(n580), .A2(n367), .ZN(n618) );
  INV_X1 U450 ( .A(n681), .ZN(n385) );
  INV_X1 U451 ( .A(n682), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n590), .B(KEYINPUT39), .ZN(n615) );
  NOR2_X1 U453 ( .A1(n585), .A2(n618), .ZN(n582) );
  INV_X1 U454 ( .A(n621), .ZN(n585) );
  INV_X1 U455 ( .A(KEYINPUT34), .ZN(n452) );
  NOR2_X1 U456 ( .A1(n597), .A2(n596), .ZN(n598) );
  INV_X1 U457 ( .A(KEYINPUT1), .ZN(n481) );
  NOR2_X1 U458 ( .A1(n722), .A2(G902), .ZN(n523) );
  NAND2_X1 U459 ( .A1(n428), .A2(n429), .ZN(n363) );
  OR2_X1 U460 ( .A1(n727), .A2(G902), .ZN(n439) );
  XNOR2_X1 U461 ( .A(n492), .B(KEYINPUT25), .ZN(n438) );
  BUF_X1 U462 ( .A(n665), .Z(n372) );
  INV_X1 U463 ( .A(G953), .ZN(n755) );
  NOR2_X1 U464 ( .A1(n769), .A2(n611), .ZN(n612) );
  INV_X1 U465 ( .A(KEYINPUT47), .ZN(n376) );
  NOR2_X1 U466 ( .A1(G953), .A2(G237), .ZN(n469) );
  NAND2_X1 U467 ( .A1(G953), .A2(G902), .ZN(n572) );
  INV_X1 U468 ( .A(KEYINPUT86), .ZN(n447) );
  INV_X1 U469 ( .A(n679), .ZN(n411) );
  NAND2_X1 U470 ( .A1(n416), .A2(n414), .ZN(n399) );
  INV_X1 U471 ( .A(n416), .ZN(n400) );
  XNOR2_X1 U472 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n466) );
  XOR2_X1 U473 ( .A(G146), .B(G137), .Z(n467) );
  XNOR2_X1 U474 ( .A(n514), .B(n471), .ZN(n478) );
  INV_X1 U475 ( .A(KEYINPUT48), .ZN(n374) );
  XNOR2_X1 U476 ( .A(n445), .B(KEYINPUT66), .ZN(n747) );
  INV_X1 U477 ( .A(KEYINPUT4), .ZN(n445) );
  NOR2_X1 U478 ( .A1(n392), .A2(n394), .ZN(n391) );
  NAND2_X1 U479 ( .A1(n505), .A2(n395), .ZN(n393) );
  NAND2_X1 U480 ( .A1(n625), .A2(KEYINPUT78), .ZN(n389) );
  XOR2_X1 U481 ( .A(G104), .B(G140), .Z(n526) );
  XNOR2_X1 U482 ( .A(G143), .B(G113), .ZN(n525) );
  XNOR2_X1 U483 ( .A(G122), .B(KEYINPUT12), .ZN(n527) );
  XOR2_X1 U484 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n528) );
  XNOR2_X1 U485 ( .A(n478), .B(n477), .ZN(n743) );
  INV_X1 U486 ( .A(n482), .ZN(n477) );
  XNOR2_X1 U487 ( .A(n747), .B(n472), .ZN(n479) );
  XNOR2_X1 U488 ( .A(KEYINPUT65), .B(G101), .ZN(n472) );
  XNOR2_X1 U489 ( .A(n592), .B(KEYINPUT106), .ZN(n682) );
  NOR2_X1 U490 ( .A1(n663), .A2(n681), .ZN(n538) );
  XNOR2_X1 U491 ( .A(n444), .B(n443), .ZN(n731) );
  INV_X1 U492 ( .A(G110), .ZN(n443) );
  XNOR2_X1 U493 ( .A(G107), .B(G104), .ZN(n444) );
  XOR2_X1 U494 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n498) );
  XNOR2_X1 U495 ( .A(n479), .B(n731), .ZN(n503) );
  NAND2_X1 U496 ( .A1(G234), .A2(G237), .ZN(n494) );
  INV_X1 U497 ( .A(n415), .ZN(n401) );
  AND2_X1 U498 ( .A1(n588), .A2(n364), .ZN(n604) );
  NOR2_X1 U499 ( .A1(n589), .A2(n365), .ZN(n364) );
  NAND2_X1 U500 ( .A1(n405), .A2(n403), .ZN(n402) );
  NOR2_X1 U501 ( .A1(n415), .A2(n404), .ZN(n403) );
  XNOR2_X1 U502 ( .A(n537), .B(n368), .ZN(n566) );
  XNOR2_X1 U503 ( .A(n536), .B(n369), .ZN(n368) );
  INV_X1 U504 ( .A(G475), .ZN(n369) );
  AND2_X1 U505 ( .A1(n561), .A2(n597), .ZN(n437) );
  XNOR2_X1 U506 ( .A(n489), .B(n366), .ZN(n727) );
  XNOR2_X1 U507 ( .A(n490), .B(n488), .ZN(n366) );
  XNOR2_X1 U508 ( .A(n520), .B(n431), .ZN(n430) );
  XNOR2_X1 U509 ( .A(n522), .B(n432), .ZN(n431) );
  XNOR2_X1 U510 ( .A(n657), .B(KEYINPUT79), .ZN(n658) );
  XNOR2_X1 U511 ( .A(n382), .B(n381), .ZN(n766) );
  INV_X1 U512 ( .A(KEYINPUT42), .ZN(n381) );
  INV_X1 U513 ( .A(KEYINPUT35), .ZN(n370) );
  INV_X1 U514 ( .A(KEYINPUT31), .ZN(n434) );
  NOR2_X1 U515 ( .A1(n564), .A2(n563), .ZN(n653) );
  NOR2_X1 U516 ( .A1(n729), .A2(n719), .ZN(n721) );
  INV_X1 U517 ( .A(n729), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n507), .B(n447), .ZN(n446) );
  INV_X1 U519 ( .A(n446), .ZN(n414) );
  XOR2_X1 U520 ( .A(n501), .B(n502), .Z(n355) );
  AND2_X1 U521 ( .A1(n419), .A2(n427), .ZN(n356) );
  XOR2_X1 U522 ( .A(n480), .B(G146), .Z(n357) );
  AND2_X1 U523 ( .A1(n399), .A2(n410), .ZN(n358) );
  AND2_X1 U524 ( .A1(n524), .A2(G210), .ZN(n359) );
  AND2_X1 U525 ( .A1(n560), .A2(n562), .ZN(n360) );
  OR2_X1 U526 ( .A1(n574), .A2(n511), .ZN(n361) );
  XNOR2_X1 U527 ( .A(G902), .B(KEYINPUT15), .ZN(n625) );
  INV_X1 U528 ( .A(KEYINPUT78), .ZN(n395) );
  XNOR2_X2 U529 ( .A(n362), .B(n571), .ZN(n448) );
  NAND2_X1 U530 ( .A1(n569), .A2(n570), .ZN(n362) );
  NOR2_X2 U531 ( .A1(n706), .A2(n729), .ZN(n707) );
  NAND2_X1 U532 ( .A1(n378), .A2(n624), .ZN(n394) );
  INV_X1 U533 ( .A(n557), .ZN(n436) );
  NAND2_X1 U534 ( .A1(n665), .A2(n666), .ZN(n557) );
  NAND2_X1 U535 ( .A1(n384), .A2(n614), .ZN(n375) );
  NOR2_X1 U536 ( .A1(n683), .A2(n648), .ZN(n377) );
  INV_X1 U537 ( .A(n662), .ZN(n577) );
  INV_X1 U538 ( .A(n558), .ZN(n428) );
  XNOR2_X1 U539 ( .A(n375), .B(n374), .ZN(n378) );
  NAND2_X1 U540 ( .A1(n651), .A2(n595), .ZN(n367) );
  XNOR2_X1 U541 ( .A(n538), .B(KEYINPUT98), .ZN(n429) );
  XNOR2_X1 U542 ( .A(n470), .B(n359), .ZN(n383) );
  XNOR2_X1 U543 ( .A(n383), .B(n475), .ZN(n629) );
  NAND2_X1 U544 ( .A1(n356), .A2(n420), .ZN(n371) );
  NAND2_X1 U545 ( .A1(n436), .A2(n669), .ZN(n674) );
  XNOR2_X1 U546 ( .A(n373), .B(n534), .ZN(n716) );
  XNOR2_X1 U547 ( .A(n533), .B(n535), .ZN(n373) );
  XNOR2_X1 U548 ( .A(n377), .B(n376), .ZN(n611) );
  NAND2_X1 U549 ( .A1(n676), .A2(n610), .ZN(n382) );
  OR2_X2 U550 ( .A1(n708), .A2(G902), .ZN(n458) );
  NOR2_X1 U551 ( .A1(n674), .A2(n558), .ZN(n435) );
  AND2_X1 U552 ( .A1(n387), .A2(n613), .ZN(n384) );
  XNOR2_X1 U553 ( .A(n453), .B(n452), .ZN(n451) );
  INV_X1 U554 ( .A(n761), .ZN(n387) );
  XNOR2_X2 U555 ( .A(G116), .B(KEYINPUT85), .ZN(n461) );
  NAND2_X1 U556 ( .A1(n391), .A2(n388), .ZN(n628) );
  AND2_X1 U557 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U558 ( .A1(n448), .A2(KEYINPUT78), .ZN(n390) );
  NOR2_X1 U559 ( .A1(n448), .A2(n393), .ZN(n392) );
  NAND2_X1 U560 ( .A1(n396), .A2(n409), .ZN(n408) );
  INV_X1 U561 ( .A(n510), .ZN(n404) );
  NOR2_X1 U562 ( .A1(n702), .A2(n413), .ZN(n412) );
  NAND2_X1 U563 ( .A1(n418), .A2(n427), .ZN(n417) );
  AND2_X1 U564 ( .A1(n437), .A2(n560), .ZN(n639) );
  NAND2_X1 U565 ( .A1(n654), .A2(KEYINPUT91), .ZN(n419) );
  INV_X1 U566 ( .A(n654), .ZN(n422) );
  NAND2_X1 U567 ( .A1(n437), .A2(n360), .ZN(n423) );
  NOR2_X1 U568 ( .A1(n654), .A2(n562), .ZN(n425) );
  INV_X1 U569 ( .A(n437), .ZN(n426) );
  INV_X1 U570 ( .A(n683), .ZN(n427) );
  XNOR2_X2 U571 ( .A(n435), .B(n434), .ZN(n654) );
  NOR2_X1 U572 ( .A1(n448), .A2(G953), .ZN(n736) );
  XNOR2_X2 U573 ( .A(n450), .B(KEYINPUT77), .ZN(n499) );
  XNOR2_X2 U574 ( .A(G143), .B(G128), .ZN(n450) );
  NAND2_X1 U575 ( .A1(n451), .A2(n603), .ZN(n548) );
  NAND2_X1 U576 ( .A1(n561), .A2(n687), .ZN(n453) );
  AND2_X1 U577 ( .A1(n456), .A2(n455), .ZN(G54) );
  XNOR2_X1 U578 ( .A(n457), .B(n712), .ZN(n456) );
  NAND2_X1 U579 ( .A1(n711), .A2(G469), .ZN(n457) );
  XNOR2_X2 U580 ( .A(n458), .B(G469), .ZN(n599) );
  XNOR2_X1 U581 ( .A(n659), .B(n658), .ZN(n661) );
  NOR2_X2 U582 ( .A1(n632), .A2(n729), .ZN(n635) );
  XNOR2_X1 U583 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U584 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U585 ( .A(KEYINPUT59), .B(KEYINPUT83), .ZN(n460) );
  INV_X1 U586 ( .A(KEYINPUT3), .ZN(n462) );
  INV_X1 U587 ( .A(n531), .ZN(n471) );
  XNOR2_X1 U588 ( .A(KEYINPUT30), .B(KEYINPUT103), .ZN(n586) );
  XNOR2_X1 U589 ( .A(n479), .B(n473), .ZN(n474) );
  XNOR2_X1 U590 ( .A(n495), .B(G122), .ZN(n496) );
  XNOR2_X1 U591 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U592 ( .A(n509), .B(KEYINPUT19), .ZN(n510) );
  XNOR2_X1 U593 ( .A(n629), .B(KEYINPUT62), .ZN(n630) );
  XNOR2_X1 U594 ( .A(n716), .B(n460), .ZN(n717) );
  XNOR2_X1 U595 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U596 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U597 ( .A1(G952), .A2(n755), .ZN(n729) );
  INV_X1 U598 ( .A(KEYINPUT45), .ZN(n571) );
  XNOR2_X1 U599 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U600 ( .A(n497), .B(n468), .Z(n470) );
  XOR2_X1 U601 ( .A(KEYINPUT75), .B(n469), .Z(n524) );
  XOR2_X1 U602 ( .A(KEYINPUT74), .B(KEYINPUT89), .Z(n473) );
  XNOR2_X1 U603 ( .A(n478), .B(n474), .ZN(n475) );
  NOR2_X1 U604 ( .A1(n629), .A2(G902), .ZN(n476) );
  XNOR2_X2 U605 ( .A(G472), .B(n476), .ZN(n597) );
  XOR2_X1 U606 ( .A(n597), .B(KEYINPUT6), .Z(n552) );
  NAND2_X1 U607 ( .A1(G227), .A2(n755), .ZN(n480) );
  XNOR2_X1 U608 ( .A(G119), .B(n482), .ZN(n490) );
  XOR2_X1 U609 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n484) );
  XNOR2_X1 U610 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U611 ( .A(n745), .B(n485), .ZN(n489) );
  NAND2_X1 U612 ( .A1(n755), .A2(G234), .ZN(n487) );
  XNOR2_X1 U613 ( .A(n487), .B(n486), .ZN(n519) );
  NAND2_X1 U614 ( .A1(n519), .A2(G221), .ZN(n488) );
  NAND2_X1 U615 ( .A1(G234), .A2(n625), .ZN(n491) );
  XNOR2_X1 U616 ( .A(KEYINPUT20), .B(n491), .ZN(n512) );
  NAND2_X1 U617 ( .A1(n512), .A2(G217), .ZN(n492) );
  NOR2_X1 U618 ( .A1(n545), .A2(n577), .ZN(n493) );
  NAND2_X1 U619 ( .A1(n552), .A2(n493), .ZN(n539) );
  XNOR2_X1 U620 ( .A(KEYINPUT14), .B(n494), .ZN(n693) );
  INV_X1 U621 ( .A(n625), .ZN(n505) );
  XOR2_X1 U622 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n495) );
  NAND2_X1 U623 ( .A1(G224), .A2(n755), .ZN(n502) );
  XNOR2_X1 U624 ( .A(n506), .B(KEYINPUT73), .ZN(n508) );
  NAND2_X1 U625 ( .A1(G210), .A2(n508), .ZN(n507) );
  NAND2_X1 U626 ( .A1(G214), .A2(n508), .ZN(n679) );
  INV_X1 U627 ( .A(G952), .ZN(n696) );
  NOR2_X1 U628 ( .A1(G953), .A2(n696), .ZN(n574) );
  NOR2_X1 U629 ( .A1(G898), .A2(n572), .ZN(n511) );
  NAND2_X1 U630 ( .A1(G221), .A2(n512), .ZN(n513) );
  XNOR2_X1 U631 ( .A(KEYINPUT21), .B(n513), .ZN(n663) );
  INV_X1 U632 ( .A(n514), .ZN(n518) );
  XNOR2_X1 U633 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U634 ( .A(n518), .B(n517), .ZN(n521) );
  NAND2_X1 U635 ( .A1(G217), .A2(n519), .ZN(n520) );
  XOR2_X1 U636 ( .A(n523), .B(G478), .Z(n565) );
  INV_X1 U637 ( .A(n565), .ZN(n563) );
  NAND2_X1 U638 ( .A1(G214), .A2(n524), .ZN(n535) );
  XNOR2_X1 U639 ( .A(n526), .B(n525), .ZN(n530) );
  XNOR2_X1 U640 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U641 ( .A(n530), .B(n529), .ZN(n534) );
  XNOR2_X1 U642 ( .A(n531), .B(KEYINPUT11), .ZN(n532) );
  XNOR2_X1 U643 ( .A(n745), .B(n532), .ZN(n533) );
  NOR2_X1 U644 ( .A1(G902), .A2(n716), .ZN(n537) );
  XNOR2_X1 U645 ( .A(KEYINPUT94), .B(KEYINPUT13), .ZN(n536) );
  NAND2_X1 U646 ( .A1(n563), .A2(n566), .ZN(n681) );
  NAND2_X1 U647 ( .A1(n545), .A2(n597), .ZN(n541) );
  NOR2_X1 U648 ( .A1(n553), .A2(n541), .ZN(n542) );
  NAND2_X1 U649 ( .A1(n662), .A2(n542), .ZN(n643) );
  NAND2_X1 U650 ( .A1(n765), .A2(n643), .ZN(n544) );
  NOR2_X1 U651 ( .A1(KEYINPUT44), .A2(KEYINPUT81), .ZN(n543) );
  XNOR2_X1 U652 ( .A(n544), .B(n543), .ZN(n549) );
  NOR2_X1 U653 ( .A1(n557), .A2(n552), .ZN(n546) );
  INV_X1 U654 ( .A(n566), .ZN(n564) );
  NAND2_X1 U655 ( .A1(n564), .A2(n565), .ZN(n547) );
  XNOR2_X1 U656 ( .A(n547), .B(KEYINPUT101), .ZN(n603) );
  NAND2_X1 U657 ( .A1(n549), .A2(n759), .ZN(n551) );
  NAND2_X1 U658 ( .A1(n551), .A2(n550), .ZN(n570) );
  INV_X1 U659 ( .A(n552), .ZN(n578) );
  NOR2_X1 U660 ( .A1(n578), .A2(n553), .ZN(n555) );
  NOR2_X1 U661 ( .A1(n662), .A2(n372), .ZN(n554) );
  NAND2_X1 U662 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U663 ( .A(KEYINPUT99), .B(n556), .ZN(n760) );
  INV_X1 U664 ( .A(KEYINPUT91), .ZN(n562) );
  INV_X1 U665 ( .A(n597), .ZN(n669) );
  NAND2_X1 U666 ( .A1(n599), .A2(n666), .ZN(n559) );
  INV_X1 U667 ( .A(n589), .ZN(n560) );
  XOR2_X1 U668 ( .A(KEYINPUT97), .B(n653), .Z(n616) );
  NOR2_X1 U669 ( .A1(n566), .A2(n565), .ZN(n651) );
  NOR2_X1 U670 ( .A1(n616), .A2(n651), .ZN(n683) );
  XNOR2_X1 U671 ( .A(n568), .B(KEYINPUT100), .ZN(n569) );
  NOR2_X1 U672 ( .A1(G900), .A2(n572), .ZN(n573) );
  NOR2_X1 U673 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U674 ( .A(n693), .ZN(n575) );
  NOR2_X1 U675 ( .A1(n576), .A2(n575), .ZN(n595) );
  INV_X1 U676 ( .A(n651), .ZN(n649) );
  NOR2_X1 U677 ( .A1(n577), .A2(n663), .ZN(n594) );
  AND2_X1 U678 ( .A1(n594), .A2(n578), .ZN(n579) );
  NAND2_X1 U679 ( .A1(n579), .A2(n679), .ZN(n580) );
  XNOR2_X1 U680 ( .A(KEYINPUT36), .B(KEYINPUT82), .ZN(n581) );
  XNOR2_X1 U681 ( .A(n582), .B(n581), .ZN(n583) );
  NAND2_X1 U682 ( .A1(n372), .A2(n583), .ZN(n584) );
  NAND2_X1 U683 ( .A1(n669), .A2(n679), .ZN(n587) );
  NAND2_X1 U684 ( .A1(n678), .A2(n604), .ZN(n590) );
  NAND2_X1 U685 ( .A1(n678), .A2(n679), .ZN(n592) );
  NAND2_X1 U686 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U687 ( .A(KEYINPUT28), .B(n598), .Z(n601) );
  XNOR2_X1 U688 ( .A(n599), .B(KEYINPUT105), .ZN(n600) );
  NOR2_X1 U689 ( .A1(n601), .A2(n600), .ZN(n610) );
  XNOR2_X1 U690 ( .A(n602), .B(KEYINPUT46), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n603), .A2(n621), .ZN(n606) );
  INV_X1 U692 ( .A(n604), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U694 ( .A(n607), .B(KEYINPUT104), .ZN(n769) );
  INV_X1 U695 ( .A(n608), .ZN(n609) );
  NAND2_X1 U696 ( .A1(n610), .A2(n609), .ZN(n648) );
  XNOR2_X1 U697 ( .A(KEYINPUT72), .B(n612), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n617), .B(KEYINPUT108), .ZN(n768) );
  NOR2_X1 U700 ( .A1(n372), .A2(n618), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n619), .B(KEYINPUT43), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U703 ( .A(KEYINPUT102), .B(n622), .ZN(n763) );
  INV_X1 U704 ( .A(n763), .ZN(n623) );
  XOR2_X1 U705 ( .A(KEYINPUT80), .B(n625), .Z(n626) );
  NAND2_X1 U706 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U707 ( .A1(KEYINPUT2), .A2(n659), .ZN(n713) );
  NAND2_X1 U708 ( .A1(n711), .A2(G472), .ZN(n631) );
  XNOR2_X1 U709 ( .A(KEYINPUT84), .B(KEYINPUT109), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(KEYINPUT63), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n635), .B(n634), .ZN(G57) );
  XOR2_X1 U712 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n637) );
  NAND2_X1 U713 ( .A1(n639), .A2(n651), .ZN(n636) );
  XNOR2_X1 U714 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U715 ( .A(G104), .B(n638), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n641) );
  NAND2_X1 U717 ( .A1(n639), .A2(n653), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U719 ( .A(G107), .B(n642), .ZN(G9) );
  XNOR2_X1 U720 ( .A(G110), .B(KEYINPUT112), .ZN(n644) );
  XNOR2_X1 U721 ( .A(n644), .B(n643), .ZN(G12) );
  INV_X1 U722 ( .A(n653), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n645), .A2(n648), .ZN(n647) );
  XNOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .ZN(n646) );
  XNOR2_X1 U725 ( .A(n647), .B(n646), .ZN(G30) );
  NOR2_X1 U726 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U727 ( .A(G146), .B(n650), .Z(G48) );
  NAND2_X1 U728 ( .A1(n354), .A2(n651), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n652), .B(G113), .ZN(G15) );
  NAND2_X1 U730 ( .A1(n354), .A2(n653), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n655), .B(KEYINPUT114), .ZN(n656) );
  XNOR2_X1 U732 ( .A(G116), .B(n656), .ZN(G18) );
  INV_X1 U733 ( .A(KEYINPUT2), .ZN(n657) );
  NAND2_X1 U734 ( .A1(n687), .A2(n676), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n698) );
  AND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U737 ( .A(KEYINPUT49), .B(n664), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n666), .A2(n372), .ZN(n668) );
  XNOR2_X1 U739 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(n670) );
  NOR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U744 ( .A(KEYINPUT51), .B(n675), .Z(n677) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n690) );
  NOR2_X1 U746 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n685) );
  NOR2_X1 U748 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U750 ( .A(KEYINPUT117), .B(n686), .ZN(n688) );
  NAND2_X1 U751 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U752 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U753 ( .A(n691), .B(KEYINPUT52), .ZN(n692) );
  XNOR2_X1 U754 ( .A(KEYINPUT118), .B(n692), .ZN(n694) );
  NAND2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U757 ( .A(n699), .B(KEYINPUT119), .ZN(n700) );
  NOR2_X1 U758 ( .A1(G953), .A2(n700), .ZN(n701) );
  XNOR2_X1 U759 ( .A(KEYINPUT53), .B(n701), .ZN(G75) );
  NAND2_X1 U760 ( .A1(n711), .A2(G210), .ZN(n705) );
  XOR2_X1 U761 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n703) );
  XNOR2_X1 U762 ( .A(n707), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U763 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n708), .B(KEYINPUT57), .ZN(n709) );
  XNOR2_X1 U765 ( .A(n710), .B(n709), .ZN(n712) );
  AND2_X1 U766 ( .A1(G475), .A2(n713), .ZN(n714) );
  NAND2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n718) );
  XNOR2_X1 U768 ( .A(KEYINPUT64), .B(KEYINPUT60), .ZN(n720) );
  XNOR2_X1 U769 ( .A(n721), .B(n720), .ZN(G60) );
  XOR2_X1 U770 ( .A(n722), .B(KEYINPUT121), .Z(n724) );
  NAND2_X1 U771 ( .A1(n711), .A2(G478), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U773 ( .A1(n729), .A2(n725), .ZN(G63) );
  NAND2_X1 U774 ( .A1(G217), .A2(n711), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U776 ( .A1(n729), .A2(n728), .ZN(G66) );
  XNOR2_X1 U777 ( .A(n730), .B(KEYINPUT123), .ZN(n732) );
  XNOR2_X1 U778 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(G101), .ZN(n735) );
  NOR2_X1 U780 ( .A1(n755), .A2(G898), .ZN(n734) );
  NOR2_X1 U781 ( .A1(n735), .A2(n734), .ZN(n742) );
  XOR2_X1 U782 ( .A(KEYINPUT122), .B(n736), .Z(n740) );
  NAND2_X1 U783 ( .A1(G953), .A2(G224), .ZN(n737) );
  XNOR2_X1 U784 ( .A(KEYINPUT61), .B(n737), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n738), .A2(G898), .ZN(n739) );
  NAND2_X1 U786 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U787 ( .A(n742), .B(n741), .ZN(G69) );
  XOR2_X1 U788 ( .A(n743), .B(KEYINPUT124), .Z(n744) );
  XNOR2_X1 U789 ( .A(n745), .B(n744), .ZN(n746) );
  XOR2_X1 U790 ( .A(n747), .B(n746), .Z(n751) );
  INV_X1 U791 ( .A(n751), .ZN(n748) );
  XOR2_X1 U792 ( .A(n748), .B(n394), .Z(n749) );
  NOR2_X1 U793 ( .A1(G953), .A2(n749), .ZN(n750) );
  XNOR2_X1 U794 ( .A(KEYINPUT125), .B(n750), .ZN(n758) );
  XOR2_X1 U795 ( .A(G227), .B(n751), .Z(n752) );
  NAND2_X1 U796 ( .A1(n752), .A2(G900), .ZN(n753) );
  XOR2_X1 U797 ( .A(KEYINPUT126), .B(n753), .Z(n754) );
  NOR2_X1 U798 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U799 ( .A(KEYINPUT127), .B(n756), .ZN(n757) );
  NAND2_X1 U800 ( .A1(n758), .A2(n757), .ZN(G72) );
  XNOR2_X1 U801 ( .A(G122), .B(n759), .ZN(G24) );
  XOR2_X1 U802 ( .A(G101), .B(n760), .Z(G3) );
  XNOR2_X1 U803 ( .A(n761), .B(G125), .ZN(n762) );
  XNOR2_X1 U804 ( .A(n762), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U805 ( .A(G140), .B(KEYINPUT115), .ZN(n764) );
  XNOR2_X1 U806 ( .A(n764), .B(n763), .ZN(G42) );
  XNOR2_X1 U807 ( .A(n765), .B(G119), .ZN(G21) );
  XOR2_X1 U808 ( .A(n766), .B(G137), .Z(G39) );
  XOR2_X1 U809 ( .A(G131), .B(n767), .Z(G33) );
  XNOR2_X1 U810 ( .A(G134), .B(n768), .ZN(G36) );
  XNOR2_X1 U811 ( .A(G143), .B(KEYINPUT113), .ZN(n770) );
  XNOR2_X1 U812 ( .A(n770), .B(n769), .ZN(G45) );
endmodule

