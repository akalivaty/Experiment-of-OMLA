

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(n452), .B(n451), .ZN(n518) );
  XNOR2_X1 U325 ( .A(n395), .B(n312), .ZN(n533) );
  XOR2_X1 U326 ( .A(KEYINPUT93), .B(n425), .Z(n531) );
  XNOR2_X1 U327 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U328 ( .A(n403), .B(n317), .ZN(n318) );
  XNOR2_X1 U329 ( .A(n407), .B(n406), .ZN(n410) );
  XNOR2_X1 U330 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U331 ( .A(n450), .B(KEYINPUT37), .ZN(n451) );
  INV_X1 U332 ( .A(KEYINPUT108), .ZN(n453) );
  XNOR2_X1 U333 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U334 ( .A(n453), .B(KEYINPUT38), .ZN(n454) );
  XNOR2_X1 U335 ( .A(n329), .B(n328), .ZN(n578) );
  NOR2_X1 U336 ( .A1(n533), .A2(n475), .ZN(n568) );
  XOR2_X1 U337 ( .A(n473), .B(KEYINPUT28), .Z(n526) );
  XNOR2_X1 U338 ( .A(n455), .B(n454), .ZN(n503) );
  XNOR2_X1 U339 ( .A(n476), .B(G190GAT), .ZN(n477) );
  XNOR2_X1 U340 ( .A(n456), .B(G43GAT), .ZN(n457) );
  XNOR2_X1 U341 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U344 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n292) );
  XNOR2_X1 U345 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(n294), .ZN(n395) );
  XOR2_X1 U347 ( .A(KEYINPUT82), .B(KEYINPUT64), .Z(n296) );
  XNOR2_X1 U348 ( .A(G15GAT), .B(G120GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U350 ( .A(G183GAT), .B(KEYINPUT85), .Z(n298) );
  XNOR2_X1 U351 ( .A(KEYINPUT83), .B(KEYINPUT20), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(n300), .B(n299), .Z(n311) );
  XOR2_X1 U354 ( .A(G127GAT), .B(G176GAT), .Z(n302) );
  XNOR2_X1 U355 ( .A(G71GAT), .B(KEYINPUT86), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n309) );
  XOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT0), .Z(n371) );
  XOR2_X1 U358 ( .A(G190GAT), .B(G99GAT), .Z(n304) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U361 ( .A(n371), .B(n305), .Z(n307) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U364 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U366 ( .A(G71GAT), .B(G57GAT), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n313), .B(KEYINPUT13), .ZN(n354) );
  XOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .Z(n439) );
  XOR2_X1 U369 ( .A(n354), .B(n439), .Z(n321) );
  XOR2_X1 U370 ( .A(G64GAT), .B(G92GAT), .Z(n315) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n388) );
  INV_X1 U373 ( .A(KEYINPUT33), .ZN(n316) );
  XNOR2_X1 U374 ( .A(n388), .B(n316), .ZN(n319) );
  XOR2_X1 U375 ( .A(G106GAT), .B(G78GAT), .Z(n403) );
  NAND2_X1 U376 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U377 ( .A(n321), .B(n320), .ZN(n323) );
  INV_X1 U378 ( .A(KEYINPUT32), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n329) );
  XOR2_X1 U380 ( .A(G120GAT), .B(G148GAT), .Z(n365) );
  XNOR2_X1 U381 ( .A(n365), .B(KEYINPUT73), .ZN(n327) );
  XOR2_X1 U382 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n325) );
  XNOR2_X1 U383 ( .A(KEYINPUT72), .B(KEYINPUT74), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  INV_X1 U385 ( .A(n578), .ZN(n465) );
  XOR2_X1 U386 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n331) );
  XNOR2_X1 U387 ( .A(G8GAT), .B(G1GAT), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n348) );
  XOR2_X1 U389 ( .A(G197GAT), .B(G141GAT), .Z(n333) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G113GAT), .ZN(n332) );
  XNOR2_X1 U391 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U392 ( .A(G29GAT), .B(G36GAT), .Z(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n344) );
  XNOR2_X1 U394 ( .A(KEYINPUT66), .B(KEYINPUT29), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n336), .B(KEYINPUT67), .ZN(n337) );
  XOR2_X1 U396 ( .A(n337), .B(KEYINPUT30), .Z(n342) );
  XOR2_X1 U397 ( .A(G43GAT), .B(G50GAT), .Z(n339) );
  XNOR2_X1 U398 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n435) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(G22GAT), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n340), .B(KEYINPUT69), .ZN(n356) );
  XNOR2_X1 U402 ( .A(n435), .B(n356), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n346) );
  NAND2_X1 U405 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U406 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U407 ( .A(n348), .B(n347), .Z(n535) );
  INV_X1 U408 ( .A(n535), .ZN(n573) );
  NAND2_X1 U409 ( .A1(n465), .A2(n573), .ZN(n490) );
  XOR2_X1 U410 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n350) );
  XNOR2_X1 U411 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n364) );
  XNOR2_X1 U413 ( .A(G1GAT), .B(G127GAT), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n351), .B(G155GAT), .ZN(n366) );
  XOR2_X1 U415 ( .A(G64GAT), .B(n366), .Z(n353) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n355) );
  XOR2_X1 U418 ( .A(n355), .B(n354), .Z(n358) );
  XNOR2_X1 U419 ( .A(n356), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U421 ( .A(n359), .B(KEYINPUT12), .Z(n362) );
  XNOR2_X1 U422 ( .A(G8GAT), .B(G183GAT), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n360), .B(G211GAT), .ZN(n392) );
  XNOR2_X1 U424 ( .A(n392), .B(KEYINPUT79), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n581) );
  XOR2_X1 U427 ( .A(n366), .B(n365), .Z(n373) );
  XNOR2_X1 U428 ( .A(G29GAT), .B(G134GAT), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n367), .B(KEYINPUT77), .ZN(n434) );
  XOR2_X1 U430 ( .A(KEYINPUT4), .B(n434), .Z(n369) );
  NAND2_X1 U431 ( .A1(G225GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U435 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n375) );
  XNOR2_X1 U436 ( .A(G85GAT), .B(G57GAT), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U438 ( .A(n377), .B(n376), .Z(n385) );
  XOR2_X1 U439 ( .A(KEYINPUT2), .B(G162GAT), .Z(n379) );
  XNOR2_X1 U440 ( .A(KEYINPUT88), .B(KEYINPUT3), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U442 ( .A(G141GAT), .B(n380), .Z(n414) );
  XOR2_X1 U443 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n382) );
  XNOR2_X1 U444 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n414), .B(n383), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n425) );
  XOR2_X1 U448 ( .A(G36GAT), .B(G190GAT), .Z(n438) );
  XOR2_X1 U449 ( .A(KEYINPUT94), .B(n438), .Z(n387) );
  NAND2_X1 U450 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U451 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U452 ( .A(n389), .B(n388), .Z(n394) );
  XOR2_X1 U453 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n391) );
  XNOR2_X1 U454 ( .A(G197GAT), .B(G218GAT), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n408) );
  XNOR2_X1 U456 ( .A(n408), .B(n392), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n521) );
  XNOR2_X1 U459 ( .A(n521), .B(KEYINPUT95), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n397), .B(KEYINPUT27), .ZN(n422) );
  XOR2_X1 U461 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n399) );
  XNOR2_X1 U462 ( .A(G22GAT), .B(G148GAT), .ZN(n398) );
  XOR2_X1 U463 ( .A(n399), .B(n398), .Z(n412) );
  XOR2_X1 U464 ( .A(G155GAT), .B(G211GAT), .Z(n401) );
  XNOR2_X1 U465 ( .A(G50GAT), .B(KEYINPUT24), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n403), .B(n402), .ZN(n407) );
  AND2_X1 U468 ( .A1(G228GAT), .A2(G233GAT), .ZN(n405) );
  INV_X1 U469 ( .A(G204GAT), .ZN(n404) );
  XNOR2_X1 U470 ( .A(n408), .B(KEYINPUT22), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U472 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U473 ( .A(n414), .B(n413), .Z(n473) );
  NAND2_X1 U474 ( .A1(n422), .A2(n526), .ZN(n532) );
  NOR2_X1 U475 ( .A1(n531), .A2(n532), .ZN(n415) );
  AND2_X1 U476 ( .A1(n533), .A2(n415), .ZN(n417) );
  INV_X1 U477 ( .A(KEYINPUT96), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n428) );
  NOR2_X1 U479 ( .A1(n533), .A2(n521), .ZN(n418) );
  NOR2_X1 U480 ( .A1(n473), .A2(n418), .ZN(n419) );
  XNOR2_X1 U481 ( .A(KEYINPUT25), .B(n419), .ZN(n424) );
  XOR2_X1 U482 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n421) );
  NAND2_X1 U483 ( .A1(n473), .A2(n533), .ZN(n420) );
  XNOR2_X1 U484 ( .A(n421), .B(n420), .ZN(n572) );
  INV_X1 U485 ( .A(n572), .ZN(n423) );
  NAND2_X1 U486 ( .A1(n423), .A2(n422), .ZN(n551) );
  NAND2_X1 U487 ( .A1(n424), .A2(n551), .ZN(n426) );
  NAND2_X1 U488 ( .A1(n426), .A2(n425), .ZN(n427) );
  NAND2_X1 U489 ( .A1(n428), .A2(n427), .ZN(n487) );
  XOR2_X1 U490 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n430) );
  XNOR2_X1 U491 ( .A(KEYINPUT78), .B(KEYINPUT10), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n447) );
  XOR2_X1 U493 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n432) );
  NAND2_X1 U494 ( .A1(G232GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U496 ( .A(n433), .B(KEYINPUT76), .Z(n437) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U499 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U500 ( .A(G106GAT), .B(G92GAT), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U502 ( .A(n443), .B(n442), .Z(n445) );
  XNOR2_X1 U503 ( .A(G162GAT), .B(G218GAT), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n485) );
  INV_X1 U506 ( .A(n485), .ZN(n557) );
  XNOR2_X1 U507 ( .A(n557), .B(KEYINPUT106), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n448), .B(KEYINPUT36), .ZN(n583) );
  NAND2_X1 U509 ( .A1(n487), .A2(n583), .ZN(n449) );
  NOR2_X1 U510 ( .A1(n581), .A2(n449), .ZN(n452) );
  INV_X1 U511 ( .A(KEYINPUT107), .ZN(n450) );
  NOR2_X1 U512 ( .A1(n490), .A2(n518), .ZN(n455) );
  NOR2_X1 U513 ( .A1(n533), .A2(n503), .ZN(n458) );
  XNOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n456) );
  XOR2_X1 U515 ( .A(KEYINPUT41), .B(n578), .Z(n565) );
  AND2_X1 U516 ( .A1(n565), .A2(n573), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT46), .ZN(n460) );
  XOR2_X1 U518 ( .A(n581), .B(KEYINPUT117), .Z(n569) );
  NOR2_X1 U519 ( .A1(n460), .A2(n569), .ZN(n461) );
  NAND2_X1 U520 ( .A1(n461), .A2(n485), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT47), .ZN(n469) );
  NAND2_X1 U522 ( .A1(n583), .A2(n581), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT45), .B(KEYINPUT118), .Z(n463) );
  XNOR2_X1 U524 ( .A(n464), .B(n463), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n573), .A2(n467), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT48), .ZN(n530) );
  NOR2_X1 U529 ( .A1(n521), .A2(n530), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT54), .B(n471), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n472), .A2(n531), .ZN(n571) );
  NOR2_X1 U532 ( .A1(n473), .A2(n571), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n474), .B(KEYINPUT55), .ZN(n475) );
  NAND2_X1 U534 ( .A1(n568), .A2(n557), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n476) );
  INV_X1 U536 ( .A(G29GAT), .ZN(n482) );
  NOR2_X1 U537 ( .A1(n503), .A2(n531), .ZN(n480) );
  XNOR2_X1 U538 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(G1328GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n484) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n493) );
  AND2_X1 U544 ( .A1(n485), .A2(n581), .ZN(n486) );
  XNOR2_X1 U545 ( .A(KEYINPUT16), .B(n486), .ZN(n488) );
  NAND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(KEYINPUT98), .ZN(n505) );
  NOR2_X1 U548 ( .A1(n490), .A2(n505), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n491), .B(KEYINPUT99), .ZN(n499) );
  NOR2_X1 U550 ( .A1(n531), .A2(n499), .ZN(n492) );
  XOR2_X1 U551 ( .A(n493), .B(n492), .Z(G1324GAT) );
  NOR2_X1 U552 ( .A1(n521), .A2(n499), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT102), .B(n494), .Z(n495) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n495), .ZN(G1325GAT) );
  NOR2_X1 U555 ( .A1(n533), .A2(n499), .ZN(n497) );
  XNOR2_X1 U556 ( .A(KEYINPUT103), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n498), .Z(G1326GAT) );
  NOR2_X1 U559 ( .A1(n526), .A2(n499), .ZN(n500) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(n500), .Z(n501) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n501), .ZN(G1327GAT) );
  NOR2_X1 U562 ( .A1(n521), .A2(n503), .ZN(n502) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U564 ( .A1(n526), .A2(n503), .ZN(n504) );
  XOR2_X1 U565 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  NAND2_X1 U566 ( .A1(n535), .A2(n565), .ZN(n517) );
  OR2_X1 U567 ( .A1(n505), .A2(n517), .ZN(n512) );
  NOR2_X1 U568 ( .A1(n531), .A2(n512), .ZN(n507) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NOR2_X1 U572 ( .A1(n521), .A2(n512), .ZN(n509) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n509), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n533), .A2(n512), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n526), .ZN(n516) );
  XOR2_X1 U578 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n514) );
  XNOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U583 ( .A(KEYINPUT114), .B(n519), .Z(n525) );
  NOR2_X1 U584 ( .A1(n531), .A2(n525), .ZN(n520) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n520), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n521), .A2(n525), .ZN(n522) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n522), .Z(G1337GAT) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n524) );
  NOR2_X1 U589 ( .A1(n533), .A2(n525), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  XNOR2_X1 U591 ( .A(KEYINPUT116), .B(KEYINPUT44), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n549) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n549), .A2(n534), .ZN(n542) );
  NOR2_X1 U598 ( .A1(n535), .A2(n542), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(KEYINPUT119), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  INV_X1 U601 ( .A(n565), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n538), .A2(n542), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT120), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n544) );
  INV_X1 U607 ( .A(n542), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n546), .A2(n569), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U612 ( .A1(n546), .A2(n557), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  INV_X1 U614 ( .A(n549), .ZN(n550) );
  NOR2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n558), .A2(n573), .ZN(n552) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U619 ( .A1(n558), .A2(n565), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n581), .A2(n558), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n568), .A2(n573), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n563) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(n564), .Z(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n565), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n584) );
  NAND2_X1 U638 ( .A1(n573), .A2(n584), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

