//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n541, new_n542, new_n543,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g023(.A(G2106), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n453), .A2(new_n449), .B1(new_n457), .B2(new_n454), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n461), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n461), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OAI21_X1  g053(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NOR3_X1   g055(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G112), .B2(new_n461), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n476), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT70), .Z(G162));
  NAND4_X1  g059(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n461), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT72), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT72), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n473), .A2(new_n487), .A3(G138), .A4(new_n461), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(KEYINPUT71), .A2(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT71), .A2(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n461), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n485), .A2(KEYINPUT72), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n506), .A2(new_n512), .ZN(G166));
  AOI22_X1  g088(.A1(new_n507), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(new_n503), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n510), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  OR3_X1    g096(.A1(new_n516), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n516), .B2(new_n520), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(G168));
  AOI22_X1  g099(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n505), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  INV_X1    g102(.A(G52), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n508), .A2(new_n527), .B1(new_n510), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G171));
  AOI22_X1  g105(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n505), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G81), .ZN(new_n534));
  INV_X1    g109(.A(G43), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n508), .A2(new_n534), .B1(new_n510), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  AND3_X1   g113(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G36), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT74), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(G188));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n507), .A2(G53), .A3(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n548), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT76), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n551), .B1(new_n546), .B2(KEYINPUT9), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n546), .A2(KEYINPUT75), .A3(KEYINPUT9), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n549), .A2(new_n550), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n515), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n508), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(G651), .B1(new_n558), .B2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n554), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND2_X1  g138(.A1(new_n558), .A2(G87), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n507), .A2(G543), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(G288));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n508), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n565), .A2(G48), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n501), .B2(new_n502), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n503), .A2(new_n507), .A3(KEYINPUT78), .A4(G86), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n571), .A2(new_n572), .A3(new_n578), .A4(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n505), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  INV_X1    g158(.A(G47), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n508), .A2(new_n583), .B1(new_n510), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT79), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n503), .A2(new_n507), .A3(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n515), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G54), .B2(new_n565), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT80), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n589), .B1(new_n597), .B2(G868), .ZN(G321));
  NOR2_X1   g174(.A1(G299), .A2(G868), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g176(.A(new_n600), .B1(G868), .B2(G168), .ZN(G280));
  XNOR2_X1  g177(.A(KEYINPUT81), .B(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n597), .B1(G860), .B2(new_n603), .ZN(G148));
  INV_X1    g179(.A(new_n537), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n597), .A2(new_n603), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT82), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n606), .B1(new_n608), .B2(G868), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n475), .A2(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n475), .A2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n477), .A2(G123), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2443), .B(G2446), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT83), .ZN(new_n638));
  OAI21_X1  g213(.A(G14), .B1(new_n634), .B2(new_n636), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n646), .A2(KEYINPUT84), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(KEYINPUT84), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(KEYINPUT17), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n647), .B(new_n648), .C1(new_n643), .C2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n644), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n651), .A2(new_n642), .A3(new_n641), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n643), .A3(new_n641), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  AOI211_X1 g242(.A(new_n665), .B(new_n667), .C1(new_n660), .C2(new_n664), .ZN(new_n668));
  XOR2_X1   g243(.A(G1981), .B(G1986), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n586), .A2(G16), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G16), .B2(G24), .ZN(new_n678));
  INV_X1    g253(.A(G1986), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n475), .A2(G131), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n477), .A2(G119), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n461), .A2(G107), .ZN(new_n683));
  OAI21_X1  g258(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  MUX2_X1   g260(.A(G25), .B(new_n685), .S(G29), .Z(new_n686));
  XOR2_X1   g261(.A(KEYINPUT35), .B(G1991), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  AOI211_X1 g264(.A(new_n680), .B(new_n689), .C1(new_n679), .C2(new_n678), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G23), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n691), .A2(G6), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G305), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G16), .A2(G22), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G166), .B2(G16), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT88), .B(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n698), .B2(new_n700), .ZN(new_n707));
  OAI21_X1  g282(.A(KEYINPUT34), .B1(new_n702), .B2(new_n707), .ZN(new_n708));
  OR3_X1    g283(.A1(new_n702), .A2(new_n707), .A3(KEYINPUT34), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n690), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT36), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G35), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT98), .Z(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G162), .B2(new_n712), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT29), .B(G2090), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G29), .A2(G32), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n475), .A2(G141), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n477), .A2(G129), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT26), .Z(new_n723));
  NAND4_X1  g298(.A1(new_n719), .A2(new_n720), .A3(new_n721), .A4(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  AOI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(G29), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT27), .B(G1996), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2078), .ZN(new_n729));
  NOR2_X1   g304(.A1(G164), .A2(new_n712), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G27), .B2(new_n712), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n717), .B(new_n728), .C1(new_n729), .C2(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT92), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n712), .A2(G26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n475), .A2(G140), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT90), .Z(new_n738));
  OR2_X1    g313(.A1(new_n461), .A2(G116), .ZN(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n477), .A2(G128), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n736), .B1(new_n743), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2067), .ZN(new_n745));
  NOR2_X1   g320(.A1(G171), .A2(new_n691), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G5), .B2(new_n691), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n712), .A2(G33), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT93), .B(KEYINPUT25), .Z(new_n751));
  NAND3_X1  g326(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n475), .A2(G139), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n753), .B(new_n754), .C1(new_n461), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(G29), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n747), .A2(new_n748), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G16), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n537), .B2(G16), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G1341), .ZN(new_n761));
  INV_X1    g336(.A(G34), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n712), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G160), .B2(new_n712), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n761), .B1(G2084), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n745), .A2(new_n758), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n747), .A2(new_n748), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT97), .Z(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G21), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G168), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n729), .B2(new_n731), .ZN(new_n775));
  INV_X1    g350(.A(new_n757), .ZN(new_n776));
  AOI22_X1  g351(.A1(G2072), .A2(new_n776), .B1(new_n760), .B2(G1341), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n621), .A2(new_n712), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT31), .B(G11), .Z(new_n779));
  INV_X1    g354(.A(G28), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(KEYINPUT30), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n781), .A2(KEYINPUT96), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(KEYINPUT96), .ZN(new_n783));
  OR3_X1    g358(.A1(new_n780), .A2(KEYINPUT95), .A3(KEYINPUT30), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT95), .B1(new_n780), .B2(KEYINPUT30), .ZN(new_n785));
  AND4_X1   g360(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n778), .A2(new_n779), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n777), .B(new_n787), .C1(G2084), .C2(new_n766), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n768), .A2(new_n770), .A3(new_n775), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n691), .A2(G4), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n597), .B2(new_n691), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1348), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n691), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT23), .Z(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G299), .B2(G16), .ZN(new_n795));
  INV_X1    g370(.A(G1956), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n711), .A2(new_n732), .A3(new_n789), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n710), .A2(KEYINPUT36), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(G311));
  XNOR2_X1  g376(.A(G311), .B(KEYINPUT99), .ZN(G150));
  AOI22_X1  g377(.A1(new_n558), .A2(G93), .B1(new_n565), .B2(G55), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(new_n505), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n537), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(KEYINPUT100), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n605), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n597), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n813), .A2(new_n814), .A3(G860), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n808), .A2(G860), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT37), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n815), .A2(new_n817), .ZN(G145));
  XOR2_X1   g393(.A(new_n612), .B(new_n685), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n477), .A2(G130), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT102), .ZN(new_n821));
  INV_X1    g396(.A(G118), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n822), .A2(KEYINPUT103), .A3(G2105), .ZN(new_n823));
  AOI21_X1  g398(.A(KEYINPUT103), .B1(new_n822), .B2(G2105), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n475), .A2(G142), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n821), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n819), .B(new_n828), .Z(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT104), .Z(new_n830));
  MUX2_X1   g405(.A(new_n725), .B(new_n724), .S(new_n756), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n743), .B(G164), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(G162), .B(G160), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(new_n621), .Z(new_n837));
  INV_X1    g412(.A(new_n829), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  OR3_X1    g414(.A1(new_n834), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G37), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n830), .A2(new_n833), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n837), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g420(.A(new_n586), .B(G288), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT107), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(G166), .B(G305), .Z(new_n850));
  OR2_X1    g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n847), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(new_n852), .A3(new_n850), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n855));
  INV_X1    g430(.A(new_n596), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G299), .ZN(new_n857));
  MUX2_X1   g432(.A(new_n855), .B(KEYINPUT41), .S(new_n857), .Z(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n608), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n860), .A2(new_n809), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n809), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT106), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n608), .B(new_n809), .Z(new_n865));
  INV_X1    g440(.A(new_n857), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n863), .A2(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT106), .B1(new_n865), .B2(new_n859), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n854), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n865), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n863), .A2(new_n864), .ZN(new_n871));
  INV_X1    g446(.A(new_n854), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n865), .A2(KEYINPUT106), .A3(new_n859), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n870), .A2(new_n871), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n875));
  AND3_X1   g450(.A1(new_n869), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n875), .B1(new_n869), .B2(new_n874), .ZN(new_n877));
  OAI21_X1  g452(.A(G868), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G868), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n808), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(G295));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n880), .ZN(G331));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n883));
  XNOR2_X1  g458(.A(G168), .B(G171), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n809), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n857), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n858), .B2(new_n885), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n887), .A2(new_n872), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n872), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n841), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n866), .A2(new_n855), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(KEYINPUT41), .B2(new_n857), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n872), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n841), .A4(new_n888), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n883), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI211_X1 g476(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n891), .C2(new_n898), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n896), .A2(new_n841), .A3(new_n888), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT44), .B1(new_n904), .B2(new_n897), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n901), .A2(new_n902), .B1(new_n903), .B2(new_n905), .ZN(G397));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n907));
  INV_X1    g482(.A(G1384), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT45), .B1(new_n499), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(G160), .A2(G40), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n486), .A2(new_n488), .A3(KEYINPUT4), .ZN(new_n912));
  AND2_X1   g487(.A1(KEYINPUT71), .A2(G114), .ZN(new_n913));
  NOR2_X1   g488(.A1(KEYINPUT71), .A2(G114), .ZN(new_n914));
  OAI21_X1  g489(.A(G2105), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n494), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n498), .A2(new_n490), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n908), .B1(new_n912), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G40), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n468), .A2(new_n471), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(KEYINPUT112), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n908), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n911), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n773), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT113), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(KEYINPUT113), .A3(new_n773), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n919), .A2(KEYINPUT50), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n499), .A2(new_n932), .A3(new_n908), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n923), .A3(new_n933), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(G2084), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n929), .A2(G168), .A3(new_n930), .A4(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G8), .ZN(new_n937));
  NAND2_X1  g512(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT119), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT51), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n936), .A2(new_n939), .A3(new_n940), .A4(G8), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(G8), .A3(G286), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n947));
  INV_X1    g522(.A(G2090), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n931), .A2(new_n948), .A3(new_n923), .A4(new_n933), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n910), .B1(new_n919), .B2(new_n920), .ZN(new_n951));
  AOI21_X1  g526(.A(G1971), .B1(new_n951), .B2(new_n925), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1971), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n485), .A2(KEYINPUT72), .A3(new_n497), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n495), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n956), .B2(new_n489), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n923), .B1(new_n957), .B2(KEYINPUT45), .ZN(new_n958));
  INV_X1    g533(.A(new_n925), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n960), .A2(KEYINPUT110), .A3(new_n949), .ZN(new_n961));
  NAND2_X1  g536(.A1(G303), .A2(G8), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT55), .Z(new_n963));
  NAND4_X1  g538(.A1(new_n953), .A2(new_n961), .A3(G8), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(G8), .B1(new_n950), .B2(new_n952), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n962), .B(KEYINPUT55), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n693), .A2(G1976), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n499), .A2(new_n908), .A3(new_n923), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(G8), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT52), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  INV_X1    g547(.A(new_n970), .ZN(new_n973));
  INV_X1    g548(.A(G1976), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT52), .B1(G288), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n971), .A2(new_n972), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G48), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n508), .A2(new_n570), .B1(new_n510), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n577), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n573), .B(KEYINPUT77), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n505), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(G1981), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G305), .B2(G1981), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT49), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n982), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n969), .A2(G8), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n968), .A2(new_n975), .A3(new_n969), .A4(G8), .ZN(new_n989));
  OAI22_X1  g564(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(KEYINPUT111), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n976), .A2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n964), .A2(new_n967), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n921), .A2(new_n729), .A3(new_n923), .A4(new_n925), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n993), .A2(new_n994), .B1(new_n934), .B2(new_n748), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n993), .A2(G2078), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n911), .A2(new_n924), .A3(new_n925), .A4(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G171), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT121), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n910), .A2(KEYINPUT120), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n923), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1004), .B2(new_n909), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n921), .A2(KEYINPUT121), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n925), .A2(new_n996), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n995), .A2(G301), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT54), .B1(new_n999), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n992), .B1(new_n1010), .B2(KEYINPUT122), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n995), .A2(G301), .A3(new_n1008), .ZN(new_n1013));
  AOI21_X1  g588(.A(G301), .B1(new_n995), .B2(new_n997), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT122), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n934), .A2(new_n748), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n994), .A2(new_n993), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1008), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1018), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n995), .A2(G301), .A3(new_n997), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(KEYINPUT54), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT123), .B1(new_n1018), .B2(G171), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1011), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT60), .ZN(new_n1025));
  INV_X1    g600(.A(G1348), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n923), .B1(new_n957), .B2(new_n932), .ZN(new_n1027));
  INV_X1    g602(.A(new_n933), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G2067), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n957), .A2(new_n1030), .A3(new_n923), .ZN(new_n1031));
  AND4_X1   g606(.A1(new_n1025), .A2(new_n1029), .A3(new_n856), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1025), .B1(new_n1033), .B2(new_n596), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(new_n856), .A3(new_n1031), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n554), .A2(new_n1037), .A3(new_n559), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n554), .B2(new_n559), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n934), .A2(new_n796), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT115), .B(KEYINPUT56), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(G2072), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n951), .A2(new_n925), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1040), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(new_n1040), .A3(new_n1044), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(KEYINPUT61), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(KEYINPUT116), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1041), .A2(new_n1040), .A3(new_n1050), .A4(new_n1044), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1045), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1036), .B(new_n1048), .C1(new_n1052), .C2(KEYINPUT61), .ZN(new_n1053));
  INV_X1    g628(.A(G1996), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n951), .A2(new_n1054), .A3(new_n925), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT58), .B(G1341), .Z(new_n1056));
  NAND2_X1  g631(.A1(new_n969), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT117), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n537), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT118), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1055), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1060), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1065), .B(new_n537), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1064), .A2(KEYINPUT59), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1062), .B2(new_n537), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1068), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1053), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1045), .B1(new_n856), .B2(new_n1033), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1075), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n946), .B(new_n1024), .C1(new_n1074), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n944), .A2(G8), .A3(G168), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n964), .A2(new_n991), .A3(new_n967), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT114), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1079), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n953), .A2(G8), .A3(new_n961), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1078), .B1(new_n1084), .B2(new_n966), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1083), .A2(new_n964), .A3(new_n991), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n1078), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n974), .B(new_n693), .C1(new_n987), .C2(new_n988), .ZN(new_n1090));
  OR2_X1    g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n988), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n964), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n991), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1077), .A2(new_n1089), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1077), .A2(KEYINPUT124), .A3(new_n1089), .A4(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n946), .A2(KEYINPUT62), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT125), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n942), .A2(new_n1101), .A3(new_n943), .A4(new_n945), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1080), .A2(new_n999), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1099), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT125), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1097), .A2(new_n1098), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n743), .A2(G2067), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n738), .A2(new_n1030), .A3(new_n742), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n921), .A2(new_n910), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(G1996), .A3(new_n724), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n921), .A2(G1996), .A3(new_n910), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n725), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n685), .A2(new_n688), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n685), .A2(new_n688), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1111), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n586), .B(new_n679), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1120), .B1(new_n1111), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1107), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1111), .A2(new_n724), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1112), .A2(KEYINPUT127), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT127), .B1(new_n1112), .B2(new_n1124), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1114), .B(KEYINPUT46), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT47), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1109), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1111), .B1(new_n1131), .B2(KEYINPUT126), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(KEYINPUT126), .B2(new_n1131), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1120), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1111), .A2(new_n679), .A3(new_n586), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT48), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1129), .B(new_n1133), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1123), .A2(new_n1137), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g713(.A(new_n459), .ZN(new_n1140));
  NOR4_X1   g714(.A1(G229), .A2(new_n1140), .A3(G401), .A4(G227), .ZN(new_n1141));
  NAND3_X1  g715(.A1(new_n844), .A2(new_n1141), .A3(new_n899), .ZN(G225));
  INV_X1    g716(.A(G225), .ZN(G308));
endmodule


