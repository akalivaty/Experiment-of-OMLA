//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G116), .A2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  INV_X1    g0008(.A(G244), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n213), .B1(new_n201), .B2(new_n214), .C1(new_n203), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n212), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n217), .B1(G1), .B2(G20), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT1), .Z(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G1), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n224), .A2(new_n221), .A3(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT0), .Z(new_n227));
  NOR3_X1   g0027(.A1(new_n219), .A2(new_n223), .A3(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n230), .B(new_n231), .Z(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G257), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT64), .B(G250), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  INV_X1    g0038(.A(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT65), .B(G107), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(KEYINPUT9), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n204), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n221), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT8), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n202), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT67), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n253), .B1(new_n255), .B2(new_n252), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n221), .A2(G33), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n248), .B1(new_n249), .B2(new_n251), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n222), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n224), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n258), .A2(new_n260), .B1(new_n201), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n224), .B2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  AND3_X1   g0066(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n264), .B1(new_n263), .B2(new_n266), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n247), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n263), .A2(new_n266), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT68), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n263), .A2(new_n264), .A3(new_n266), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(KEYINPUT9), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n250), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G223), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G222), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n283), .C1(G77), .C2(new_n278), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n224), .B1(G41), .B2(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n222), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n250), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n285), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n284), .B(new_n288), .C1(new_n214), .C2(new_n292), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT66), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(KEYINPUT66), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G200), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n295), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G190), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n274), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n274), .A2(new_n301), .A3(new_n296), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT12), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n262), .B(new_n203), .C1(KEYINPUT70), .C2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(KEYINPUT12), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n262), .A2(KEYINPUT70), .A3(new_n304), .A4(new_n203), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n265), .A2(G68), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n203), .A2(G20), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n312), .B1(new_n257), .B2(new_n208), .C1(new_n201), .C2(new_n251), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n313), .B2(new_n260), .ZN(new_n314));
  AND3_X1   g0114(.A1(new_n313), .A2(new_n311), .A3(new_n260), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n309), .B(new_n310), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT71), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT13), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n214), .A2(new_n280), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n278), .B(new_n319), .C1(G232), .C2(new_n280), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n287), .B1(new_n322), .B2(new_n283), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n292), .A2(new_n215), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n318), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n291), .B1(new_n320), .B2(new_n321), .ZN(new_n327));
  NOR4_X1   g0127(.A1(new_n327), .A2(new_n324), .A3(KEYINPUT13), .A4(new_n287), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT69), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT69), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(G200), .C1(new_n326), .C2(new_n328), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n317), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(G190), .ZN(new_n335));
  OAI21_X1  g0135(.A(G169), .B1(new_n326), .B2(new_n328), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(KEYINPUT14), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n329), .A2(G179), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n339), .B(G169), .C1(new_n326), .C2(new_n328), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n334), .A2(new_n335), .B1(new_n341), .B2(new_n317), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT3), .A2(G33), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(G232), .B2(new_n280), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n215), .B2(new_n280), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n283), .C1(G107), .C2(new_n278), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n288), .C1(new_n209), .C2(new_n292), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n262), .A2(new_n208), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n265), .A2(G77), .ZN(new_n353));
  XOR2_X1   g0153(.A(KEYINPUT15), .B(G87), .Z(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT8), .B(G58), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n355), .A2(new_n257), .B1(new_n251), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(G20), .B2(G77), .ZN(new_n358));
  INV_X1    g0158(.A(new_n260), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n352), .B(new_n353), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n351), .B(new_n360), .C1(G179), .C2(new_n349), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n270), .B1(new_n297), .B2(G169), .ZN(new_n362));
  AOI21_X1  g0162(.A(G179), .B1(new_n294), .B2(new_n295), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n360), .B1(new_n349), .B2(G200), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n349), .ZN(new_n367));
  AND4_X1   g0167(.A1(new_n342), .A2(new_n361), .A3(new_n364), .A4(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT18), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n214), .A2(G1698), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n278), .B(new_n370), .C1(G223), .C2(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G33), .A2(G87), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n291), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n291), .A2(G232), .A3(new_n285), .ZN(new_n374));
  INV_X1    g0174(.A(G179), .ZN(new_n375));
  NOR4_X1   g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .A4(new_n287), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n373), .A2(new_n374), .A3(new_n287), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n376), .B1(new_n378), .B2(G169), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT7), .B1(new_n345), .B2(new_n221), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n221), .A4(new_n277), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT74), .ZN(new_n384));
  INV_X1    g0184(.A(G159), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n251), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n202), .A2(KEYINPUT67), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT67), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G58), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n387), .A2(new_n389), .A3(G68), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G58), .B2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n386), .B1(new_n391), .B2(G20), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n276), .A2(new_n221), .A3(new_n277), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(new_n381), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT74), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n397), .A3(G68), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n384), .A2(new_n392), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n395), .A2(KEYINPUT72), .A3(new_n381), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n381), .B2(KEYINPUT72), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT16), .B(new_n392), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT73), .ZN(new_n405));
  INV_X1    g0205(.A(new_n403), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT72), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n396), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(KEYINPUT16), .A4(new_n392), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n401), .A2(new_n260), .A3(new_n405), .A4(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n265), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n256), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n256), .B2(new_n262), .ZN(new_n414));
  AOI211_X1 g0214(.A(new_n369), .B(new_n379), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n405), .A2(new_n260), .A3(new_n410), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n399), .A2(new_n400), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n379), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT18), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n377), .A2(new_n366), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n377), .B2(G200), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n411), .A2(new_n414), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n411), .A2(KEYINPUT17), .A3(new_n414), .A4(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n421), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n303), .A2(new_n368), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT75), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n303), .A2(new_n368), .A3(new_n429), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G107), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n224), .A2(new_n435), .A3(G13), .A4(G20), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT25), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n224), .A2(G33), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n359), .A2(new_n261), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n437), .B1(new_n440), .B2(G107), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n221), .B(G87), .C1(new_n343), .C2(new_n344), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT22), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n278), .A2(KEYINPUT22), .A3(new_n221), .A4(G87), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT23), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT82), .B1(new_n221), .B2(G107), .ZN(new_n448));
  NAND2_X1  g0248(.A1(KEYINPUT82), .A2(KEYINPUT23), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G116), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n447), .A2(new_n448), .B1(new_n451), .B2(new_n221), .ZN(new_n452));
  NAND3_X1  g0252(.A1(KEYINPUT82), .A2(KEYINPUT23), .A3(G107), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n445), .A2(new_n446), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(KEYINPUT24), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n454), .A2(KEYINPUT24), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n260), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT82), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(G20), .B2(new_n435), .ZN(new_n461));
  AOI22_X1  g0261(.A1(KEYINPUT82), .A2(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n461), .A2(KEYINPUT23), .B1(new_n462), .B2(G20), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n444), .B2(new_n443), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(new_n453), .A4(new_n446), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n454), .A2(KEYINPUT24), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(KEYINPUT83), .A3(new_n260), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n442), .B1(new_n459), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n278), .B1(G257), .B2(new_n280), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G250), .A2(G1698), .ZN(new_n472));
  INV_X1    g0272(.A(G294), .ZN(new_n473));
  OAI22_X1  g0273(.A1(new_n471), .A2(new_n472), .B1(new_n250), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT5), .A2(G41), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n479), .A2(new_n291), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n474), .A2(new_n283), .B1(G264), .B2(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n479), .A2(new_n286), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n330), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(G190), .B2(new_n483), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n470), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(KEYINPUT83), .B1(new_n468), .B2(new_n260), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n458), .B(new_n359), .C1(new_n466), .C2(new_n467), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n441), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(G169), .B1(new_n481), .B2(new_n482), .ZN(new_n490));
  INV_X1    g0290(.A(new_n483), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n375), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n221), .B(G68), .C1(new_n343), .C2(new_n344), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT19), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n210), .A2(new_n496), .A3(new_n435), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n321), .A2(new_n221), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n321), .A2(KEYINPUT19), .A3(G20), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT77), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT77), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n503), .B(new_n494), .C1(new_n499), .C2(new_n500), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n260), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n354), .A2(new_n261), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n355), .B2(new_n439), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n291), .B(G250), .C1(G1), .C2(new_n475), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n476), .A2(G274), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n276), .A2(new_n277), .B1(new_n209), .B2(G1698), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n215), .A2(new_n280), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n512), .A2(new_n513), .B1(G33), .B2(G116), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n510), .B(new_n511), .C1(new_n514), .C2(new_n291), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n350), .ZN(new_n516));
  INV_X1    g0316(.A(new_n515), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n375), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n486), .A2(new_n493), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n280), .A2(G257), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G264), .A2(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n343), .C2(new_n344), .ZN(new_n523));
  INV_X1    g0323(.A(G303), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n276), .A2(new_n524), .A3(new_n277), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n283), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n523), .A2(KEYINPUT79), .A3(new_n525), .A4(new_n283), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n529), .B1(new_n480), .B2(G270), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n350), .B1(new_n530), .B2(new_n482), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n262), .A2(new_n239), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n359), .A2(G116), .A3(new_n261), .A4(new_n438), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n259), .A2(new_n222), .B1(G20), .B2(new_n239), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G283), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n221), .C1(G33), .C2(new_n496), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT20), .B1(new_n534), .B2(new_n536), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n532), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT80), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n239), .A2(G20), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(new_n260), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT20), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n534), .A2(KEYINPUT20), .A3(new_n536), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT80), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(new_n532), .A4(new_n533), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n540), .A2(new_n548), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n531), .A2(new_n549), .A3(KEYINPUT21), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT21), .B1(new_n531), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n528), .A2(new_n529), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n480), .A2(G270), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n552), .A2(G179), .A3(new_n482), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n548), .B2(new_n540), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT81), .ZN(new_n557));
  INV_X1    g0357(.A(new_n549), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n530), .A2(new_n482), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G200), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n560), .C1(new_n366), .C2(new_n559), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n531), .A2(new_n549), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n531), .A2(new_n549), .A3(KEYINPUT21), .ZN(new_n566));
  INV_X1    g0366(.A(new_n555), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n561), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT81), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n515), .A2(new_n366), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n515), .A2(G200), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n440), .A2(G87), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n572), .A2(new_n507), .A3(new_n505), .A4(new_n573), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n574), .A2(KEYINPUT78), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(KEYINPUT78), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n571), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT4), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(G1698), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n579), .B(G244), .C1(new_n344), .C2(new_n343), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n209), .B1(new_n276), .B2(new_n277), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n535), .C1(new_n581), .C2(KEYINPUT4), .ZN(new_n582));
  OAI21_X1  g0382(.A(G250), .B1(new_n343), .B2(new_n344), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n280), .B1(new_n583), .B2(KEYINPUT4), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n283), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n480), .A2(G257), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n482), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT76), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n585), .A2(new_n589), .A3(new_n482), .A4(new_n586), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(G200), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n261), .A2(G97), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n439), .A2(new_n496), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n396), .A2(G107), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n221), .A2(new_n250), .A3(G77), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n435), .A2(KEYINPUT6), .A3(G97), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n496), .A2(new_n435), .ZN(new_n597));
  NOR2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n599), .B2(KEYINPUT6), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G20), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n594), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  AOI211_X1 g0402(.A(new_n592), .B(new_n593), .C1(new_n602), .C2(new_n260), .ZN(new_n603));
  INV_X1    g0403(.A(new_n587), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G190), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n591), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n592), .B1(new_n602), .B2(new_n260), .ZN(new_n607));
  INV_X1    g0407(.A(new_n593), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n375), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n587), .A2(new_n350), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n577), .A2(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n434), .A2(new_n520), .A3(new_n570), .A4(new_n614), .ZN(G372));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n577), .A2(new_n616), .A3(new_n612), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n493), .A2(new_n556), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n574), .A2(new_n571), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n470), .B2(new_n485), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n618), .A2(new_n606), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n612), .A2(new_n619), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(KEYINPUT26), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n617), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n519), .ZN(new_n625));
  OR2_X1    g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n434), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n364), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n303), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n300), .A2(KEYINPUT84), .A3(new_n302), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n415), .A2(new_n420), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n361), .B1(new_n334), .B2(new_n335), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n317), .B2(new_n341), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n428), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n628), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n627), .A2(new_n637), .ZN(G369));
  INV_X1    g0438(.A(G13), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n224), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n556), .A2(new_n558), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n549), .A2(new_n646), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n570), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G330), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n489), .A2(new_n492), .A3(new_n647), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n486), .B1(new_n470), .B2(new_n647), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(new_n493), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n556), .A2(new_n646), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n654), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(new_n660), .ZN(G399));
  NOR2_X1   g0461(.A1(new_n497), .A2(G116), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT85), .Z(new_n663));
  INV_X1    g0463(.A(new_n225), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n663), .A2(new_n224), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n220), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(new_n665), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n668), .B(KEYINPUT28), .Z(new_n669));
  NAND4_X1  g0469(.A1(new_n570), .A2(new_n520), .A3(new_n614), .A4(new_n647), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n554), .A2(new_n515), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(new_n491), .A3(new_n585), .A4(new_n586), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT30), .Z(new_n673));
  NAND3_X1  g0473(.A1(new_n483), .A2(new_n375), .A3(new_n515), .ZN(new_n674));
  AOI211_X1 g0474(.A(new_n604), .B(new_n674), .C1(new_n482), .C2(new_n530), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n646), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n676), .A2(KEYINPUT31), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n682), .B(new_n647), .C1(new_n624), .C2(new_n625), .ZN(new_n683));
  INV_X1    g0483(.A(new_n612), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT78), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n574), .B(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n616), .B(new_n684), .C1(new_n686), .C2(new_n571), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT26), .B1(new_n612), .B2(new_n619), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n687), .A2(new_n519), .A3(new_n688), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n606), .A2(KEYINPUT86), .A3(new_n612), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT86), .B1(new_n606), .B2(new_n612), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n618), .B(new_n620), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n646), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n683), .B1(new_n682), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n681), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n669), .B1(new_n695), .B2(G1), .ZN(G364));
  NAND2_X1  g0496(.A1(new_n640), .A2(G45), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT87), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G1), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(new_n665), .ZN(new_n701));
  INV_X1    g0501(.A(new_n652), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n650), .A2(new_n651), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n701), .ZN(new_n705));
  NOR2_X1   g0505(.A1(G13), .A2(G33), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G20), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n222), .B1(G20), .B2(new_n350), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n664), .A2(new_n278), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n667), .A2(new_n475), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n711), .B(new_n712), .C1(new_n245), .C2(new_n475), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n278), .A2(new_n225), .A3(G355), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n713), .B(new_n714), .C1(G116), .C2(new_n225), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n650), .A2(new_n708), .B1(new_n710), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n221), .A2(new_n366), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n330), .A2(G179), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n210), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n221), .A2(G190), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT88), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n722), .A2(G179), .A3(new_n330), .ZN(new_n723));
  AOI211_X1 g0523(.A(new_n345), .B(new_n720), .C1(new_n723), .C2(G107), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT89), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n375), .A2(G200), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n375), .A2(new_n330), .ZN(new_n728));
  AND2_X1   g0528(.A1(new_n728), .A2(new_n721), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n727), .A2(new_n254), .B1(new_n729), .B2(G68), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n721), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G179), .A2(G200), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n221), .B1(new_n732), .B2(G190), .ZN(new_n733));
  OAI221_X1 g0533(.A(new_n730), .B1(new_n208), .B2(new_n731), .C1(new_n496), .C2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT32), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n722), .A2(G179), .A3(G200), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n737), .B2(new_n385), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n736), .A2(KEYINPUT32), .A3(G159), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n717), .A2(new_n728), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n725), .B(new_n740), .C1(new_n201), .C2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n727), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(G283), .A2(new_n723), .B1(new_n736), .B2(G329), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n731), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G326), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n741), .A2(new_n749), .B1(new_n719), .B2(new_n524), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT33), .B(G317), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n748), .B(new_n750), .C1(new_n729), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n733), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n278), .B1(new_n753), .B2(G294), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n746), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n742), .B1(new_n745), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n709), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n705), .B1(new_n716), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n704), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT90), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(G396));
  INV_X1    g0561(.A(new_n723), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n203), .ZN(new_n763));
  INV_X1    g0563(.A(G132), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n278), .B1(new_n255), .B2(new_n733), .C1(new_n737), .C2(new_n764), .ZN(new_n765));
  AOI22_X1  g0565(.A1(new_n727), .A2(G143), .B1(new_n729), .B2(G150), .ZN(new_n766));
  INV_X1    g0566(.A(G137), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n766), .B1(new_n767), .B2(new_n741), .C1(new_n385), .C2(new_n731), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT91), .Z(new_n769));
  AOI211_X1 g0569(.A(new_n763), .B(new_n765), .C1(new_n769), .C2(KEYINPUT34), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n770), .B1(KEYINPUT34), .B2(new_n769), .C1(new_n201), .C2(new_n719), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n345), .B1(new_n731), .B2(new_n239), .ZN(new_n772));
  INV_X1    g0572(.A(new_n741), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G303), .B1(new_n729), .B2(G283), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n774), .B1(new_n435), .B2(new_n719), .C1(new_n473), .C2(new_n743), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n772), .B(new_n775), .C1(G97), .C2(new_n753), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n776), .B1(new_n210), .B2(new_n762), .C1(new_n747), .C2(new_n737), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n771), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n705), .B1(new_n778), .B2(new_n709), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n709), .A2(new_n706), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(new_n208), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n360), .A2(new_n646), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n367), .A2(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(new_n361), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n361), .A2(new_n646), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n779), .B(new_n781), .C1(new_n707), .C2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n647), .B(new_n786), .C1(new_n624), .C2(new_n625), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(KEYINPUT92), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n680), .B(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n786), .B1(new_n626), .B2(new_n647), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n790), .B(new_n791), .Z(new_n792));
  OAI21_X1  g0592(.A(new_n787), .B1(new_n792), .B2(new_n701), .ZN(G384));
  NAND2_X1  g0593(.A1(new_n317), .A2(new_n646), .ZN(new_n794));
  AOI21_X1  g0594(.A(KEYINPUT93), .B1(new_n342), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n316), .B(KEYINPUT71), .Z(new_n796));
  OAI21_X1  g0596(.A(G200), .B1(new_n326), .B2(new_n328), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n797), .A2(KEYINPUT69), .ZN(new_n798));
  INV_X1    g0598(.A(new_n333), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n335), .B(new_n796), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n341), .A2(new_n317), .ZN(new_n801));
  AND4_X1   g0601(.A1(KEYINPUT93), .A2(new_n800), .A3(new_n801), .A4(new_n794), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n795), .A2(new_n802), .B1(new_n801), .B2(new_n647), .ZN(new_n803));
  AND4_X1   g0603(.A1(new_n677), .A2(new_n803), .A3(new_n678), .A4(new_n786), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n400), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n405), .A2(new_n806), .A3(new_n410), .A4(new_n260), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n414), .ZN(new_n808));
  INV_X1    g0608(.A(new_n644), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n421), .B2(new_n428), .ZN(new_n812));
  XOR2_X1   g0612(.A(new_n644), .B(KEYINPUT94), .Z(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n418), .B1(new_n419), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n816), .A3(new_n424), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n808), .A2(new_n419), .ZN(new_n818));
  AND3_X1   g0618(.A1(new_n810), .A2(new_n818), .A3(new_n424), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n817), .B1(new_n819), .B2(new_n816), .ZN(new_n820));
  AOI21_X1  g0620(.A(KEYINPUT38), .B1(new_n812), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n812), .A2(KEYINPUT38), .A3(new_n820), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(KEYINPUT95), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT95), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n812), .A2(KEYINPUT38), .A3(new_n820), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n825), .B1(new_n826), .B2(new_n821), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n804), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT40), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(KEYINPUT97), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(KEYINPUT97), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n828), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT96), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n823), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n418), .A2(new_n814), .ZN(new_n837));
  INV_X1    g0637(.A(new_n428), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n633), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n424), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n411), .A2(new_n414), .B1(new_n379), .B2(new_n813), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT37), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n842), .A2(new_n817), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n836), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n812), .A2(new_n820), .A3(KEYINPUT96), .A4(KEYINPUT38), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n835), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n804), .A2(KEYINPUT40), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n833), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n434), .A2(new_n679), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n849), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G330), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT39), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n826), .A2(new_n821), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n853), .B2(new_n846), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n801), .A2(new_n646), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n421), .A2(new_n813), .ZN(new_n858));
  INV_X1    g0658(.A(new_n785), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n788), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n824), .A2(new_n827), .A3(new_n860), .A4(new_n803), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n434), .A2(new_n694), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n863), .A2(new_n637), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n862), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n852), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n224), .B2(new_n640), .ZN(new_n867));
  OAI211_X1 g0667(.A(G20), .B(new_n289), .C1(new_n600), .C2(KEYINPUT35), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n239), .B(new_n868), .C1(KEYINPUT35), .C2(new_n600), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  NAND3_X1  g0670(.A1(new_n390), .A2(G77), .A3(new_n667), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(G50), .B2(new_n203), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(G1), .A3(new_n639), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n867), .A2(new_n870), .A3(new_n873), .ZN(G367));
  OAI22_X1  g0674(.A1(new_n690), .A2(new_n691), .B1(new_n603), .B2(new_n647), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n684), .A2(new_n646), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n657), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT42), .ZN(new_n881));
  INV_X1    g0681(.A(new_n875), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n659), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT99), .Z(new_n884));
  NAND2_X1  g0684(.A1(new_n508), .A2(new_n573), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n646), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n519), .B1(new_n887), .B2(new_n619), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n519), .B2(new_n887), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n881), .B1(new_n659), .B2(new_n882), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n612), .B1(new_n875), .B2(new_n493), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n892), .B1(new_n893), .B2(new_n647), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n884), .A2(new_n891), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT100), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n891), .B1(new_n884), .B2(new_n894), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT43), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n889), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n879), .A2(KEYINPUT101), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n880), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI211_X1 g0702(.A(KEYINPUT101), .B(new_n879), .C1(new_n896), .C2(new_n899), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n665), .B(KEYINPUT41), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n656), .B(new_n658), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT106), .Z(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n652), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(KEYINPUT106), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n652), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n695), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OR3_X1    g0714(.A1(new_n660), .A2(KEYINPUT44), .A3(new_n877), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT44), .B1(new_n660), .B2(new_n877), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT45), .Z(new_n919));
  NAND3_X1  g0719(.A1(new_n660), .A2(new_n877), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n919), .ZN(new_n921));
  INV_X1    g0721(.A(new_n660), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n921), .B1(new_n922), .B2(new_n878), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n917), .A2(KEYINPUT104), .A3(new_n920), .A4(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n657), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n923), .A2(new_n915), .A3(new_n916), .A4(new_n920), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT104), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT105), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n926), .A2(new_n925), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n914), .B(new_n932), .C1(new_n930), .C2(new_n929), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n906), .B1(new_n933), .B2(new_n695), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n904), .B1(new_n934), .B2(new_n700), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n723), .A2(G97), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n773), .A2(G311), .B1(new_n727), .B2(G303), .ZN(new_n937));
  INV_X1    g0737(.A(G317), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n936), .B(new_n937), .C1(new_n737), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n719), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(G116), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT46), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n278), .B1(new_n753), .B2(G107), .ZN(new_n943));
  INV_X1    g0743(.A(G283), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n942), .B(new_n943), .C1(new_n944), .C2(new_n731), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n939), .B(new_n945), .C1(G294), .C2(new_n729), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT107), .Z(new_n947));
  OAI22_X1  g0747(.A1(new_n208), .A2(new_n762), .B1(new_n737), .B2(new_n767), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(G68), .B2(new_n753), .ZN(new_n949));
  INV_X1    g0749(.A(new_n731), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n773), .A2(G143), .B1(new_n950), .B2(G50), .ZN(new_n951));
  OAI221_X1 g0751(.A(new_n951), .B1(new_n249), .B2(new_n743), .C1(new_n255), .C2(new_n719), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G159), .B2(new_n729), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n278), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n947), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n705), .B1(new_n956), .B2(new_n709), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n236), .A2(new_n711), .B1(new_n664), .B2(new_n354), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n710), .ZN(new_n959));
  INV_X1    g0759(.A(new_n708), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n957), .B(new_n959), .C1(new_n960), .C2(new_n890), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n935), .A2(new_n961), .ZN(G387));
  INV_X1    g0762(.A(new_n709), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n719), .A2(new_n473), .B1(new_n733), .B2(new_n944), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT111), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n727), .A2(G317), .B1(new_n729), .B2(G311), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n524), .B2(new_n731), .C1(new_n744), .C2(new_n741), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT48), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT112), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n967), .A2(new_n968), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT49), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n723), .A2(G116), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n970), .A2(KEYINPUT49), .A3(new_n971), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n278), .B1(new_n736), .B2(G326), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n950), .A2(G68), .B1(new_n727), .B2(G50), .ZN(new_n979));
  INV_X1    g0779(.A(new_n729), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n979), .B1(new_n256), .B2(new_n980), .C1(new_n355), .C2(new_n733), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n345), .B1(new_n940), .B2(G77), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n936), .B(new_n982), .C1(new_n737), .C2(new_n249), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT110), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n984), .B2(new_n983), .C1(new_n385), .C2(new_n741), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n963), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n663), .A2(new_n225), .A3(new_n278), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT108), .ZN(new_n989));
  INV_X1    g0789(.A(new_n232), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n989), .B1(new_n990), .B2(new_n475), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n232), .A2(KEYINPUT108), .A3(G45), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n991), .A2(new_n711), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n356), .A2(G50), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT109), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n475), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(KEYINPUT50), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n203), .A2(new_n208), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n663), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n988), .B1(G107), .B2(new_n225), .C1(new_n993), .C2(new_n1000), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n705), .B(new_n987), .C1(new_n710), .C2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT113), .Z(new_n1003));
  OR2_X1    g0803(.A1(new_n656), .A2(new_n960), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n911), .A2(new_n700), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n665), .B1(new_n911), .B2(new_n695), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n914), .B2(new_n1006), .ZN(G393));
  AND2_X1   g0807(.A1(new_n926), .A2(new_n925), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n912), .A2(new_n913), .B1(new_n931), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n933), .A2(new_n1009), .A3(new_n665), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n700), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n1008), .A2(new_n931), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n773), .A2(G150), .B1(new_n727), .B2(G159), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT51), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n210), .C2(new_n762), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n731), .A2(new_n356), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n345), .B(new_n1017), .C1(G50), .C2(new_n729), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n203), .B2(new_n719), .C1(new_n208), .C2(new_n733), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(G143), .C2(new_n736), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n731), .A2(new_n473), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n345), .B1(new_n980), .B2(new_n524), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G116), .C2(new_n753), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n743), .A2(new_n747), .B1(new_n938), .B2(new_n741), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT52), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G107), .A2(new_n723), .B1(new_n736), .B2(G322), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G283), .B2(new_n940), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n709), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n709), .B(new_n708), .C1(new_n242), .C2(new_n711), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n664), .A2(G97), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n705), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n1032), .C1(new_n877), .C2(new_n960), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1012), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT114), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT114), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1012), .A2(new_n1036), .A3(new_n1033), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1010), .A2(new_n1038), .ZN(G390));
  NAND3_X1  g0839(.A1(new_n434), .A2(G330), .A3(new_n679), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1040), .A2(new_n863), .A3(new_n637), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n677), .A2(new_n678), .A3(new_n786), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1042), .A2(G330), .A3(new_n803), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n646), .B(new_n784), .C1(new_n689), .C2(new_n692), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT116), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n785), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n689), .A2(new_n692), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n784), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n647), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT116), .B1(new_n1050), .B2(new_n859), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n803), .B1(new_n1042), .B2(G330), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n1044), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1042), .A2(G330), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n803), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1057), .A2(new_n1043), .B1(new_n859), .B2(new_n788), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1041), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT117), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n856), .B(KEYINPUT115), .Z(new_n1061));
  NAND2_X1  g0861(.A1(new_n846), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1052), .B2(new_n803), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n846), .A2(new_n853), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n854), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n860), .A2(new_n803), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n856), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1064), .A2(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1060), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1046), .B1(new_n1045), .B2(new_n785), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1050), .A2(KEYINPUT116), .A3(new_n859), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n803), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1072), .A2(new_n846), .A3(new_n1061), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n856), .B1(new_n860), .B2(new_n803), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1073), .B(KEYINPUT117), .C1(new_n855), .C2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1069), .A2(new_n1075), .A3(new_n1043), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1068), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1077), .A2(KEYINPUT117), .A3(new_n1073), .A4(new_n1044), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1059), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n665), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1059), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT119), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1011), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n762), .A2(new_n201), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  AOI211_X1 g0888(.A(new_n345), .B(new_n1087), .C1(new_n950), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(G125), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n737), .C1(new_n767), .C2(new_n980), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n743), .A2(new_n764), .B1(new_n1092), .B2(new_n741), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT118), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n385), .B2(new_n733), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n940), .A2(G150), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT53), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1091), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n203), .A2(new_n762), .B1(new_n737), .B2(new_n473), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n727), .A2(G116), .B1(new_n729), .B2(G107), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n496), .B2(new_n731), .C1(new_n944), .C2(new_n741), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n345), .B1(new_n733), .B2(new_n208), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1099), .A2(new_n720), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n709), .B1(new_n1098), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n701), .B(new_n1104), .C1(new_n855), .C2(new_n707), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n256), .B2(new_n780), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1085), .B1(new_n1086), .B2(new_n1106), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n1086), .A2(new_n1085), .A3(new_n1106), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1084), .A2(new_n1107), .A3(new_n1108), .ZN(G378));
  NAND3_X1  g0909(.A1(new_n848), .A2(G330), .A3(new_n862), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n857), .A2(new_n858), .A3(new_n861), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n833), .A2(G330), .A3(new_n847), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n630), .A2(new_n364), .A3(new_n631), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT121), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT121), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n630), .A2(new_n1118), .A3(new_n364), .A4(new_n631), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n267), .A2(new_n268), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n809), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1115), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1121), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1114), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1110), .A2(new_n1113), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1130), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n290), .B(new_n345), .C1(new_n719), .C2(new_n208), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n773), .A2(G116), .B1(new_n727), .B2(G107), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1136), .B1(new_n496), .B2(new_n980), .C1(new_n355), .C2(new_n731), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(G68), .C2(new_n753), .ZN(new_n1138));
  OAI221_X1 g0938(.A(new_n1138), .B1(new_n944), .B2(new_n737), .C1(new_n255), .C2(new_n762), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT58), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n201), .B1(new_n343), .B2(G41), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n741), .A2(new_n1090), .B1(new_n733), .B2(new_n249), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n940), .A2(new_n1088), .B1(new_n727), .B2(G128), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n767), .B2(new_n731), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G132), .C2(new_n729), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT59), .ZN(new_n1146));
  AOI21_X1  g0946(.A(G41), .B1(new_n736), .B2(G124), .ZN(new_n1147));
  AOI21_X1  g0947(.A(G33), .B1(new_n723), .B2(G159), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1140), .A2(new_n1141), .A3(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1134), .A2(new_n706), .B1(new_n709), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n705), .B1(new_n201), .B2(new_n780), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT120), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1133), .A2(new_n700), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1131), .A2(new_n1132), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT122), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n1041), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1041), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1079), .A2(KEYINPUT122), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1156), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n665), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n1157), .A3(new_n1041), .ZN(new_n1164));
  OAI21_X1  g0964(.A(KEYINPUT122), .B1(new_n1079), .B2(new_n1160), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT57), .B1(new_n1166), .B2(new_n1133), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1154), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT123), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1134), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1110), .A2(new_n1113), .A3(new_n1130), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1162), .B(new_n665), .C1(new_n1174), .C2(KEYINPUT57), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT123), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n1154), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1169), .A2(new_n1177), .ZN(G375));
  NOR2_X1   g0978(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n780), .A2(new_n203), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n803), .A2(new_n707), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n278), .B1(new_n723), .B2(G77), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT125), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n355), .A2(new_n733), .B1(new_n496), .B2(new_n719), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n727), .A2(G283), .B1(new_n729), .B2(G116), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n473), .B2(new_n741), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1185), .B(new_n1187), .C1(G303), .C2(new_n736), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1184), .B(new_n1188), .C1(new_n435), .C2(new_n731), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1092), .A2(new_n737), .B1(new_n762), .B2(new_n255), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n773), .A2(G132), .B1(new_n729), .B2(new_n1088), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n249), .B2(new_n731), .C1(new_n385), .C2(new_n719), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n278), .B1(new_n733), .B2(new_n201), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n767), .B2(new_n743), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n963), .B1(new_n1189), .B2(new_n1195), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1182), .A2(new_n705), .A3(new_n1196), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1180), .A2(new_n700), .B1(new_n1181), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1179), .A2(new_n1160), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n905), .B(KEYINPUT124), .Z(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1059), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1198), .A2(new_n1202), .ZN(G381));
  AND3_X1   g1003(.A1(new_n1175), .A2(new_n1176), .A3(new_n1154), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1176), .B1(new_n1175), .B2(new_n1154), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1204), .A2(new_n1205), .A3(G378), .ZN(new_n1206));
  INV_X1    g1006(.A(G390), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n935), .A3(new_n961), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G393), .A2(G396), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1208), .A2(G384), .A3(G381), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1206), .A2(new_n1211), .ZN(G407));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n645), .ZN(new_n1213));
  INV_X1    g1013(.A(G378), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1169), .A2(new_n1214), .A3(new_n1177), .ZN(new_n1215));
  OAI21_X1  g1015(.A(G213), .B1(new_n1213), .B2(new_n1215), .ZN(G409));
  NAND2_X1  g1016(.A1(new_n1208), .A2(KEYINPUT127), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1207), .B1(new_n935), .B2(new_n961), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT126), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1210), .B2(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1210), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1217), .A2(new_n1218), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G387), .A2(G390), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(new_n1221), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1224), .A2(new_n1225), .A3(KEYINPUT127), .A4(new_n1208), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT61), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1214), .B1(new_n1175), .B2(new_n1154), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1133), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1154), .B1(new_n1230), .B2(new_n1200), .ZN(new_n1231));
  INV_X1    g1031(.A(G213), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1231), .A2(G378), .B1(new_n1232), .B2(G343), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT60), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1199), .A2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1179), .A2(KEYINPUT60), .A3(new_n1160), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1235), .A2(new_n665), .A3(new_n1059), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1198), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(G384), .A3(new_n1198), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1229), .A2(new_n1233), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT62), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1228), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n645), .A2(G213), .A3(G2897), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1242), .B(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1229), .B2(new_n1233), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1168), .A2(G378), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1173), .B2(new_n1011), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1174), .B2(new_n1201), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1252), .A2(new_n1214), .B1(G213), .B2(new_n645), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1242), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1249), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT62), .B1(new_n1248), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1227), .B1(new_n1245), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1248), .A2(new_n1255), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(KEYINPUT63), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1228), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(KEYINPUT63), .B2(new_n1243), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1257), .B1(new_n1260), .B2(new_n1262), .ZN(G405));
  AND3_X1   g1063(.A1(new_n1215), .A2(new_n1242), .A3(new_n1249), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1242), .B1(new_n1215), .B2(new_n1249), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1264), .A2(new_n1265), .A3(new_n1227), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1254), .B1(new_n1206), .B2(new_n1229), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1215), .A2(new_n1242), .A3(new_n1249), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1261), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1266), .A2(new_n1269), .ZN(G402));
endmodule


