

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  NOR2_X1 U321 ( .A1(n529), .A2(n446), .ZN(n561) );
  XOR2_X1 U322 ( .A(n405), .B(n352), .Z(n289) );
  XNOR2_X1 U323 ( .A(n420), .B(KEYINPUT123), .ZN(n421) );
  INV_X1 U324 ( .A(KEYINPUT68), .ZN(n355) );
  XNOR2_X1 U325 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U326 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U327 ( .A(n358), .B(n357), .ZN(n359) );
  INV_X1 U328 ( .A(G190GAT), .ZN(n447) );
  XNOR2_X1 U329 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U330 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT84), .B(G176GAT), .Z(n291) );
  NAND2_X1 U332 ( .A1(G227GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U333 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U334 ( .A(KEYINPUT20), .B(G190GAT), .Z(n293) );
  XNOR2_X1 U335 ( .A(G43GAT), .B(G99GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U337 ( .A(n295), .B(n294), .Z(n300) );
  XOR2_X1 U338 ( .A(KEYINPUT18), .B(KEYINPUT83), .Z(n297) );
  XNOR2_X1 U339 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(KEYINPUT17), .B(n298), .Z(n419) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(n419), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U344 ( .A(G15GAT), .B(G127GAT), .Z(n390) );
  XOR2_X1 U345 ( .A(n301), .B(n390), .Z(n305) );
  XOR2_X1 U346 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n303) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G134GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n323) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n371) );
  XNOR2_X1 U350 ( .A(n323), .B(n371), .ZN(n304) );
  XOR2_X1 U351 ( .A(n305), .B(n304), .Z(n476) );
  INV_X1 U352 ( .A(n476), .ZN(n529) );
  XOR2_X1 U353 ( .A(G85GAT), .B(G155GAT), .Z(n307) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(G162GAT), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U356 ( .A(KEYINPUT6), .B(G148GAT), .Z(n309) );
  XNOR2_X1 U357 ( .A(G120GAT), .B(G127GAT), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U359 ( .A(n311), .B(n310), .Z(n316) );
  XOR2_X1 U360 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n313) );
  NAND2_X1 U361 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U363 ( .A(KEYINPUT5), .B(n314), .ZN(n315) );
  XNOR2_X1 U364 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U365 ( .A(G57GAT), .B(KEYINPUT92), .Z(n318) );
  XNOR2_X1 U366 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U368 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n322) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n430) );
  XNOR2_X1 U372 ( .A(n323), .B(n430), .ZN(n324) );
  XOR2_X1 U373 ( .A(n325), .B(n324), .Z(n514) );
  INV_X1 U374 ( .A(n514), .ZN(n542) );
  XOR2_X1 U375 ( .A(KEYINPUT73), .B(KEYINPUT71), .Z(n327) );
  XNOR2_X1 U376 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n327), .B(n326), .ZN(n332) );
  XNOR2_X1 U378 ( .A(G36GAT), .B(G190GAT), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n328), .B(G218GAT), .ZN(n415) );
  XOR2_X1 U380 ( .A(KEYINPUT75), .B(n415), .Z(n330) );
  XOR2_X1 U381 ( .A(G50GAT), .B(G162GAT), .Z(n433) );
  XNOR2_X1 U382 ( .A(G134GAT), .B(n433), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n343) );
  XOR2_X1 U385 ( .A(KEYINPUT72), .B(KEYINPUT74), .Z(n334) );
  NAND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U388 ( .A(n335), .B(KEYINPUT9), .Z(n341) );
  XOR2_X1 U389 ( .A(G29GAT), .B(G43GAT), .Z(n337) );
  XNOR2_X1 U390 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n354) );
  XOR2_X1 U392 ( .A(G92GAT), .B(G85GAT), .Z(n339) );
  XNOR2_X1 U393 ( .A(G99GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n366) );
  XNOR2_X1 U395 ( .A(n354), .B(n366), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n552) );
  XOR2_X1 U398 ( .A(G1GAT), .B(G15GAT), .Z(n345) );
  XNOR2_X1 U399 ( .A(G141GAT), .B(G113GAT), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U401 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n347) );
  XNOR2_X1 U402 ( .A(KEYINPUT67), .B(KEYINPUT30), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n360) );
  XOR2_X1 U405 ( .A(G169GAT), .B(G8GAT), .Z(n405) );
  XOR2_X1 U406 ( .A(G22GAT), .B(G197GAT), .Z(n351) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G50GAT), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  NAND2_X1 U409 ( .A1(G229GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n289), .B(n353), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n354), .B(KEYINPUT65), .ZN(n356) );
  XOR2_X1 U412 ( .A(n360), .B(n359), .Z(n565) );
  INV_X1 U413 ( .A(n565), .ZN(n555) );
  XOR2_X1 U414 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n362) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U417 ( .A(n363), .B(KEYINPUT31), .Z(n368) );
  XOR2_X1 U418 ( .A(G64GAT), .B(KEYINPUT70), .Z(n365) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(G204GAT), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n406) );
  XNOR2_X1 U421 ( .A(n406), .B(n366), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n368), .B(n367), .ZN(n370) );
  XNOR2_X1 U423 ( .A(G57GAT), .B(KEYINPUT69), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n369), .B(KEYINPUT13), .ZN(n388) );
  XOR2_X1 U425 ( .A(n370), .B(n388), .Z(n373) );
  XOR2_X1 U426 ( .A(G148GAT), .B(G78GAT), .Z(n427) );
  XNOR2_X1 U427 ( .A(n371), .B(n427), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n570) );
  XOR2_X1 U429 ( .A(n570), .B(KEYINPUT41), .Z(n557) );
  NAND2_X1 U430 ( .A1(n555), .A2(n557), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n374), .B(KEYINPUT46), .ZN(n395) );
  XOR2_X1 U432 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n376) );
  XNOR2_X1 U433 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n394) );
  XOR2_X1 U435 ( .A(G78GAT), .B(G211GAT), .Z(n378) );
  XNOR2_X1 U436 ( .A(G183GAT), .B(G71GAT), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U438 ( .A(KEYINPUT77), .B(G64GAT), .Z(n380) );
  XNOR2_X1 U439 ( .A(G1GAT), .B(G8GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U441 ( .A(n382), .B(n381), .Z(n387) );
  XOR2_X1 U442 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n384) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U445 ( .A(KEYINPUT15), .B(n385), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U447 ( .A(n389), .B(n388), .Z(n392) );
  XOR2_X1 U448 ( .A(G22GAT), .B(G155GAT), .Z(n432) );
  XNOR2_X1 U449 ( .A(n390), .B(n432), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U451 ( .A(n394), .B(n393), .Z(n574) );
  INV_X1 U452 ( .A(n574), .ZN(n453) );
  NAND2_X1 U453 ( .A1(n395), .A2(n453), .ZN(n396) );
  NOR2_X1 U454 ( .A1(n552), .A2(n396), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n397), .B(KEYINPUT47), .ZN(n403) );
  XOR2_X1 U456 ( .A(KEYINPUT45), .B(KEYINPUT117), .Z(n399) );
  XNOR2_X1 U457 ( .A(KEYINPUT76), .B(n552), .ZN(n537) );
  XNOR2_X1 U458 ( .A(KEYINPUT36), .B(n537), .ZN(n576) );
  NAND2_X1 U459 ( .A1(n574), .A2(n576), .ZN(n398) );
  XNOR2_X1 U460 ( .A(n399), .B(n398), .ZN(n400) );
  NOR2_X1 U461 ( .A1(n570), .A2(n400), .ZN(n401) );
  NAND2_X1 U462 ( .A1(n401), .A2(n565), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n403), .A2(n402), .ZN(n404) );
  XNOR2_X1 U464 ( .A(KEYINPUT48), .B(n404), .ZN(n541) );
  XOR2_X1 U465 ( .A(n406), .B(n405), .Z(n408) );
  NAND2_X1 U466 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U468 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n410) );
  XNOR2_X1 U469 ( .A(G92GAT), .B(KEYINPUT94), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U471 ( .A(n412), .B(n411), .Z(n417) );
  XOR2_X1 U472 ( .A(G211GAT), .B(KEYINPUT21), .Z(n414) );
  XNOR2_X1 U473 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n438) );
  XNOR2_X1 U475 ( .A(n438), .B(n415), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U477 ( .A(n419), .B(n418), .Z(n516) );
  INV_X1 U478 ( .A(n516), .ZN(n473) );
  NAND2_X1 U479 ( .A1(n541), .A2(n473), .ZN(n422) );
  XOR2_X1 U480 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n420) );
  NOR2_X1 U481 ( .A1(n542), .A2(n423), .ZN(n564) );
  XOR2_X1 U482 ( .A(KEYINPUT91), .B(KEYINPUT85), .Z(n425) );
  XNOR2_X1 U483 ( .A(KEYINPUT22), .B(KEYINPUT90), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n426), .B(G106GAT), .Z(n429) );
  XNOR2_X1 U486 ( .A(n427), .B(G218GAT), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U488 ( .A(n431), .B(n430), .Z(n435) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n444) );
  XOR2_X1 U491 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n437) );
  XNOR2_X1 U492 ( .A(KEYINPUT23), .B(KEYINPUT87), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n442) );
  XOR2_X1 U494 ( .A(G204GAT), .B(n438), .Z(n440) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U497 ( .A(n442), .B(n441), .Z(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n461) );
  NAND2_X1 U499 ( .A1(n564), .A2(n461), .ZN(n445) );
  XOR2_X1 U500 ( .A(KEYINPUT55), .B(n445), .Z(n446) );
  NAND2_X1 U501 ( .A1(n561), .A2(n537), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n448) );
  XOR2_X1 U503 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n452) );
  XNOR2_X1 U504 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n472) );
  NOR2_X1 U506 ( .A1(n537), .A2(n453), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(KEYINPUT16), .ZN(n468) );
  XNOR2_X1 U508 ( .A(KEYINPUT27), .B(KEYINPUT97), .ZN(n455) );
  XOR2_X1 U509 ( .A(n455), .B(n516), .Z(n460) );
  XNOR2_X1 U510 ( .A(KEYINPUT64), .B(KEYINPUT28), .ZN(n456) );
  XOR2_X1 U511 ( .A(n456), .B(n461), .Z(n479) );
  INV_X1 U512 ( .A(n479), .ZN(n523) );
  NAND2_X1 U513 ( .A1(n542), .A2(n523), .ZN(n457) );
  NOR2_X1 U514 ( .A1(n460), .A2(n457), .ZN(n527) );
  NAND2_X1 U515 ( .A1(n529), .A2(n527), .ZN(n467) );
  NAND2_X1 U516 ( .A1(n476), .A2(n473), .ZN(n458) );
  NAND2_X1 U517 ( .A1(n461), .A2(n458), .ZN(n459) );
  XOR2_X1 U518 ( .A(KEYINPUT25), .B(n459), .Z(n464) );
  INV_X1 U519 ( .A(n460), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n461), .A2(n476), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U522 ( .A1(n463), .A2(n563), .ZN(n544) );
  NAND2_X1 U523 ( .A1(n464), .A2(n544), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n465), .A2(n514), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n484) );
  NAND2_X1 U526 ( .A1(n468), .A2(n484), .ZN(n469) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(n469), .Z(n502) );
  NOR2_X1 U528 ( .A1(n570), .A2(n565), .ZN(n489) );
  NAND2_X1 U529 ( .A1(n502), .A2(n489), .ZN(n470) );
  XNOR2_X1 U530 ( .A(n470), .B(KEYINPUT99), .ZN(n480) );
  NAND2_X1 U531 ( .A1(n542), .A2(n480), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U533 ( .A1(n473), .A2(n480), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT102), .ZN(n475) );
  XNOR2_X1 U535 ( .A(G8GAT), .B(n475), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U537 ( .A1(n480), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n482) );
  NAND2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n483), .ZN(G1327GAT) );
  NAND2_X1 U543 ( .A1(n576), .A2(n484), .ZN(n485) );
  NOR2_X1 U544 ( .A1(n574), .A2(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT106), .B(n488), .ZN(n512) );
  NAND2_X1 U548 ( .A1(n489), .A2(n512), .ZN(n491) );
  XOR2_X1 U549 ( .A(KEYINPUT38), .B(KEYINPUT107), .Z(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n499) );
  NOR2_X1 U551 ( .A1(n499), .A2(n514), .ZN(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT39), .B(KEYINPUT108), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n516), .A2(n499), .ZN(n495) );
  XOR2_X1 U556 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  XNOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n497) );
  NOR2_X1 U558 ( .A1(n529), .A2(n499), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n499), .A2(n523), .ZN(n500) );
  XOR2_X1 U562 ( .A(KEYINPUT110), .B(n500), .Z(n501) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  AND2_X1 U564 ( .A1(n565), .A2(n557), .ZN(n513) );
  NAND2_X1 U565 ( .A1(n513), .A2(n502), .ZN(n508) );
  NOR2_X1 U566 ( .A1(n514), .A2(n508), .ZN(n503) );
  XOR2_X1 U567 ( .A(G57GAT), .B(n503), .Z(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U569 ( .A1(n516), .A2(n508), .ZN(n505) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n529), .A2(n508), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1334GAT) );
  NOR2_X1 U574 ( .A1(n523), .A2(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n512), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n514), .A2(n522), .ZN(n515) );
  XOR2_X1 U580 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n522), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G92GAT), .B(KEYINPUT113), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n522), .ZN(n519) );
  XOR2_X1 U585 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(KEYINPUT44), .Z(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(KEYINPUT115), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n525) );
  NOR2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(n525), .B(n524), .Z(n526) );
  XNOR2_X1 U591 ( .A(KEYINPUT114), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n541), .A2(n527), .ZN(n528) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n538), .A2(n555), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT118), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U598 ( .A1(n538), .A2(n557), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U601 ( .A1(n538), .A2(n574), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n553), .A2(n555), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n545), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n549) );
  XOR2_X1 U612 ( .A(KEYINPUT52), .B(KEYINPUT120), .Z(n547) );
  NAND2_X1 U613 ( .A1(n553), .A2(n557), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT121), .Z(n551) );
  NAND2_X1 U617 ( .A1(n553), .A2(n574), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n561), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  NAND2_X1 U624 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n574), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n569) );
  NOR2_X1 U630 ( .A1(n565), .A2(n569), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n572) );
  INV_X1 U635 ( .A(n569), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n573), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

