//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n467), .A2(G137), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n466), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT70), .ZN(G160));
  AND4_X1   g054(.A1(new_n468), .A2(new_n469), .A3(new_n464), .A4(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT71), .Z(new_n482));
  NAND4_X1  g057(.A1(new_n469), .A2(new_n464), .A3(G2105), .A4(new_n466), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  AND4_X1   g067(.A1(G2105), .A2(new_n469), .A3(new_n464), .A4(new_n466), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G126), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n469), .A2(new_n464), .A3(new_n466), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n471), .A2(new_n466), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT73), .B1(new_n505), .B2(G651), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT6), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(new_n509), .B1(new_n505), .B2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT74), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT74), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XOR2_X1   g090(.A(KEYINPUT75), .B(G88), .Z(new_n516));
  NAND3_X1  g091(.A1(new_n510), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n510), .A2(G50), .A3(G543), .ZN(new_n518));
  INV_X1    g093(.A(G62), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n519), .B1(new_n513), .B2(new_n514), .ZN(new_n520));
  AND2_X1   g095(.A1(G75), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(G651), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n517), .A2(new_n518), .A3(new_n522), .A4(KEYINPUT76), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(G166));
  AND2_X1   g102(.A1(new_n510), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n506), .A2(new_n509), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n505), .A2(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(new_n515), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G89), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n536), .A2(new_n537), .B1(new_n515), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n529), .A2(new_n534), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND3_X1  g116(.A1(new_n510), .A2(G52), .A3(G543), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT77), .B(G90), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n510), .A2(new_n515), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n542), .B(new_n544), .C1(new_n508), .C2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n528), .A2(G43), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n508), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n533), .A2(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g130(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n556));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND4_X1  g134(.A1(new_n530), .A2(G53), .A3(G543), .A4(new_n531), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n510), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n510), .A2(G91), .A3(new_n515), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n513), .B2(new_n514), .ZN(new_n566));
  AND2_X1   g141(.A1(G78), .A2(G543), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n562), .A2(new_n563), .A3(new_n564), .A4(new_n568), .ZN(G299));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n546), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G77), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(new_n515), .ZN(new_n573));
  INV_X1    g148(.A(G64), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n576), .A2(KEYINPUT79), .A3(new_n544), .A4(new_n542), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n571), .A2(new_n577), .ZN(G301));
  INV_X1    g153(.A(G166), .ZN(G303));
  NAND2_X1  g154(.A1(new_n533), .A2(G87), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND3_X1  g158(.A1(new_n510), .A2(G86), .A3(new_n515), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n586), .B1(new_n513), .B2(new_n514), .ZN(new_n587));
  AND2_X1   g162(.A1(G73), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n584), .A2(new_n585), .A3(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n528), .A2(G47), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n508), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n533), .A2(G85), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n591), .A2(new_n593), .A3(KEYINPUT80), .A4(new_n594), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(G290));
  AND2_X1   g174(.A1(new_n515), .A2(G66), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT81), .ZN(new_n602));
  OAI21_X1  g177(.A(G651), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n528), .A2(G54), .ZN(new_n604));
  AND3_X1   g179(.A1(new_n510), .A2(G92), .A3(new_n515), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n605), .A2(KEYINPUT10), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n603), .B(new_n604), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  MUX2_X1   g184(.A(new_n609), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g185(.A(new_n609), .B(G301), .S(G868), .Z(G321));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G299), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(G168), .B2(new_n612), .ZN(G280));
  NAND2_X1  g190(.A1(new_n604), .A2(new_n603), .ZN(new_n616));
  INV_X1    g191(.A(new_n608), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n606), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  OR3_X1    g195(.A1(new_n609), .A2(KEYINPUT82), .A3(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT82), .B1(new_n609), .B2(G559), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  MUX2_X1   g198(.A(new_n552), .B(new_n623), .S(G868), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n499), .A2(new_n476), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n480), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n468), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT72), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n483), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n630), .B1(new_n631), .B2(new_n632), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n629), .A2(new_n637), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  AND3_X1   g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n656), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n659), .A3(new_n656), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  MUX2_X1   g255(.A(new_n680), .B(new_n679), .S(new_n672), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n683), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n682), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  AND3_X1   g266(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n686), .B2(new_n690), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  NAND3_X1  g269(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n480), .A2(G139), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n698), .B(new_n699), .C1(new_n468), .C2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G33), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G2072), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n480), .A2(G141), .ZN(new_n706));
  NAND3_X1  g281(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT26), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n709), .A2(new_n710), .B1(G105), .B2(new_n476), .ZN(new_n711));
  INV_X1    g286(.A(G129), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n706), .B(new_n711), .C1(new_n634), .C2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(G29), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n703), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(G160), .A2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G34), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(G29), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G2084), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT95), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n716), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n553), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G16), .B2(G19), .ZN(new_n727));
  INV_X1    g302(.A(G1341), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G16), .ZN(new_n730));
  NOR2_X1   g305(.A1(G171), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G5), .B2(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(G1961), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G27), .A2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G164), .B2(G29), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(G2078), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n729), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n704), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n704), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT29), .B(G2090), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n730), .A2(G21), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G168), .B2(new_n730), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n720), .A2(new_n721), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n618), .A2(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G4), .B2(G16), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n704), .B1(new_n755), .B2(G28), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n756), .A2(KEYINPUT97), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(G28), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n756), .B2(KEYINPUT97), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n754), .B1(new_n757), .B2(new_n759), .C1(new_n636), .C2(new_n704), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n733), .B2(new_n732), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n727), .A2(new_n728), .B1(G2078), .B2(new_n736), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n752), .A2(new_n750), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n714), .A2(new_n715), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n744), .A2(new_n753), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n704), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  OR2_X1    g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT90), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n480), .A2(G140), .ZN(new_n772));
  INV_X1    g347(.A(G128), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n771), .B(new_n772), .C1(new_n634), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT91), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n768), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n730), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  INV_X1    g356(.A(G299), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n730), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT98), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1956), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n716), .A2(new_n787), .A3(new_n723), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n725), .A2(new_n766), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n704), .A2(G25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n484), .A2(G119), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT85), .ZN(new_n792));
  OAI21_X1  g367(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n793));
  INV_X1    g368(.A(G107), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G2105), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n480), .B2(G131), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(new_n704), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT86), .Z(new_n799));
  XOR2_X1   g374(.A(KEYINPUT35), .B(G1991), .Z(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n798), .B(KEYINPUT86), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(new_n800), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT88), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT32), .B(G1981), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n730), .A2(G22), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT89), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G166), .B2(new_n730), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G1971), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(G1971), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n810), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n730), .A2(G23), .ZN(new_n817));
  INV_X1    g392(.A(G288), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n730), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT33), .B(G1976), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n807), .B2(new_n809), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n816), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n805), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G16), .A2(G24), .ZN(new_n827));
  XOR2_X1   g402(.A(G290), .B(KEYINPUT87), .Z(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G16), .ZN(new_n829));
  INV_X1    g404(.A(G1986), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n823), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT36), .B1(new_n826), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n834), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n802), .A2(new_n804), .B1(KEYINPUT34), .B2(new_n824), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n789), .B1(new_n835), .B2(new_n839), .ZN(G311));
  INV_X1    g415(.A(new_n789), .ZN(new_n841));
  NOR3_X1   g416(.A1(new_n826), .A2(new_n834), .A3(KEYINPUT36), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n838), .B1(new_n836), .B2(new_n837), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(G150));
  NOR2_X1   g419(.A1(new_n609), .A2(new_n619), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n528), .A2(G55), .ZN(new_n847));
  XOR2_X1   g422(.A(KEYINPUT99), .B(G93), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n533), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n849), .C1(new_n508), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n552), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n846), .B(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n854), .A2(new_n855), .A3(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n851), .A2(G860), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n856), .A2(new_n858), .ZN(G145));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  INV_X1    g435(.A(G118), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(G2105), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(new_n480), .B2(G142), .ZN(new_n863));
  INV_X1    g438(.A(G130), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n634), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT100), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n627), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n701), .B(new_n713), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n627), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n866), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n775), .A2(G164), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n775), .A2(G164), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n797), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n877), .ZN(new_n879));
  INV_X1    g454(.A(new_n797), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n875), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n870), .A2(new_n873), .A3(new_n878), .A4(new_n881), .ZN(new_n884));
  XNOR2_X1  g459(.A(G160), .B(new_n636), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G162), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n883), .B2(new_n884), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(G395));
  XNOR2_X1  g468(.A(new_n553), .B(new_n851), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n623), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n622), .A4(new_n621), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT102), .B1(new_n618), .B2(G299), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n609), .A2(new_n902), .A3(new_n782), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n618), .A2(G299), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n618), .B2(G299), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n609), .A2(new_n782), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n899), .A2(new_n900), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n899), .A2(new_n900), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n904), .A2(new_n909), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT103), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n917), .B2(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(G290), .A2(G288), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n597), .A2(new_n598), .A3(new_n818), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  XNOR2_X1  g497(.A(G166), .B(G305), .ZN(new_n923));
  OR3_X1    g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n920), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n818), .B1(new_n597), .B2(new_n598), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(KEYINPUT104), .A3(new_n920), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n923), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT42), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n924), .A2(new_n929), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n932), .ZN(new_n935));
  NAND2_X1  g510(.A1(KEYINPUT105), .A2(KEYINPUT42), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n918), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n933), .A2(new_n937), .ZN(new_n939));
  INV_X1    g514(.A(new_n911), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n940), .B(KEYINPUT103), .C1(new_n914), .C2(new_n916), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n941), .B2(new_n913), .ZN(new_n942));
  OAI21_X1  g517(.A(G868), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n851), .A2(new_n612), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(G295));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n944), .ZN(G331));
  NAND3_X1  g521(.A1(G168), .A2(new_n571), .A3(new_n577), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT106), .B1(G286), .B2(G171), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(G301), .A2(KEYINPUT106), .A3(G168), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n852), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n894), .A2(new_n949), .A3(new_n950), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(KEYINPUT107), .A3(new_n953), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n951), .A2(KEYINPUT107), .A3(new_n852), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n916), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n901), .A2(new_n903), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT41), .B1(new_n904), .B2(new_n909), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n957), .A2(new_n908), .B1(new_n958), .B2(KEYINPUT108), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n958), .A2(KEYINPUT108), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n959), .A2(new_n960), .B1(new_n953), .B2(new_n952), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n934), .B1(new_n956), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n907), .A2(new_n910), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n954), .A2(new_n955), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(new_n915), .A3(new_n953), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n930), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n966), .A3(new_n888), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n964), .A2(new_n965), .ZN(new_n970));
  AOI21_X1  g545(.A(G37), .B1(new_n970), .B2(new_n934), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT43), .B1(new_n971), .B2(new_n966), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n968), .B1(new_n971), .B2(new_n966), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(G397));
  NAND2_X1  g553(.A1(new_n776), .A2(G2067), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n775), .A2(new_n778), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n713), .B(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT109), .B(G1384), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n503), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n470), .A2(new_n475), .A3(G40), .A4(new_n477), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n983), .A2(KEYINPUT110), .A3(new_n989), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n880), .A2(new_n801), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n797), .A2(new_n800), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n993), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n989), .ZN(new_n998));
  NOR2_X1   g573(.A1(G290), .A2(G1986), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G290), .A2(G1986), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1004), .A2(KEYINPUT116), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(KEYINPUT116), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT117), .Z(new_n1007));
  AND3_X1   g582(.A1(G299), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1007), .B1(G299), .B2(new_n1005), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n499), .B2(new_n500), .ZN(new_n1012));
  INV_X1    g587(.A(new_n490), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(G114), .B2(new_n468), .ZN(new_n1014));
  INV_X1    g589(.A(G126), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n483), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1011), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(new_n988), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n1011), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1956), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n988), .B1(new_n1017), .B2(new_n986), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT45), .B(new_n984), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT56), .B(G2072), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1010), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n988), .B1(new_n1017), .B2(KEYINPUT50), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1021), .A2(KEYINPUT111), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1021), .A2(KEYINPUT111), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n750), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1017), .A2(new_n988), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n778), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n609), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1024), .A2(new_n1010), .A3(new_n1028), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1029), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n503), .A2(new_n1040), .A3(new_n1020), .A4(new_n1011), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1021), .A2(KEYINPUT111), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1348), .B1(new_n1043), .B2(new_n1030), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1036), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n618), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT60), .B1(new_n1037), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT61), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1024), .A2(new_n1010), .A3(new_n1028), .ZN(new_n1049));
  OAI211_X1 g624(.A(KEYINPUT121), .B(new_n1048), .C1(new_n1049), .C2(new_n1029), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1025), .A2(new_n981), .A3(new_n1026), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(new_n728), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1017), .B2(new_n988), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n553), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT119), .B(new_n1051), .C1(new_n1057), .C2(KEYINPUT120), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(new_n1059), .A3(new_n553), .ZN(new_n1060));
  AOI211_X1 g635(.A(KEYINPUT120), .B(new_n552), .C1(new_n1052), .C2(new_n1055), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1060), .B(KEYINPUT59), .C1(new_n1061), .C2(new_n1059), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1047), .A2(new_n1050), .A3(new_n1058), .A4(new_n1062), .ZN(new_n1063));
  OR4_X1    g638(.A1(KEYINPUT60), .A2(new_n1044), .A3(new_n609), .A4(new_n1045), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1010), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1068), .B2(new_n1038), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1069), .B2(new_n1048), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1039), .B1(new_n1063), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1017), .A2(new_n986), .ZN(new_n1072));
  INV_X1    g647(.A(G2078), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT45), .B(new_n1011), .C1(new_n1012), .C2(new_n1016), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1072), .A2(new_n1019), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT125), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT125), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1025), .A2(new_n1077), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1072), .A2(new_n1019), .A3(new_n1026), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(G2078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1033), .A2(new_n733), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1079), .A2(G301), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n988), .A2(new_n1080), .A3(G2078), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n987), .A2(new_n1026), .A3(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1083), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1084), .B(KEYINPUT54), .C1(new_n1087), .C2(new_n546), .ZN(new_n1088));
  OAI21_X1  g663(.A(G8), .B1(new_n1017), .B2(new_n988), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT112), .B(G86), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n510), .A2(new_n515), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n585), .A2(new_n1092), .A3(new_n589), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G1981), .ZN(new_n1094));
  INV_X1    g669(.A(G1981), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n584), .A2(new_n585), .A3(new_n589), .A4(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1089), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1094), .A2(KEYINPUT49), .A3(new_n1096), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n580), .A2(G1976), .A3(new_n581), .A4(new_n582), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(G8), .C1(new_n988), .C2(new_n1017), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1098), .A2(new_n1099), .B1(KEYINPUT52), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1089), .ZN(new_n1103));
  INV_X1    g678(.A(G1976), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT52), .B1(G288), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1103), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G8), .ZN(new_n1107));
  INV_X1    g682(.A(G1971), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1081), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G2090), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1030), .A2(new_n1110), .A3(new_n1021), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1107), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n525), .A2(G8), .A3(new_n526), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT55), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n525), .A2(KEYINPUT55), .A3(G8), .A4(new_n526), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1102), .B(new_n1106), .C1(new_n1112), .C2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1043), .A2(new_n1110), .A3(new_n1030), .ZN(new_n1119));
  AOI221_X4 g694(.A(new_n1107), .B1(new_n1115), .B2(new_n1116), .C1(new_n1119), .C2(new_n1109), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1088), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1123));
  INV_X1    g698(.A(G301), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1083), .A2(G301), .A3(new_n1082), .A4(new_n1086), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT54), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1071), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1121), .A2(new_n1130), .A3(new_n1124), .A4(new_n1123), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1043), .A2(new_n721), .A3(new_n1030), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1025), .A2(new_n1074), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n747), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G8), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  NAND2_X1  g713(.A1(G286), .A2(G8), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT122), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1107), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT123), .B1(new_n1143), .B2(new_n1140), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1142), .A2(KEYINPUT51), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1144), .B2(KEYINPUT51), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1132), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1144), .A2(KEYINPUT51), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1142), .A2(KEYINPUT51), .A3(new_n1144), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT124), .A4(new_n1146), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1129), .A2(new_n1131), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  AOI211_X1 g727(.A(G1976), .B(G288), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1096), .B(KEYINPUT113), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1103), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1107), .B1(new_n1119), .B2(new_n1109), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1117), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1097), .A2(new_n1090), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(new_n1103), .A3(new_n1099), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1101), .A2(KEYINPUT52), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1106), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1155), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1107), .B(G286), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1111), .ZN(new_n1164));
  AOI21_X1  g739(.A(G1971), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1165));
  OAI21_X1  g740(.A(G8), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1117), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1161), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1157), .A2(new_n1163), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT114), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT63), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1161), .B1(new_n1167), .B2(new_n1166), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1174), .A2(KEYINPUT114), .A3(new_n1157), .A4(new_n1163), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1172), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT115), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1156), .A2(new_n1117), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n1161), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1169), .B(KEYINPUT115), .C1(new_n1117), .C2(new_n1156), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1157), .A2(new_n1163), .A3(KEYINPUT63), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1162), .B1(new_n1176), .B2(new_n1183), .ZN(new_n1184));
  NOR4_X1   g759(.A1(new_n1125), .A2(new_n1118), .A3(new_n1120), .A4(new_n1130), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1148), .A2(new_n1151), .A3(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1003), .B1(new_n1152), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n979), .A2(new_n980), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n989), .B1(new_n1189), .B2(new_n713), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n989), .A2(new_n981), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT46), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1193), .A2(KEYINPUT47), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1193), .A2(KEYINPUT47), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n999), .A2(new_n989), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT48), .Z(new_n1197));
  OAI22_X1  g772(.A1(new_n1194), .A2(new_n1195), .B1(new_n997), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n998), .B1(new_n1199), .B2(new_n980), .ZN(new_n1200));
  NOR2_X1   g775(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1188), .A2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g777(.A1(new_n975), .A2(new_n976), .ZN(new_n1204));
  NOR3_X1   g778(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1205));
  OAI21_X1  g779(.A(new_n1205), .B1(new_n692), .B2(new_n693), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1206), .A2(KEYINPUT126), .ZN(new_n1207));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n1208));
  OAI211_X1 g782(.A(new_n1205), .B(new_n1208), .C1(new_n692), .C2(new_n693), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g784(.A(new_n1210), .B1(new_n889), .B2(new_n890), .ZN(new_n1211));
  NOR2_X1   g785(.A1(new_n1204), .A2(new_n1211), .ZN(G308));
  OAI221_X1 g786(.A(new_n1210), .B1(new_n890), .B2(new_n889), .C1(new_n975), .C2(new_n976), .ZN(G225));
endmodule


