

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591;

  XNOR2_X1 U320 ( .A(n400), .B(n399), .ZN(n401) );
  INV_X1 U321 ( .A(KEYINPUT92), .ZN(n399) );
  XNOR2_X1 U322 ( .A(n402), .B(n401), .ZN(n403) );
  AND2_X1 U323 ( .A1(G228GAT), .A2(G233GAT), .ZN(n288) );
  AND2_X1 U324 ( .A1(n417), .A2(n416), .ZN(n289) );
  XNOR2_X1 U325 ( .A(KEYINPUT45), .B(KEYINPUT119), .ZN(n467) );
  XNOR2_X1 U326 ( .A(n468), .B(n467), .ZN(n469) );
  INV_X1 U327 ( .A(n539), .ZN(n416) );
  XNOR2_X1 U328 ( .A(n464), .B(KEYINPUT47), .ZN(n465) );
  XNOR2_X1 U329 ( .A(n378), .B(n288), .ZN(n379) );
  XNOR2_X1 U330 ( .A(n298), .B(n406), .ZN(n299) );
  XNOR2_X1 U331 ( .A(n466), .B(n465), .ZN(n473) );
  XNOR2_X1 U332 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U333 ( .A(n300), .B(n299), .ZN(n302) );
  XNOR2_X1 U334 ( .A(n474), .B(KEYINPUT48), .ZN(n475) );
  XNOR2_X1 U335 ( .A(n387), .B(n386), .ZN(n388) );
  NOR2_X1 U336 ( .A1(n527), .A2(n479), .ZN(n576) );
  XNOR2_X1 U337 ( .A(n421), .B(KEYINPUT103), .ZN(n422) );
  XNOR2_X1 U338 ( .A(n389), .B(n388), .ZN(n480) );
  XNOR2_X1 U339 ( .A(n391), .B(n390), .ZN(n575) );
  XNOR2_X1 U340 ( .A(n306), .B(n305), .ZN(n585) );
  XOR2_X1 U341 ( .A(n332), .B(n331), .Z(n568) );
  XNOR2_X1 U342 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n490) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n459) );
  XNOR2_X1 U344 ( .A(n491), .B(n490), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n460), .B(n459), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n291) );
  XNOR2_X1 U347 ( .A(KEYINPUT79), .B(KEYINPUT15), .ZN(n290) );
  XOR2_X1 U348 ( .A(n291), .B(n290), .Z(n306) );
  XOR2_X1 U349 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n293) );
  XNOR2_X1 U350 ( .A(G71GAT), .B(G57GAT), .ZN(n292) );
  XNOR2_X1 U351 ( .A(n293), .B(n292), .ZN(n451) );
  INV_X1 U352 ( .A(KEYINPUT14), .ZN(n294) );
  XNOR2_X1 U353 ( .A(n451), .B(n294), .ZN(n296) );
  NAND2_X1 U354 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U356 ( .A(G22GAT), .B(G155GAT), .Z(n372) );
  XOR2_X1 U357 ( .A(G15GAT), .B(G127GAT), .Z(n357) );
  XOR2_X1 U358 ( .A(n372), .B(n357), .Z(n298) );
  XNOR2_X1 U359 ( .A(G8GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U360 ( .A(n297), .B(G211GAT), .ZN(n406) );
  INV_X1 U361 ( .A(G64GAT), .ZN(n301) );
  XNOR2_X1 U362 ( .A(n302), .B(n301), .ZN(n304) );
  XOR2_X1 U363 ( .A(KEYINPUT70), .B(G1GAT), .Z(n427) );
  XNOR2_X1 U364 ( .A(n427), .B(G78GAT), .ZN(n303) );
  XNOR2_X1 U365 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U366 ( .A(KEYINPUT77), .B(KEYINPUT65), .Z(n308) );
  XNOR2_X1 U367 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n307) );
  XNOR2_X1 U368 ( .A(n308), .B(n307), .ZN(n332) );
  INV_X1 U369 ( .A(G43GAT), .ZN(n309) );
  NAND2_X1 U370 ( .A1(G29GAT), .A2(n309), .ZN(n312) );
  INV_X1 U371 ( .A(G29GAT), .ZN(n310) );
  NAND2_X1 U372 ( .A1(n310), .A2(G43GAT), .ZN(n311) );
  NAND2_X1 U373 ( .A1(n312), .A2(n311), .ZN(n314) );
  XNOR2_X1 U374 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n430) );
  XNOR2_X1 U376 ( .A(G99GAT), .B(G85GAT), .ZN(n315) );
  NAND2_X1 U377 ( .A1(n315), .A2(KEYINPUT74), .ZN(n319) );
  INV_X1 U378 ( .A(n315), .ZN(n317) );
  INV_X1 U379 ( .A(KEYINPUT74), .ZN(n316) );
  NAND2_X1 U380 ( .A1(n317), .A2(n316), .ZN(n318) );
  NAND2_X1 U381 ( .A1(n319), .A2(n318), .ZN(n443) );
  XNOR2_X1 U382 ( .A(n430), .B(n443), .ZN(n324) );
  XNOR2_X1 U383 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n321) );
  AND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U386 ( .A(KEYINPUT76), .B(n322), .Z(n323) );
  XNOR2_X1 U387 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .Z(n398) );
  XOR2_X1 U389 ( .A(G92GAT), .B(n398), .Z(n326) );
  XOR2_X1 U390 ( .A(G50GAT), .B(G162GAT), .Z(n373) );
  XNOR2_X1 U391 ( .A(G106GAT), .B(n373), .ZN(n325) );
  XNOR2_X1 U392 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n330) );
  XOR2_X1 U394 ( .A(G134GAT), .B(G218GAT), .Z(n329) );
  XNOR2_X1 U395 ( .A(n330), .B(n329), .ZN(n331) );
  INV_X1 U396 ( .A(n568), .ZN(n552) );
  XNOR2_X1 U397 ( .A(KEYINPUT36), .B(n552), .ZN(n588) );
  XOR2_X1 U398 ( .A(KEYINPUT0), .B(G134GAT), .Z(n334) );
  XNOR2_X1 U399 ( .A(KEYINPUT80), .B(G120GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U401 ( .A(G113GAT), .B(n335), .Z(n369) );
  XOR2_X1 U402 ( .A(G85GAT), .B(G162GAT), .Z(n338) );
  XNOR2_X1 U403 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n336), .B(KEYINPUT2), .ZN(n385) );
  XNOR2_X1 U405 ( .A(G29GAT), .B(n385), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U407 ( .A(G127GAT), .B(n339), .ZN(n352) );
  XOR2_X1 U408 ( .A(G57GAT), .B(G155GAT), .Z(n341) );
  XNOR2_X1 U409 ( .A(G1GAT), .B(G148GAT), .ZN(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U411 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n343) );
  XNOR2_X1 U412 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n342) );
  XNOR2_X1 U413 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U414 ( .A(n345), .B(n344), .Z(n350) );
  XOR2_X1 U415 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n347) );
  NAND2_X1 U416 ( .A1(G225GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U417 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U418 ( .A(KEYINPUT89), .B(n348), .ZN(n349) );
  XNOR2_X1 U419 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n369), .B(n353), .ZN(n527) );
  XNOR2_X1 U422 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n391) );
  XOR2_X1 U423 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n355) );
  XNOR2_X1 U424 ( .A(G190GAT), .B(G71GAT), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U426 ( .A(n356), .B(G99GAT), .Z(n359) );
  XNOR2_X1 U427 ( .A(G43GAT), .B(n357), .ZN(n358) );
  XNOR2_X1 U428 ( .A(n359), .B(n358), .ZN(n365) );
  XOR2_X1 U429 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n361) );
  XNOR2_X1 U430 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n361), .B(n360), .ZN(n395) );
  XOR2_X1 U432 ( .A(G176GAT), .B(n395), .Z(n363) );
  NAND2_X1 U433 ( .A1(G227GAT), .A2(G233GAT), .ZN(n362) );
  XNOR2_X1 U434 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U435 ( .A(n365), .B(n364), .Z(n371) );
  XOR2_X1 U436 ( .A(G183GAT), .B(KEYINPUT82), .Z(n367) );
  XNOR2_X1 U437 ( .A(KEYINPUT20), .B(KEYINPUT64), .ZN(n366) );
  XNOR2_X1 U438 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n539) );
  XOR2_X1 U441 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n375) );
  XNOR2_X1 U442 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U444 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n377) );
  XNOR2_X1 U445 ( .A(G211GAT), .B(G204GAT), .ZN(n376) );
  XNOR2_X1 U446 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U447 ( .A(n381), .B(KEYINPUT86), .Z(n389) );
  XOR2_X1 U448 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n383) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G218GAT), .ZN(n382) );
  XNOR2_X1 U450 ( .A(n383), .B(n382), .ZN(n394) );
  XNOR2_X1 U451 ( .A(G106GAT), .B(G78GAT), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n384), .B(G148GAT), .ZN(n452) );
  XNOR2_X1 U453 ( .A(n394), .B(n452), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n385), .B(KEYINPUT87), .ZN(n386) );
  NOR2_X1 U455 ( .A1(n539), .A2(n480), .ZN(n390) );
  XOR2_X1 U456 ( .A(G64GAT), .B(G92GAT), .Z(n393) );
  XNOR2_X1 U457 ( .A(G176GAT), .B(G204GAT), .ZN(n392) );
  XNOR2_X1 U458 ( .A(n393), .B(n392), .ZN(n456) );
  XNOR2_X1 U459 ( .A(n394), .B(n456), .ZN(n404) );
  XOR2_X1 U460 ( .A(n395), .B(KEYINPUT91), .Z(n397) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n398), .B(KEYINPUT93), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n477) );
  XOR2_X1 U466 ( .A(KEYINPUT27), .B(n477), .Z(n415) );
  NAND2_X1 U467 ( .A1(n575), .A2(n415), .ZN(n407) );
  XNOR2_X1 U468 ( .A(KEYINPUT97), .B(n407), .ZN(n411) );
  INV_X1 U469 ( .A(n477), .ZN(n529) );
  NAND2_X1 U470 ( .A1(n539), .A2(n529), .ZN(n408) );
  NAND2_X1 U471 ( .A1(n480), .A2(n408), .ZN(n409) );
  XNOR2_X1 U472 ( .A(KEYINPUT25), .B(n409), .ZN(n410) );
  NOR2_X1 U473 ( .A1(n411), .A2(n410), .ZN(n412) );
  NOR2_X1 U474 ( .A1(n527), .A2(n412), .ZN(n413) );
  XOR2_X1 U475 ( .A(KEYINPUT98), .B(n413), .Z(n419) );
  XNOR2_X1 U476 ( .A(n480), .B(KEYINPUT67), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n414), .B(KEYINPUT28), .ZN(n533) );
  NAND2_X1 U478 ( .A1(n527), .A2(n415), .ZN(n556) );
  NOR2_X1 U479 ( .A1(n533), .A2(n556), .ZN(n538) );
  XNOR2_X1 U480 ( .A(n538), .B(KEYINPUT94), .ZN(n417) );
  XNOR2_X1 U481 ( .A(KEYINPUT95), .B(n289), .ZN(n418) );
  NAND2_X1 U482 ( .A1(n419), .A2(n418), .ZN(n494) );
  NAND2_X1 U483 ( .A1(n588), .A2(n494), .ZN(n420) );
  NOR2_X1 U484 ( .A1(n585), .A2(n420), .ZN(n423) );
  XNOR2_X1 U485 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n526) );
  XOR2_X1 U487 ( .A(G15GAT), .B(G113GAT), .Z(n425) );
  XNOR2_X1 U488 ( .A(G36GAT), .B(G50GAT), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U490 ( .A(n426), .B(G141GAT), .Z(n429) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n434) );
  XOR2_X1 U493 ( .A(n430), .B(KEYINPUT71), .Z(n432) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U496 ( .A(n434), .B(n433), .Z(n442) );
  XOR2_X1 U497 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n436) );
  XNOR2_X1 U498 ( .A(G22GAT), .B(G197GAT), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U500 ( .A(KEYINPUT72), .B(G8GAT), .Z(n438) );
  XNOR2_X1 U501 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n577) );
  INV_X1 U505 ( .A(KEYINPUT32), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n444), .B(n443), .ZN(n446) );
  NAND2_X1 U507 ( .A1(G230GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U509 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n448) );
  XNOR2_X1 U510 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n447) );
  XNOR2_X1 U511 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U512 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U514 ( .A(n454), .B(n453), .Z(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n582) );
  NOR2_X1 U516 ( .A1(n577), .A2(n582), .ZN(n495) );
  NAND2_X1 U517 ( .A1(n526), .A2(n495), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT38), .ZN(n458) );
  XNOR2_X1 U519 ( .A(KEYINPUT105), .B(n458), .ZN(n508) );
  NAND2_X1 U520 ( .A1(n508), .A2(n539), .ZN(n460) );
  XNOR2_X1 U521 ( .A(KEYINPUT41), .B(n582), .ZN(n560) );
  NOR2_X1 U522 ( .A1(n577), .A2(n560), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n461), .B(KEYINPUT46), .ZN(n462) );
  XNOR2_X1 U524 ( .A(KEYINPUT116), .B(n585), .ZN(n572) );
  NOR2_X1 U525 ( .A1(n462), .A2(n572), .ZN(n463) );
  NAND2_X1 U526 ( .A1(n463), .A2(n568), .ZN(n466) );
  XOR2_X1 U527 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n464) );
  NAND2_X1 U528 ( .A1(n588), .A2(n585), .ZN(n468) );
  NAND2_X1 U529 ( .A1(n469), .A2(n577), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n582), .A2(n470), .ZN(n471) );
  XNOR2_X1 U531 ( .A(KEYINPUT120), .B(n471), .ZN(n472) );
  NOR2_X1 U532 ( .A1(n473), .A2(n472), .ZN(n476) );
  INV_X1 U533 ( .A(KEYINPUT121), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(n537) );
  NOR2_X1 U535 ( .A1(n537), .A2(n477), .ZN(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT54), .B(n478), .Z(n479) );
  NAND2_X1 U537 ( .A1(n480), .A2(n576), .ZN(n481) );
  XNOR2_X1 U538 ( .A(n481), .B(KEYINPUT55), .ZN(n482) );
  NAND2_X1 U539 ( .A1(n482), .A2(n539), .ZN(n483) );
  XNOR2_X1 U540 ( .A(KEYINPUT126), .B(n483), .ZN(n570) );
  XOR2_X1 U541 ( .A(KEYINPUT109), .B(n560), .Z(n543) );
  NOR2_X1 U542 ( .A1(n570), .A2(n543), .ZN(n486) );
  XNOR2_X1 U543 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G176GAT), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1349GAT) );
  NAND2_X1 U546 ( .A1(n508), .A2(n527), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT39), .B(KEYINPUT106), .Z(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(G29GAT), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(G1328GAT) );
  INV_X1 U550 ( .A(n570), .ZN(n573) );
  NAND2_X1 U551 ( .A1(n573), .A2(n552), .ZN(n491) );
  XNOR2_X1 U552 ( .A(KEYINPUT100), .B(KEYINPUT34), .ZN(n500) );
  XOR2_X1 U553 ( .A(G1GAT), .B(KEYINPUT101), .Z(n498) );
  NAND2_X1 U554 ( .A1(n568), .A2(n585), .ZN(n492) );
  XOR2_X1 U555 ( .A(KEYINPUT16), .B(n492), .Z(n493) );
  AND2_X1 U556 ( .A1(n494), .A2(n493), .ZN(n512) );
  NAND2_X1 U557 ( .A1(n495), .A2(n512), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT99), .B(n496), .ZN(n505) );
  NAND2_X1 U559 ( .A1(n505), .A2(n527), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1324GAT) );
  NAND2_X1 U562 ( .A1(n505), .A2(n529), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n503) );
  NAND2_X1 U565 ( .A1(n505), .A2(n539), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G15GAT), .B(n504), .ZN(G1326GAT) );
  NAND2_X1 U568 ( .A1(n505), .A2(n533), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n529), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n507), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT107), .Z(n510) );
  NAND2_X1 U573 ( .A1(n533), .A2(n508), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(G1331GAT) );
  INV_X1 U575 ( .A(n577), .ZN(n541) );
  NOR2_X1 U576 ( .A1(n543), .A2(n541), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(KEYINPUT110), .ZN(n525) );
  AND2_X1 U578 ( .A1(n512), .A2(n525), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n527), .A2(n521), .ZN(n516) );
  XOR2_X1 U580 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n514) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1332GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n518) );
  NAND2_X1 U585 ( .A1(n521), .A2(n529), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U587 ( .A(G64GAT), .B(n519), .ZN(G1333GAT) );
  NAND2_X1 U588 ( .A1(n521), .A2(n539), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT114), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U591 ( .A1(n521), .A2(n533), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U593 ( .A(G78GAT), .B(n524), .ZN(G1335GAT) );
  AND2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n534), .A2(n527), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  XOR2_X1 U597 ( .A(G92GAT), .B(KEYINPUT115), .Z(n531) );
  NAND2_X1 U598 ( .A1(n534), .A2(n529), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n534), .A2(n539), .ZN(n532) );
  XNOR2_X1 U601 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U602 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n535), .B(KEYINPUT44), .ZN(n536) );
  XNOR2_X1 U604 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  BUF_X1 U605 ( .A(n537), .Z(n557) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U607 ( .A1(n557), .A2(n540), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n541), .A2(n553), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U610 ( .A(n553), .ZN(n544) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n548) );
  XOR2_X1 U612 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n546) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT50), .B(KEYINPUT124), .Z(n550) );
  NAND2_X1 U617 ( .A1(n553), .A2(n572), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(G127GAT), .B(n551), .Z(G1342GAT) );
  XOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n575), .A2(n558), .ZN(n567) );
  NOR2_X1 U625 ( .A1(n577), .A2(n567), .ZN(n559) );
  XOR2_X1 U626 ( .A(G141GAT), .B(n559), .Z(G1344GAT) );
  NOR2_X1 U627 ( .A1(n567), .A2(n560), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT52), .B(KEYINPUT125), .Z(n562) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1345GAT) );
  INV_X1 U632 ( .A(n585), .ZN(n565) );
  NOR2_X1 U633 ( .A1(n565), .A2(n567), .ZN(n566) );
  XOR2_X1 U634 ( .A(G155GAT), .B(n566), .Z(G1346GAT) );
  NOR2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n569), .Z(G1347GAT) );
  NOR2_X1 U637 ( .A1(n577), .A2(n570), .ZN(n571) );
  XOR2_X1 U638 ( .A(G169GAT), .B(n571), .Z(G1348GAT) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n581) );
  NOR2_X1 U642 ( .A1(n577), .A2(n581), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n581), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n589), .A2(n585), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(n590), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

