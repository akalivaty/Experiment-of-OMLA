//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT83), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G104), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT83), .A3(G107), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n194), .A2(KEYINPUT3), .A3(G104), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT3), .B1(new_n194), .B2(G104), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n195), .B(new_n197), .C1(new_n198), .C2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G101), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n196), .B2(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n194), .A2(KEYINPUT3), .A3(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G101), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n205), .A2(new_n206), .A3(new_n195), .A4(new_n197), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(KEYINPUT4), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  AOI22_X1  g028(.A1(new_n210), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n200), .A2(new_n219), .A3(G101), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n194), .A2(G104), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n196), .A2(G107), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n207), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(new_n210), .A3(new_n212), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n227), .A2(new_n210), .A3(new_n212), .A4(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT1), .B1(new_n211), .B2(G146), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n233), .A2(G128), .B1(new_n210), .B2(new_n212), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n225), .A2(new_n236), .A3(KEYINPUT10), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n221), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(KEYINPUT84), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT84), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n210), .A2(new_n240), .A3(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(G128), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n210), .A2(new_n212), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n243), .B1(new_n230), .B2(new_n231), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n207), .A2(new_n224), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT85), .B1(new_n246), .B2(KEYINPUT10), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT10), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n248), .B(new_n249), .C1(new_n244), .C2(new_n245), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n238), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G137), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT11), .A2(G134), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(G134), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G134), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G137), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G131), .ZN(new_n264));
  AOI21_X1  g078(.A(G131), .B1(new_n261), .B2(G137), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n257), .A2(new_n260), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n192), .B1(new_n251), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n242), .A2(new_n243), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n232), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n225), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n248), .B1(new_n272), .B2(new_n249), .ZN(new_n273));
  INV_X1    g087(.A(new_n250), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(KEYINPUT86), .B(new_n267), .C1(new_n275), .C2(new_n238), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n251), .A2(new_n268), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n280));
  XNOR2_X1  g094(.A(G110), .B(G140), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT82), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n283), .A2(G227), .ZN(new_n284));
  XOR2_X1   g098(.A(new_n282), .B(new_n284), .Z(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n279), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n275), .A2(new_n267), .A3(new_n238), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(new_n269), .B2(new_n276), .ZN(new_n289));
  OAI21_X1  g103(.A(KEYINPUT87), .B1(new_n289), .B2(new_n285), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n288), .A2(new_n286), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n225), .A2(new_n236), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n267), .B1(new_n292), .B2(new_n246), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n293), .B(KEYINPUT12), .Z(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n287), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G469), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n190), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n285), .B1(new_n294), .B2(new_n278), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n299), .B1(new_n277), .B2(new_n291), .ZN(new_n300));
  OAI21_X1  g114(.A(G469), .B1(new_n300), .B2(G902), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n191), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G214), .B1(G237), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G119), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT66), .A3(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(G119), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n307), .A3(G116), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G113), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n312), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n245), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G122), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(KEYINPUT8), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT89), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n316), .B1(new_n314), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n310), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT89), .A3(KEYINPUT5), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n312), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT90), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n225), .B1(new_n326), .B2(new_n327), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n319), .B(new_n321), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n234), .B1(new_n230), .B2(new_n231), .ZN(new_n331));
  OR2_X1    g145(.A1(KEYINPUT78), .A2(G125), .ZN(new_n332));
  NAND2_X1  g146(.A1(KEYINPUT78), .A2(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n218), .A2(new_n334), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT88), .B(G224), .Z(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G953), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(KEYINPUT7), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n312), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n310), .A2(new_n311), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n208), .A2(new_n344), .A3(new_n220), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n318), .A2(new_n225), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n320), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(KEYINPUT7), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n335), .A2(new_n336), .A3(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n341), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n330), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(G210), .B1(G237), .B2(G902), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n346), .ZN(new_n353));
  INV_X1    g167(.A(new_n320), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n347), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n337), .B(new_n340), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n353), .A2(new_n358), .A3(new_n354), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n351), .A2(new_n352), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n352), .B1(new_n351), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n303), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(KEYINPUT91), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(G237), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n283), .A3(G214), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(new_n211), .ZN(new_n370));
  NAND2_X1  g184(.A1(KEYINPUT18), .A2(G131), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n370), .B(new_n371), .Z(new_n372));
  XNOR2_X1  g186(.A(G125), .B(G140), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G146), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n376));
  XNOR2_X1  g190(.A(KEYINPUT76), .B(G140), .ZN(new_n377));
  INV_X1    g191(.A(G125), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n332), .A2(G140), .A3(new_n333), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(KEYINPUT76), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT77), .B(G125), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n380), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n375), .B1(new_n385), .B2(G146), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n372), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n379), .A2(new_n384), .A3(KEYINPUT16), .A4(new_n380), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT16), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n334), .A2(new_n389), .A3(new_n381), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n209), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n388), .A2(G146), .A3(new_n390), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT79), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n395), .A3(new_n209), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n370), .B(G131), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n370), .A2(G131), .ZN(new_n399));
  MUX2_X1   g213(.A(new_n398), .B(new_n399), .S(KEYINPUT17), .Z(new_n400));
  AOI21_X1  g214(.A(new_n387), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g215(.A(G113), .B(G122), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(new_n196), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n387), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n385), .A2(KEYINPUT19), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(KEYINPUT19), .B2(new_n374), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n393), .B(new_n398), .C1(new_n407), .C2(G146), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n403), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n366), .B(new_n367), .C1(new_n404), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n401), .B2(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(new_n367), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n401), .A2(new_n403), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n190), .B1(new_n404), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G475), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n283), .A2(G952), .ZN(new_n419));
  NAND2_X1  g233(.A1(G234), .A2(G237), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(G902), .A3(G953), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(G898), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G116), .B(G122), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT14), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n305), .A2(KEYINPUT14), .A3(G122), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(G107), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT92), .Z(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n194), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n211), .A2(G128), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n226), .A2(G143), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n261), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n261), .B1(new_n434), .B2(new_n435), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n427), .B(new_n194), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n435), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n434), .A2(new_n443), .ZN(new_n446));
  OAI21_X1  g260(.A(G134), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n447), .A3(new_n436), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT75), .B(G217), .Z(new_n449));
  NAND3_X1  g263(.A1(new_n189), .A2(new_n283), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n450), .ZN(new_n452));
  INV_X1    g266(.A(new_n448), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n452), .B1(new_n440), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n454), .A3(new_n190), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n455), .B(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n418), .A2(new_n426), .A3(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n302), .A2(new_n365), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT72), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g276(.A(G131), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n254), .A2(G137), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n261), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n466), .B2(new_n258), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n257), .A2(new_n260), .A3(new_n265), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n258), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n253), .A2(new_n255), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n261), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n266), .B(KEYINPUT67), .C1(new_n472), .C2(new_n463), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(new_n473), .A3(new_n236), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n217), .B1(new_n264), .B2(new_n266), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n344), .B1(new_n477), .B2(KEYINPUT71), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT71), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n461), .B(KEYINPUT28), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(KEYINPUT71), .ZN(new_n482));
  INV_X1    g296(.A(new_n344), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT28), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT72), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT68), .B1(new_n477), .B2(new_n344), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n266), .B1(new_n472), .B2(new_n463), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n331), .B1(new_n489), .B2(new_n462), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n475), .B1(new_n490), .B2(new_n473), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT68), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n492), .A3(new_n483), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n477), .A2(new_n344), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(KEYINPUT28), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n487), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n500));
  NAND3_X1  g314(.A1(new_n368), .A2(new_n283), .A3(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(G101), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n502), .B(new_n503), .Z(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT29), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n499), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n492), .B1(new_n491), .B2(new_n483), .ZN(new_n509));
  AND4_X1   g323(.A1(new_n492), .A2(new_n474), .A3(new_n476), .A4(new_n483), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n489), .A2(new_n331), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n344), .B1(new_n512), .B2(new_n475), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT28), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n483), .B1(new_n491), .B2(new_n479), .ZN(new_n517));
  INV_X1    g331(.A(new_n480), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n485), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n461), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n484), .A2(KEYINPUT72), .A3(new_n485), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n516), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT74), .B1(new_n522), .B2(new_n505), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n474), .B2(new_n476), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n512), .A2(new_n475), .A3(KEYINPUT30), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n344), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n494), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n505), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n523), .A2(new_n506), .A3(new_n529), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n522), .A2(KEYINPUT74), .A3(new_n505), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n508), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G472), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n504), .B1(new_n487), .B2(new_n516), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n494), .A2(new_n504), .A3(new_n527), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n494), .A2(KEYINPUT31), .A3(new_n504), .A4(new_n527), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT73), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n522), .A2(new_n505), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n538), .A2(new_n539), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n534), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n547), .ZN(new_n549));
  AOI211_X1 g363(.A(KEYINPUT32), .B(new_n549), .C1(new_n541), .C2(new_n545), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n533), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G234), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n449), .B1(new_n552), .B2(G902), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n226), .A2(G119), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n307), .A2(G128), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n226), .A2(KEYINPUT23), .A3(G119), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G110), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n557), .A2(new_n554), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT24), .B(G110), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n394), .A2(new_n396), .A3(new_n565), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n559), .A2(new_n560), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n564), .A2(new_n562), .ZN(new_n568));
  OAI221_X1 g382(.A(new_n393), .B1(G146), .B2(new_n374), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n187), .A2(new_n552), .A3(G953), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n570), .B(new_n571), .Z(new_n572));
  AND3_X1   g386(.A1(new_n566), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n572), .B1(new_n566), .B2(new_n569), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT25), .B1(new_n575), .B2(new_n190), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT80), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n553), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n574), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n566), .A2(new_n569), .A3(new_n572), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n190), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n575), .B(KEYINPUT81), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n553), .A2(new_n190), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n460), .A2(new_n551), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT93), .B(G101), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G3));
  AOI221_X4 g407(.A(KEYINPUT73), .B1(new_n538), .B2(new_n539), .C1(new_n522), .C2(new_n505), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n190), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n547), .B1(new_n594), .B2(new_n595), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n590), .A2(new_n302), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n303), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n351), .A2(new_n360), .ZN(new_n603));
  INV_X1    g417(.A(new_n352), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n602), .B1(new_n605), .B2(new_n361), .ZN(new_n606));
  INV_X1    g420(.A(new_n426), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n450), .A2(KEYINPUT94), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n441), .A2(new_n448), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(KEYINPUT94), .B(new_n450), .C1(new_n440), .C2(new_n453), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT33), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT95), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n609), .A2(new_n610), .A3(new_n613), .A4(KEYINPUT33), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n451), .A2(new_n454), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n456), .A2(G902), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n612), .A2(new_n614), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n455), .A2(new_n456), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n418), .A2(new_n606), .A3(new_n607), .A4(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n601), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n196), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT96), .B(KEYINPUT34), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  AOI22_X1  g440(.A1(new_n410), .A2(new_n413), .B1(new_n416), .B2(G475), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n426), .B(KEYINPUT97), .Z(new_n628));
  NAND4_X1  g442(.A1(new_n606), .A2(new_n627), .A3(new_n458), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n601), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  INV_X1    g447(.A(new_n588), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n566), .A2(new_n569), .ZN(new_n635));
  INV_X1    g449(.A(new_n572), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n578), .A2(new_n585), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n460), .A2(new_n599), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  AND2_X1   g457(.A1(new_n302), .A2(new_n640), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n551), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n421), .B(KEYINPUT99), .Z(new_n646));
  OR2_X1    g460(.A1(KEYINPUT98), .A2(G900), .ZN(new_n647));
  NAND2_X1  g461(.A1(KEYINPUT98), .A2(G900), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n424), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n627), .A2(new_n458), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n364), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XOR2_X1   g468(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n650), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n302), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT101), .Z(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n660));
  INV_X1    g474(.A(G472), .ZN(new_n661));
  INV_X1    g475(.A(new_n496), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n536), .B1(new_n662), .B2(new_n504), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n663), .B2(new_n190), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n665), .B1(new_n548), .B2(new_n550), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(new_n639), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n362), .A2(new_n363), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n418), .A2(new_n458), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n669), .A2(new_n602), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n659), .A2(new_n660), .A3(new_n667), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  AOI21_X1  g487(.A(new_n627), .B1(new_n619), .B2(new_n618), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n650), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n364), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n645), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  NAND2_X1  g492(.A1(new_n598), .A2(KEYINPUT32), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n546), .A2(new_n534), .A3(new_n547), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n679), .A2(new_n680), .B1(G472), .B2(new_n532), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n589), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n296), .A2(new_n190), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G469), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n298), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n685), .A2(new_n191), .A3(new_n621), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  INV_X1    g503(.A(new_n298), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n297), .B1(new_n296), .B2(new_n190), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n690), .A2(new_n629), .A3(new_n691), .A4(new_n191), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n682), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  INV_X1    g508(.A(new_n191), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n684), .A2(new_n695), .A3(new_n298), .A4(new_n606), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n551), .A2(new_n459), .A3(new_n640), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NOR2_X1   g513(.A1(new_n685), .A2(new_n191), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n670), .A2(new_n364), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(new_n628), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n498), .A2(new_n505), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n549), .B1(new_n703), .B2(new_n544), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n596), .B2(G472), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n700), .A2(new_n702), .A3(new_n590), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  NAND2_X1  g521(.A1(new_n418), .A2(new_n620), .ZN(new_n708));
  INV_X1    g522(.A(new_n650), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n704), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n597), .A2(new_n640), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT102), .B1(new_n712), .B2(new_n696), .ZN(new_n713));
  AOI211_X1 g527(.A(new_n639), .B(new_n704), .C1(new_n596), .C2(G472), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n697), .A3(new_n715), .A4(new_n710), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n681), .B2(new_n589), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n298), .A2(KEYINPUT103), .A3(new_n301), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT103), .B1(new_n298), .B2(new_n301), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n362), .A2(new_n363), .A3(new_n602), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n695), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n551), .A2(KEYINPUT104), .A3(new_n590), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n675), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n720), .A2(new_n725), .A3(new_n726), .A4(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(new_n551), .A3(new_n590), .A4(new_n710), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n727), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G131), .ZN(G33));
  INV_X1    g547(.A(new_n651), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n590), .A2(new_n725), .A3(new_n551), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n261), .ZN(G36));
  OR2_X1    g550(.A1(new_n300), .A2(KEYINPUT45), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n300), .A2(KEYINPUT45), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(G469), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(G469), .A2(G902), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n298), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n742), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n743), .A2(KEYINPUT106), .A3(new_n298), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n695), .A3(new_n656), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n627), .A2(new_n620), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT43), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n599), .A2(new_n639), .A3(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n759), .A2(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(KEYINPUT107), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n723), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT108), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n760), .A2(new_n764), .A3(new_n723), .A4(new_n761), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n758), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n252), .ZN(G39));
  NAND4_X1  g581(.A1(new_n681), .A2(new_n589), .A3(new_n710), .A4(new_n723), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT109), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n751), .A2(KEYINPUT47), .A3(new_n695), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT47), .B1(new_n751), .B2(new_n695), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n772), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n770), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n769), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  NAND3_X1  g594(.A1(new_n684), .A2(new_n191), .A3(new_n298), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n776), .A2(new_n770), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n755), .A2(new_n646), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(new_n590), .A3(new_n705), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n723), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT114), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n700), .A2(new_n723), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT116), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n666), .A2(new_n589), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n422), .A3(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n418), .A3(new_n620), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n784), .A2(new_n602), .A3(new_n669), .A4(new_n700), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT50), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n789), .A2(new_n783), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT117), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n798), .A3(new_n714), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n798), .B1(new_n797), .B2(new_n714), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n787), .B(new_n795), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT51), .ZN(new_n803));
  INV_X1    g617(.A(new_n801), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n799), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n781), .B(KEYINPUT115), .Z(new_n807));
  OAI21_X1  g621(.A(new_n786), .B1(new_n777), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n806), .A3(new_n795), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT52), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n713), .A2(new_n716), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n551), .B(new_n644), .C1(new_n652), .C2(new_n676), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n670), .A2(new_n191), .A3(new_n364), .A4(new_n709), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n721), .A2(new_n722), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n666), .A2(new_n815), .A3(new_n816), .A4(new_n639), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n812), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n717), .A2(KEYINPUT52), .A3(new_n814), .A4(new_n817), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n735), .B1(new_n729), .B2(new_n731), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n590), .B(new_n551), .C1(new_n686), .C2(new_n692), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n674), .A2(KEYINPUT111), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n708), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT112), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n458), .B(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n824), .B(new_n826), .C1(new_n418), .C2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n365), .A2(new_n628), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n599), .A2(new_n829), .A3(new_n600), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n823), .A2(new_n698), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n641), .A2(new_n591), .A3(new_n706), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n627), .A3(new_n650), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT113), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n723), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(KEYINPUT113), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n712), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n645), .A2(new_n839), .B1(new_n840), .B2(new_n725), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n822), .A2(new_n834), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n811), .B1(new_n821), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n645), .A2(new_n839), .ZN(new_n845));
  INV_X1    g659(.A(new_n725), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n712), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n832), .A3(new_n833), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n819), .A2(new_n820), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT53), .A4(new_n822), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n843), .A2(new_n844), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n844), .B1(new_n843), .B2(new_n850), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n720), .A2(new_n726), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n797), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT48), .Z(new_n857));
  NAND2_X1  g671(.A1(new_n784), .A2(new_n697), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n419), .B(new_n858), .C1(new_n791), .C2(new_n708), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n810), .A2(new_n853), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(G952), .B2(G953), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n669), .A2(new_n695), .A3(new_n303), .ZN(new_n863));
  AOI211_X1 g677(.A(new_n754), .B(new_n863), .C1(KEYINPUT49), .C2(new_n685), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n864), .B(new_n790), .C1(KEYINPUT49), .C2(new_n685), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n862), .A2(new_n865), .ZN(G75));
  NOR2_X1   g680(.A1(new_n283), .A2(G952), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n190), .B1(new_n843), .B2(new_n850), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n869), .B2(G210), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n356), .A2(new_n359), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n357), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n868), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT120), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n869), .A2(new_n876), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n604), .A3(new_n878), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n874), .B(KEYINPUT121), .Z(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(KEYINPUT56), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n875), .B1(new_n879), .B2(new_n881), .ZN(G51));
  NAND2_X1  g696(.A1(new_n877), .A2(new_n878), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n883), .A2(new_n741), .ZN(new_n884));
  INV_X1    g698(.A(new_n296), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT122), .B1(new_n851), .B2(new_n852), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n843), .A2(new_n850), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT54), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n742), .B(KEYINPUT57), .Z(new_n892));
  AOI21_X1  g706(.A(new_n885), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n884), .B1(new_n893), .B2(KEYINPUT123), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n895));
  INV_X1    g709(.A(new_n892), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n886), .B2(new_n890), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n897), .B2(new_n885), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n867), .B1(new_n894), .B2(new_n898), .ZN(G54));
  NAND4_X1  g713(.A1(new_n877), .A2(KEYINPUT58), .A3(G475), .A4(new_n878), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n411), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n411), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n867), .ZN(G60));
  NAND3_X1  g717(.A1(new_n612), .A2(new_n614), .A3(new_n616), .ZN(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n891), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n904), .B1(new_n853), .B2(new_n906), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n868), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n908), .A2(KEYINPUT124), .A3(new_n868), .A4(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n843), .B2(new_n850), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n867), .B1(new_n917), .B2(new_n638), .ZN(new_n918));
  INV_X1    g732(.A(new_n587), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n917), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT125), .B1(new_n917), .B2(new_n638), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(KEYINPUT61), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n920), .B(new_n922), .ZN(G66));
  OAI21_X1  g737(.A(G953), .B1(new_n338), .B2(new_n425), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n834), .B2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n871), .B1(G898), .B2(new_n283), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  NAND2_X1  g741(.A1(new_n763), .A2(new_n765), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(new_n753), .A3(new_n757), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n753), .A2(new_n701), .A3(new_n855), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n717), .A2(new_n814), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n930), .A2(new_n822), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n779), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n525), .A2(new_n526), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT126), .Z(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n407), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n933), .A2(new_n283), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n766), .B1(new_n775), .B2(new_n778), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n682), .A2(new_n723), .A3(new_n829), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n658), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n672), .A2(new_n931), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(KEYINPUT62), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(G953), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n937), .B(G900), .C1(new_n945), .C2(new_n936), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n937), .B(new_n949), .C1(new_n945), .C2(new_n936), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(G72));
  XNOR2_X1  g765(.A(new_n528), .B(KEYINPUT127), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n938), .A2(new_n834), .A3(new_n944), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT63), .Z(new_n956));
  AOI211_X1 g770(.A(new_n505), .B(new_n953), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n953), .A2(new_n505), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n938), .A2(new_n834), .A3(new_n932), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n956), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n529), .A2(new_n536), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n887), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n868), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n957), .A2(new_n960), .A3(new_n963), .ZN(G57));
endmodule


