//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT64), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G116), .ZN(new_n217));
  INV_X1    g0017(.A(G270), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT65), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n219), .A2(new_n220), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n205), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n208), .B1(new_n211), .B2(new_n213), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT13), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT67), .B(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(new_n252), .A3(G226), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(G232), .A3(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n261), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n262), .B1(G238), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n246), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n258), .A2(new_n246), .A3(new_n265), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G169), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT14), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT14), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n272), .A3(G169), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(G179), .A3(new_n275), .A4(new_n268), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n260), .A2(KEYINPUT69), .A3(G13), .A4(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT12), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n209), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n280), .B2(new_n281), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n260), .A2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G68), .A3(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n248), .A2(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G77), .ZN(new_n295));
  INV_X1    g0095(.A(G20), .ZN(new_n296));
  OAI22_X1  g0096(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(G68), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n297), .A2(KEYINPUT75), .B1(new_n215), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n297), .A2(KEYINPUT75), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n288), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT11), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n302), .A2(new_n303), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n292), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n277), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n251), .A2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(G238), .ZN(new_n309));
  INV_X1    g0109(.A(G107), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n308), .A2(new_n309), .B1(new_n310), .B2(new_n251), .ZN(new_n311));
  INV_X1    g0111(.A(new_n251), .ZN(new_n312));
  INV_X1    g0112(.A(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT67), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n312), .A2(new_n230), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n257), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n262), .B1(G244), .B2(new_n264), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n288), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(KEYINPUT70), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n293), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n298), .B1(G20), .B2(G77), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n322), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n289), .A2(G77), .A3(new_n290), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G77), .B2(new_n282), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n321), .A2(G169), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n321), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT71), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n321), .A2(new_n340), .A3(new_n337), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n334), .A2(new_n335), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n336), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G200), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n321), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n331), .A2(new_n333), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n321), .A2(G190), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n306), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n274), .A2(G190), .A3(new_n275), .A4(new_n268), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n269), .A2(G200), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n262), .B1(G226), .B2(new_n264), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n251), .A2(new_n252), .A3(G222), .ZN(new_n356));
  INV_X1    g0156(.A(G223), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n356), .B1(new_n295), .B2(new_n251), .C1(new_n308), .C2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n257), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT68), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n337), .ZN(new_n363));
  INV_X1    g0163(.A(G150), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n328), .A2(new_n294), .B1(new_n364), .B2(new_n299), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n296), .B1(new_n201), .B2(new_n215), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n288), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n289), .A2(G50), .A3(new_n290), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n367), .B(new_n368), .C1(G50), .C2(new_n282), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n363), .B(new_n369), .C1(G169), .C2(new_n362), .ZN(new_n370));
  AND4_X1   g0170(.A1(new_n307), .A2(new_n350), .A3(new_n354), .A4(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  OR3_X1    g0172(.A1(new_n362), .A2(new_n372), .A3(new_n345), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n362), .B2(new_n345), .ZN(new_n374));
  XOR2_X1   g0174(.A(new_n369), .B(KEYINPUT9), .Z(new_n375));
  AOI21_X1  g0175(.A(new_n375), .B1(new_n362), .B2(G190), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT10), .ZN(new_n378));
  INV_X1    g0178(.A(G58), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n284), .ZN(new_n380));
  OR2_X1    g0180(.A1(new_n380), .A2(new_n201), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(G20), .B1(G159), .B2(new_n298), .ZN(new_n382));
  OR2_X1    g0182(.A1(KEYINPUT76), .A2(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT76), .A2(G33), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n247), .A3(new_n384), .ZN(new_n385));
  AND3_X1   g0185(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n296), .ZN(new_n386));
  AOI21_X1  g0186(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n249), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n385), .A2(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n382), .B1(new_n390), .B2(new_n284), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n247), .B1(new_n383), .B2(new_n384), .ZN(new_n394));
  INV_X1    g0194(.A(new_n249), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n389), .A3(new_n296), .ZN(new_n397));
  AND2_X1   g0197(.A1(KEYINPUT76), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(KEYINPUT76), .A2(G33), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT3), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n249), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT7), .B1(new_n401), .B2(G20), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(G68), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n382), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n393), .B(new_n288), .C1(new_n404), .C2(new_n392), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n328), .B1(new_n260), .B2(G20), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n283), .A2(new_n328), .B1(new_n406), .B2(new_n289), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n257), .A2(new_n263), .A3(new_n230), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n409), .A2(new_n262), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n317), .A2(new_n357), .B1(new_n216), .B2(new_n313), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n411), .A2(new_n401), .B1(G33), .B2(G87), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n412), .B2(new_n360), .ZN(new_n413));
  INV_X1    g0213(.A(G169), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT77), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n410), .B(new_n337), .C1(new_n412), .C2(new_n360), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n408), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(G190), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n413), .A2(G200), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n405), .A2(new_n407), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT18), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n408), .B(new_n429), .C1(new_n419), .C2(new_n420), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n427), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n422), .A2(new_n428), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n371), .A2(new_n378), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n283), .A2(G97), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n260), .A2(G33), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n289), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(G97), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n310), .A2(G97), .ZN(new_n441));
  INV_X1    g0241(.A(G97), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G107), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(KEYINPUT6), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT6), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(KEYINPUT78), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n441), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n446), .A2(new_n451), .A3(G20), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n298), .A2(G77), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n453), .C1(new_n390), .C2(new_n310), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n454), .A2(KEYINPUT79), .A3(new_n288), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT79), .B1(new_n454), .B2(new_n288), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n440), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n251), .A2(G250), .A3(G1698), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n401), .A2(G244), .A3(new_n252), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT4), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT4), .A2(G244), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n251), .A2(new_n252), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT80), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT80), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n360), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(KEYINPUT5), .B(G41), .ZN(new_n471));
  INV_X1    g0271(.A(G45), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(G1), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n257), .A2(new_n259), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G257), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n360), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n414), .B1(new_n470), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n469), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n314), .A2(new_n316), .A3(G244), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n249), .B2(new_n400), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n459), .B(new_n458), .C1(new_n484), .C2(KEYINPUT4), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n257), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n480), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(new_n337), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n457), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n470), .B2(new_n480), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n486), .A2(KEYINPUT81), .A3(new_n487), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT82), .A4(G200), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n486), .A2(new_n487), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G190), .ZN(new_n497));
  INV_X1    g0297(.A(new_n457), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n492), .A2(G200), .A3(new_n493), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n490), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G250), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n473), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n476), .A2(new_n473), .B1(new_n360), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n217), .B1(new_n383), .B2(new_n384), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n314), .A2(new_n316), .A3(G238), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G244), .A2(G1698), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n401), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(G179), .B(new_n506), .C1(new_n511), .C2(new_n360), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n249), .A2(new_n400), .B1(new_n508), .B2(new_n509), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n257), .B1(new_n514), .B2(new_n507), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n414), .B1(new_n515), .B2(new_n506), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT83), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n401), .A2(new_n510), .ZN(new_n518));
  INV_X1    g0318(.A(new_n507), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n360), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n506), .ZN(new_n521));
  OAI21_X1  g0321(.A(G169), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n523), .A3(new_n512), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n296), .B(G68), .C1(new_n394), .C2(new_n395), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n293), .A2(G97), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n296), .B1(new_n255), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G87), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n442), .A3(new_n310), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n322), .B1(new_n525), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n282), .B1(new_n324), .B2(new_n325), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n326), .A2(new_n289), .A3(new_n437), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n517), .A2(new_n524), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n474), .A2(new_n360), .A3(G264), .ZN(new_n538));
  INV_X1    g0338(.A(G294), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n383), .B2(new_n384), .ZN(new_n540));
  NAND2_X1  g0340(.A1(G257), .A2(G1698), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n317), .B2(new_n504), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n542), .B2(new_n401), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n477), .B(new_n538), .C1(new_n543), .C2(new_n360), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n414), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT23), .B1(new_n296), .B2(G107), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT23), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(new_n310), .A3(G20), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n296), .B(G116), .C1(new_n398), .C2(new_n399), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n296), .A2(G87), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n249), .B2(new_n250), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n550), .B(new_n551), .C1(KEYINPUT22), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(KEYINPUT22), .A2(G87), .ZN(new_n555));
  AOI211_X1 g0355(.A(G20), .B(new_n555), .C1(new_n400), .C2(new_n249), .ZN(new_n556));
  OAI21_X1  g0356(.A(KEYINPUT24), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n401), .A2(KEYINPUT22), .A3(new_n296), .A4(G87), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n549), .B1(new_n507), .B2(new_n296), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n560), .A4(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n322), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n280), .A2(new_n310), .A3(new_n281), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT25), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n564), .B(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n310), .B2(new_n438), .ZN(new_n567));
  OAI221_X1 g0367(.A(new_n545), .B1(G179), .B2(new_n544), .C1(new_n563), .C2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n563), .A2(new_n567), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n544), .A2(new_n345), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G190), .B2(new_n544), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n289), .A2(G87), .A3(new_n437), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n532), .A2(new_n573), .A3(new_n533), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n520), .B2(new_n521), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n515), .A2(G190), .A3(new_n506), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n537), .A2(new_n568), .A3(new_n572), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n438), .B2(new_n217), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n289), .A2(KEYINPUT84), .A3(G116), .A4(new_n437), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n287), .A2(new_n209), .B1(G20), .B2(new_n217), .ZN(new_n583));
  AOI21_X1  g0383(.A(G20), .B1(G33), .B2(G283), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n248), .A2(G97), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT85), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT85), .B1(new_n584), .B2(new_n585), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT20), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(KEYINPUT20), .B(new_n583), .C1(new_n586), .C2(new_n587), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n217), .B2(new_n283), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(G264), .A2(G1698), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n317), .B2(new_n478), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n595), .A2(new_n401), .ZN(new_n596));
  INV_X1    g0396(.A(G303), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n251), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n257), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n479), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(G270), .B1(new_n476), .B2(new_n475), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n414), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n595), .A2(new_n401), .B1(G303), .B2(new_n312), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n360), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n477), .B1(new_n218), .B2(new_n479), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n608), .A2(new_n609), .A3(new_n337), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n593), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n593), .B(new_n602), .C1(new_n604), .C2(KEYINPUT21), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n599), .A2(G190), .A3(new_n601), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n582), .A4(new_n592), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n606), .A2(new_n611), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n578), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n435), .A2(new_n503), .A3(new_n617), .ZN(G372));
  NAND4_X1  g0418(.A1(new_n568), .A2(new_n606), .A3(new_n611), .A4(new_n612), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT87), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n522), .A2(new_n512), .B1(new_n534), .B2(new_n535), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n536), .B1(new_n513), .B2(new_n516), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n577), .A3(KEYINPUT87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n572), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n503), .A2(new_n619), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT88), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n623), .A2(new_n625), .B1(new_n489), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n457), .A2(new_n481), .A3(KEYINPUT88), .A4(new_n488), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n490), .A2(new_n577), .A3(new_n537), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n622), .B1(new_n634), .B2(KEYINPUT26), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n435), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n428), .A2(new_n431), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n339), .B(new_n341), .C1(new_n334), .C2(new_n335), .ZN(new_n639));
  INV_X1    g0439(.A(new_n343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n354), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n638), .B1(new_n642), .B2(new_n307), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n422), .A2(new_n430), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n378), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n370), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n637), .A2(new_n647), .ZN(G369));
  NAND3_X1  g0448(.A1(new_n606), .A2(new_n611), .A3(new_n612), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n260), .A2(new_n296), .A3(G13), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(KEYINPUT27), .ZN(new_n651));
  XOR2_X1   g0451(.A(new_n651), .B(KEYINPUT89), .Z(new_n652));
  INV_X1    g0452(.A(G213), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n650), .B2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n593), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n660), .A2(KEYINPUT90), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n660), .B(KEYINPUT90), .C1(new_n616), .C2(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G330), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n568), .A2(new_n572), .ZN(new_n666));
  INV_X1    g0466(.A(new_n657), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n569), .A2(new_n667), .ZN(new_n668));
  OAI22_X1  g0468(.A1(new_n666), .A2(new_n668), .B1(new_n568), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n649), .A2(new_n667), .ZN(new_n671));
  OAI22_X1  g0471(.A1(new_n671), .A2(new_n666), .B1(new_n568), .B2(new_n657), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(G399));
  INV_X1    g0474(.A(new_n206), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n530), .A2(G116), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n676), .A2(new_n678), .A3(new_n260), .ZN(new_n679));
  INV_X1    g0479(.A(new_n212), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n679), .B1(new_n680), .B2(new_n676), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT28), .Z(new_n682));
  NAND2_X1  g0482(.A1(new_n636), .A2(new_n667), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n628), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n489), .A2(new_n629), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n626), .A2(KEYINPUT26), .A3(new_n687), .A4(new_n632), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT92), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT92), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n630), .A2(new_n690), .A3(KEYINPUT26), .A4(new_n632), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n537), .A2(new_n577), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n631), .B1(new_n692), .B2(new_n489), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT93), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n634), .A2(KEYINPUT93), .A3(new_n631), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n689), .A2(new_n691), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n624), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n686), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n697), .A2(KEYINPUT94), .A3(new_n624), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n657), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT29), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n685), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n515), .A2(new_n506), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n543), .A2(new_n360), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n600), .A2(G264), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n610), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n705), .B1(new_n710), .B2(new_n495), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n706), .A2(new_n337), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n599), .B2(new_n601), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n495), .A3(new_n544), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n496), .A2(new_n709), .A3(KEYINPUT30), .A4(new_n610), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n657), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n502), .A2(new_n494), .A3(new_n497), .A4(new_n498), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n617), .A2(new_n722), .A3(new_n489), .A4(new_n667), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT91), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n503), .A2(KEYINPUT91), .A3(new_n617), .A4(new_n667), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n664), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n704), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n682), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR3_X1   g0531(.A1(new_n731), .A2(new_n472), .A3(G20), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT95), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(new_n260), .A3(new_n676), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n665), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n663), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n735), .B1(G330), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n209), .B1(G20), .B2(new_n414), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n251), .A2(new_n206), .ZN(new_n744));
  INV_X1    g0544(.A(G355), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(KEYINPUT96), .B2(new_n745), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n745), .A2(KEYINPUT96), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(new_n217), .B2(new_n675), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n241), .A2(new_n472), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n401), .A2(new_n675), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n213), .B2(G45), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n748), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n740), .B(new_n743), .C1(new_n752), .C2(KEYINPUT97), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(KEYINPUT97), .B2(new_n752), .ZN(new_n754));
  INV_X1    g0554(.A(new_n734), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n296), .A2(new_n337), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n423), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT99), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n758), .A2(KEYINPUT99), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(G326), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n296), .A2(G179), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT100), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT100), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G329), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n757), .A2(G190), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n765), .A2(new_n423), .A3(G200), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n773), .A2(new_n774), .B1(new_n776), .B2(G283), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n423), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n296), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n765), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n780), .A2(G294), .B1(new_n782), .B2(G303), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n756), .A2(new_n766), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n312), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n756), .A2(G190), .A3(new_n345), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n786), .B1(G322), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n772), .A2(new_n777), .A3(new_n783), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n767), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n793), .A2(KEYINPUT32), .B1(G107), .B2(new_n776), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n794), .B1(new_n442), .B2(new_n779), .C1(new_n762), .C2(new_n215), .ZN(new_n795));
  INV_X1    g0595(.A(new_n773), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n796), .A2(new_n284), .B1(new_n793), .B2(KEYINPUT32), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n251), .B1(new_n784), .B2(new_n295), .C1(new_n529), .C2(new_n781), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n787), .B(KEYINPUT98), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n379), .B2(new_n800), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n764), .A2(new_n790), .B1(new_n795), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n755), .B1(new_n802), .B2(new_n743), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n754), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n737), .B1(new_n742), .B2(new_n804), .ZN(G396));
  INV_X1    g0605(.A(KEYINPUT101), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n641), .A2(new_n806), .B1(new_n347), .B2(new_n667), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n347), .A2(new_n667), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n344), .A2(KEYINPUT101), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n344), .A2(new_n347), .A3(new_n346), .A4(new_n348), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n683), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n807), .A2(new_n809), .A3(new_n810), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n636), .A2(new_n813), .A3(new_n667), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n725), .A2(new_n726), .ZN(new_n816));
  INV_X1    g0616(.A(new_n721), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G330), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n734), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n819), .B2(new_n815), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n743), .A2(new_n738), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n755), .B1(new_n295), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n743), .ZN(new_n824));
  INV_X1    g0624(.A(new_n784), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n251), .B1(new_n825), .B2(G116), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n826), .B1(new_n539), .B2(new_n787), .C1(new_n770), .C2(new_n785), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n782), .A2(G107), .B1(new_n776), .B2(G87), .ZN(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n442), .B2(new_n779), .C1(new_n829), .C2(new_n796), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n827), .B(new_n830), .C1(G303), .C2(new_n763), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n773), .A2(G150), .B1(new_n825), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(G143), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n832), .B1(new_n833), .B2(new_n800), .C1(new_n762), .C2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT34), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n401), .B1(new_n215), .B2(new_n781), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n779), .A2(new_n379), .B1(new_n775), .B2(new_n284), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(new_n771), .C2(G132), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n831), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n823), .B1(new_n824), .B2(new_n840), .C1(new_n813), .C2(new_n739), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n821), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n211), .A2(new_n217), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n446), .A2(new_n451), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT35), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n846), .B2(new_n845), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT36), .ZN(new_n849));
  OR3_X1    g0649(.A1(new_n212), .A2(new_n295), .A3(new_n380), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n215), .A2(G68), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n260), .B(G13), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n288), .B1(new_n404), .B2(new_n392), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n403), .B2(new_n382), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n407), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n420), .B2(new_n419), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n426), .ZN(new_n858));
  INV_X1    g0658(.A(new_n655), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n408), .A2(new_n859), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n421), .A2(new_n862), .A3(new_n863), .A4(new_n426), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n432), .A2(new_n860), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT39), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT103), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n432), .A2(new_n408), .A3(new_n859), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n421), .A2(new_n426), .A3(new_n863), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n864), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT39), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n870), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n872), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n870), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n883), .A2(new_n878), .A3(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n869), .B2(new_n870), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT103), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n307), .A2(KEYINPUT102), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n277), .A2(new_n889), .A3(new_n306), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n887), .A2(new_n667), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n344), .A2(new_n657), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n814), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n306), .A2(new_n657), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n354), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n888), .A2(new_n890), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n354), .A2(new_n276), .A3(new_n271), .A4(new_n273), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n306), .A3(new_n657), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n903), .A2(new_n871), .B1(new_n644), .B2(new_n655), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n698), .A2(new_n699), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n628), .A3(new_n701), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n667), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n684), .B1(new_n908), .B2(KEYINPUT29), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n647), .B1(new_n909), .B2(new_n434), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n905), .B(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n901), .ZN(new_n912));
  NOR3_X1   g0712(.A1(new_n727), .A2(new_n912), .A3(new_n811), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n879), .A2(new_n870), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT40), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n917), .A3(new_n871), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n434), .A2(new_n727), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n664), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n911), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(G1), .B1(new_n731), .B2(G20), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n911), .A2(new_n922), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n853), .B1(new_n925), .B2(new_n926), .ZN(G367));
  NOR2_X1   g0727(.A1(new_n733), .A2(new_n260), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n503), .B1(new_n498), .B2(new_n667), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n490), .A2(new_n657), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n930), .A2(new_n672), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT106), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n930), .A2(new_n934), .A3(new_n672), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT44), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n933), .A2(KEYINPUT44), .A3(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n930), .A2(new_n931), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT45), .B1(new_n940), .B2(new_n673), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n940), .A2(KEYINPUT45), .A3(new_n673), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n938), .B(new_n939), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n670), .B(KEYINPUT107), .Z(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT108), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n670), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n943), .A2(KEYINPUT108), .A3(new_n944), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n671), .A2(new_n666), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n671), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n669), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n665), .B(new_n954), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n729), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n676), .B(KEYINPUT41), .Z(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n929), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n940), .A2(new_n951), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT42), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n489), .B1(new_n930), .B2(new_n568), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n667), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT105), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n624), .A2(new_n574), .A3(new_n667), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT104), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n626), .B1(new_n574), .B2(new_n667), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n964), .A2(new_n965), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n964), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n965), .B1(new_n964), .B2(new_n970), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n971), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n946), .A2(new_n940), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT109), .B1(new_n959), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n975), .B(new_n976), .Z(new_n979));
  INV_X1    g0779(.A(new_n729), .ZN(new_n980));
  INV_X1    g0780(.A(new_n949), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n981), .A2(new_n945), .A3(new_n947), .ZN(new_n982));
  INV_X1    g0782(.A(new_n955), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n928), .B1(new_n984), .B2(new_n957), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT109), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n979), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n740), .A2(new_n743), .ZN(new_n989));
  INV_X1    g0789(.A(new_n750), .ZN(new_n990));
  INV_X1    g0790(.A(new_n326), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n989), .B1(new_n990), .B2(new_n236), .C1(new_n991), .C2(new_n206), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n734), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n763), .A2(G143), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n787), .A2(new_n364), .B1(new_n767), .B2(new_n834), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n312), .B(new_n995), .C1(G50), .C2(new_n825), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G68), .A2(new_n780), .B1(new_n773), .B2(G159), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n782), .A2(G58), .B1(new_n776), .B2(G77), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n994), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n780), .A2(G107), .B1(new_n776), .B2(G97), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n539), .B2(new_n796), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n763), .B2(G311), .ZN(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n784), .A2(new_n829), .B1(new_n767), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n781), .A2(new_n217), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n401), .B(new_n1004), .C1(KEYINPUT46), .C2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1002), .B(new_n1006), .C1(new_n597), .C2(new_n800), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(KEYINPUT46), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT110), .Z(new_n1009));
  OAI21_X1  g0809(.A(new_n999), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT47), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n993), .B1(new_n1011), .B2(new_n743), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n969), .B2(new_n741), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n988), .A2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n980), .A2(new_n955), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n729), .A2(new_n983), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n1016), .A3(new_n676), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n779), .A2(new_n829), .B1(new_n781), .B2(new_n539), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n800), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1019), .A2(G317), .B1(G303), .B2(new_n825), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(KEYINPUT112), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(KEYINPUT112), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n763), .A2(G322), .B1(G311), .B2(new_n773), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT48), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1018), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT49), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n767), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n401), .B1(G326), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(new_n217), .C2(new_n775), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n796), .A2(new_n328), .B1(new_n781), .B2(new_n295), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n396), .B(new_n1033), .C1(G97), .C2(new_n776), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n763), .A2(G159), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n326), .A2(new_n780), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n787), .A2(new_n215), .B1(new_n784), .B2(new_n284), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G150), .B2(new_n1030), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n824), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n744), .A2(new_n677), .B1(G107), .B2(new_n206), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n233), .A2(new_n472), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n678), .C1(G68), .C2(G77), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n328), .A2(G50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n990), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1041), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(KEYINPUT111), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n989), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(KEYINPUT111), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n734), .B1(new_n1049), .B2(new_n1050), .C1(new_n669), .C2(new_n741), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1017), .B1(new_n955), .B2(new_n928), .C1(new_n1040), .C2(new_n1051), .ZN(G393));
  INV_X1    g0852(.A(new_n676), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1016), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n982), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n943), .B(new_n670), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1055), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n929), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n989), .B1(new_n442), .B2(new_n206), .C1(new_n990), .C2(new_n244), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n734), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT113), .Z(new_n1061));
  OAI22_X1  g0861(.A1(new_n796), .A2(new_n597), .B1(new_n775), .B2(new_n310), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n251), .B1(new_n1030), .B2(G322), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n539), .B2(new_n784), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n779), .A2(new_n217), .B1(new_n781), .B2(new_n829), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n763), .A2(G317), .B1(G311), .B2(new_n788), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT52), .ZN(new_n1068));
  AND2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT114), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n762), .A2(new_n364), .B1(new_n791), .B2(new_n787), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT51), .Z(new_n1074));
  OAI221_X1 g0874(.A(new_n401), .B1(new_n833), .B2(new_n767), .C1(new_n328), .C2(new_n784), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n779), .A2(new_n295), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G68), .B2(new_n782), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n215), .B2(new_n796), .C1(new_n529), .C2(new_n775), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1074), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1071), .A2(KEYINPUT114), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1072), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1061), .B1(new_n1081), .B2(new_n824), .C1(new_n940), .C2(new_n741), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1057), .A2(new_n1058), .A3(new_n1082), .ZN(G390));
  NAND2_X1  g0883(.A1(new_n891), .A2(new_n667), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n902), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n886), .A3(new_n882), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n907), .A2(new_n667), .A3(new_n813), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n912), .B1(new_n1087), .B2(new_n894), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n914), .A2(new_n1084), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NOR4_X1   g0890(.A1(new_n727), .A2(new_n912), .A3(new_n664), .A4(new_n811), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n728), .A2(new_n813), .A3(new_n901), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1086), .B(new_n1093), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n895), .ZN(new_n1096));
  NOR3_X1   g0896(.A1(new_n727), .A2(new_n664), .A3(new_n811), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT115), .B1(new_n1097), .B2(new_n901), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n912), .B1(new_n819), .B2(new_n811), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n901), .B1(new_n728), .B2(new_n813), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1091), .B2(KEYINPUT115), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n893), .B1(new_n702), .B2(new_n813), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1101), .A2(new_n1091), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n819), .A2(new_n434), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n646), .B(new_n1108), .C1(new_n704), .C2(new_n435), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1053), .B1(new_n1095), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT116), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1094), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1089), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n1104), .B2(new_n912), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1093), .B1(new_n1115), .B2(new_n1086), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1100), .A2(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1108), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n647), .B(new_n1119), .C1(new_n909), .C2(new_n434), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1112), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  AND4_X1   g0922(.A1(new_n1112), .A2(new_n1121), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1111), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1117), .A2(new_n929), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n822), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n734), .B1(new_n329), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n887), .A2(new_n739), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n763), .A2(G283), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n284), .A2(new_n775), .B1(new_n781), .B2(new_n529), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1076), .B(new_n1130), .C1(G107), .C2(new_n773), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n771), .A2(G294), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n312), .B1(new_n787), .B2(new_n217), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G97), .B2(new_n825), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1129), .A2(new_n1131), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT54), .B(G143), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n773), .A2(G137), .B1(new_n825), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT117), .Z(new_n1139));
  NOR2_X1   g0939(.A1(new_n775), .A2(new_n215), .ZN(new_n1140));
  INV_X1    g0940(.A(G132), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n251), .B1(new_n787), .B2(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1140), .B(new_n1142), .C1(G159), .C2(new_n780), .ZN(new_n1143));
  INV_X1    g0943(.A(G128), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1139), .B(new_n1143), .C1(new_n1144), .C2(new_n762), .ZN(new_n1145));
  OR3_X1    g0945(.A1(new_n781), .A2(KEYINPUT53), .A3(new_n364), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT53), .B1(new_n781), .B2(new_n364), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1146), .B(new_n1147), .C1(new_n770), .C2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1135), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1127), .B(new_n1128), .C1(new_n743), .C2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT118), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1124), .A2(new_n1125), .A3(new_n1152), .ZN(G378));
  INV_X1    g0953(.A(KEYINPUT57), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT116), .B1(new_n1095), .B2(new_n1110), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1121), .A2(new_n1112), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1120), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n905), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n378), .A2(new_n370), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n859), .A2(new_n369), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n919), .A2(G330), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(G330), .A3(new_n919), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1158), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1158), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1154), .B1(new_n1157), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1109), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1170), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1154), .B1(new_n1174), .B2(new_n1168), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1172), .A2(new_n1176), .A3(new_n676), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1171), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1164), .A2(new_n738), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n779), .A2(new_n284), .B1(new_n781), .B2(new_n295), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n796), .A2(new_n442), .B1(new_n775), .B2(new_n379), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n763), .C2(G116), .ZN(new_n1182));
  INV_X1    g0982(.A(G41), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n396), .B(new_n1183), .C1(new_n310), .C2(new_n787), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n771), .B2(G283), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1182), .B(new_n1185), .C1(new_n991), .C2(new_n784), .ZN(new_n1186));
  XOR2_X1   g0986(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1187));
  OR2_X1    g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1189));
  AOI21_X1  g0989(.A(G41), .B1(new_n394), .B2(G33), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1188), .B(new_n1189), .C1(G50), .C2(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n787), .A2(new_n1144), .B1(new_n784), .B2(new_n834), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G132), .B2(new_n773), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n780), .A2(G150), .B1(new_n782), .B2(new_n1137), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n762), .C2(new_n1148), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n776), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n1030), .C2(G124), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n743), .B1(new_n1191), .B2(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT120), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n755), .B(new_n1203), .C1(new_n215), .C2(new_n822), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1178), .A2(new_n929), .B1(new_n1179), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1177), .A2(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n912), .A2(new_n738), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n734), .B1(G68), .B2(new_n1126), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n762), .A2(new_n1141), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT121), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n401), .B1(new_n379), .B2(new_n775), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT122), .Z(new_n1212));
  AOI22_X1  g1012(.A1(new_n1019), .A2(G137), .B1(new_n771), .B2(G128), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G159), .A2(new_n782), .B1(new_n825), .B2(G150), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G50), .A2(new_n780), .B1(new_n773), .B2(new_n1137), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n312), .B1(new_n787), .B2(new_n829), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G107), .B2(new_n825), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1036), .B(new_n1218), .C1(new_n597), .C2(new_n770), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n773), .A2(G116), .B1(new_n776), .B2(G77), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n442), .B2(new_n781), .C1(new_n762), .C2(new_n539), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n1210), .A2(new_n1216), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1208), .B1(new_n1222), .B2(new_n743), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1107), .A2(new_n929), .B1(new_n1207), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1110), .A2(new_n958), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(G381));
  INV_X1    g1027(.A(G390), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n842), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1229), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1013), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n978), .B2(new_n987), .ZN(new_n1232));
  INV_X1    g1032(.A(G378), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1230), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1234), .A2(G375), .ZN(G407));
  NOR2_X1   g1035(.A1(new_n653), .A2(G343), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G375), .C2(new_n1237), .ZN(G409));
  INV_X1    g1038(.A(KEYINPUT125), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(G387), .B2(new_n1228), .ZN(new_n1240));
  XOR2_X1   g1040(.A(G393), .B(G396), .Z(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G387), .A2(new_n1228), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1232), .A2(G390), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1240), .A2(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G387), .A2(new_n1228), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1232), .A2(G390), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1226), .B1(KEYINPUT60), .B2(new_n1110), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1118), .A2(new_n1120), .A3(KEYINPUT60), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n676), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1224), .B1(new_n1251), .B2(new_n1253), .ZN(new_n1254));
  OR2_X1    g1054(.A1(new_n1254), .A2(new_n842), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n842), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1236), .A2(G2897), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1255), .A2(G2897), .A3(new_n1236), .A4(new_n1256), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1173), .A2(new_n1178), .A3(new_n958), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G378), .B1(new_n1205), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1264));
  OAI21_X1  g1064(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n676), .B1(new_n1157), .B2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G378), .B(new_n1205), .C1(new_n1264), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT123), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1177), .A2(KEYINPUT123), .A3(G378), .A4(new_n1205), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1263), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1261), .B1(new_n1271), .B2(new_n1236), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1271), .A2(new_n1236), .A3(new_n1257), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1250), .B(new_n1272), .C1(new_n1273), .C2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1263), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1236), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1257), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1281), .A2(KEYINPUT62), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1249), .B1(new_n1275), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1284), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1245), .A2(new_n1250), .A3(new_n1248), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1261), .B(KEYINPUT124), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1273), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1281), .A2(new_n1285), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1286), .A2(new_n1290), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1283), .A2(new_n1293), .ZN(G405));
  NAND2_X1  g1094(.A1(G375), .A2(new_n1233), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1276), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT127), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1276), .A2(new_n1298), .A3(new_n1295), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1297), .A2(new_n1249), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1249), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1257), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1249), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1297), .A2(new_n1249), .A3(new_n1299), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1280), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1302), .A2(new_n1307), .ZN(G402));
endmodule


