

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725;

  NOR2_X1 U373 ( .A1(G953), .A2(G237), .ZN(n386) );
  XOR2_X1 U374 ( .A(G134), .B(n437), .Z(n450) );
  XNOR2_X1 U375 ( .A(n551), .B(n550), .ZN(n555) );
  AND2_X1 U376 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U377 ( .A1(n615), .A2(n587), .ZN(n588) );
  OR2_X1 U378 ( .A1(n601), .A2(n586), .ZN(n447) );
  INV_X4 U379 ( .A(G128), .ZN(n356) );
  AND2_X2 U380 ( .A1(n688), .A2(n414), .ZN(n415) );
  XNOR2_X1 U381 ( .A(n562), .B(n561), .ZN(n579) );
  XNOR2_X1 U382 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U383 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U384 ( .A(n453), .B(n452), .ZN(n457) );
  AND2_X1 U385 ( .A1(n593), .A2(G953), .ZN(n691) );
  INV_X1 U386 ( .A(G119), .ZN(n403) );
  INV_X1 U387 ( .A(KEYINPUT88), .ZN(n454) );
  XNOR2_X1 U388 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n434) );
  OR2_X1 U389 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U390 ( .A(n385), .B(n384), .ZN(n500) );
  XNOR2_X1 U391 ( .A(n383), .B(G478), .ZN(n384) );
  NAND2_X1 U392 ( .A1(n581), .A2(n698), .ZN(n614) );
  XNOR2_X1 U393 ( .A(n681), .B(n680), .ZN(n682) );
  XOR2_X1 U394 ( .A(G104), .B(G107), .Z(n351) );
  NAND2_X1 U395 ( .A1(n615), .A2(n698), .ZN(n352) );
  XOR2_X1 U396 ( .A(KEYINPUT74), .B(KEYINPUT19), .Z(n353) );
  NAND2_X2 U397 ( .A1(n589), .A2(n588), .ZN(n687) );
  NAND2_X1 U398 ( .A1(n527), .A2(n526), .ZN(n711) );
  XNOR2_X2 U399 ( .A(G146), .B(G125), .ZN(n435) );
  AND2_X1 U400 ( .A1(n578), .A2(n577), .ZN(n354) );
  XOR2_X1 U401 ( .A(G101), .B(G146), .Z(n355) );
  INV_X1 U402 ( .A(KEYINPUT46), .ZN(n506) );
  INV_X1 U403 ( .A(KEYINPUT44), .ZN(n561) );
  XNOR2_X1 U404 ( .A(n451), .B(n355), .ZN(n452) );
  XNOR2_X1 U405 ( .A(n464), .B(KEYINPUT109), .ZN(n465) );
  INV_X1 U406 ( .A(KEYINPUT82), .ZN(n520) );
  XNOR2_X1 U407 ( .A(n378), .B(n377), .ZN(n379) );
  AND2_X1 U408 ( .A1(n491), .A2(n636), .ZN(n492) );
  INV_X1 U409 ( .A(n724), .ZN(n526) );
  XNOR2_X1 U410 ( .A(n380), .B(n379), .ZN(n382) );
  NOR2_X1 U411 ( .A1(n514), .A2(n476), .ZN(n469) );
  INV_X1 U412 ( .A(G953), .ZN(n432) );
  BUF_X1 U413 ( .A(n432), .Z(n712) );
  XNOR2_X1 U414 ( .A(n505), .B(KEYINPUT42), .ZN(n599) );
  XNOR2_X2 U415 ( .A(n356), .B(G143), .ZN(n376) );
  XNOR2_X1 U416 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n357) );
  XNOR2_X2 U417 ( .A(n376), .B(n357), .ZN(n437) );
  XOR2_X1 U418 ( .A(KEYINPUT5), .B(G131), .Z(n359) );
  XNOR2_X1 U419 ( .A(G137), .B(G146), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n361) );
  NAND2_X1 U421 ( .A1(n386), .A2(G210), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n366) );
  XNOR2_X1 U423 ( .A(G116), .B(G113), .ZN(n363) );
  XNOR2_X1 U424 ( .A(G101), .B(KEYINPUT69), .ZN(n362) );
  XNOR2_X1 U425 ( .A(n363), .B(n362), .ZN(n365) );
  XNOR2_X1 U426 ( .A(KEYINPUT3), .B(G119), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n443) );
  XNOR2_X1 U428 ( .A(n366), .B(n443), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n450), .B(n367), .ZN(n590) );
  NOR2_X1 U430 ( .A1(n590), .A2(G902), .ZN(n369) );
  XNOR2_X1 U431 ( .A(KEYINPUT96), .B(G472), .ZN(n368) );
  XNOR2_X2 U432 ( .A(n369), .B(n368), .ZN(n623) );
  INV_X1 U433 ( .A(KEYINPUT6), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n623), .B(n370), .ZN(n572) );
  INV_X1 U435 ( .A(G902), .ZN(n414) );
  INV_X1 U436 ( .A(G237), .ZN(n371) );
  NAND2_X1 U437 ( .A1(n414), .A2(n371), .ZN(n445) );
  NAND2_X1 U438 ( .A1(n445), .A2(G214), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n372), .B(KEYINPUT86), .ZN(n634) );
  XOR2_X1 U440 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n375) );
  AND2_X1 U441 ( .A1(G234), .A2(n432), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n373), .B(KEYINPUT8), .ZN(n401) );
  NAND2_X1 U443 ( .A1(n401), .A2(G217), .ZN(n374) );
  XNOR2_X1 U444 ( .A(n375), .B(n374), .ZN(n380) );
  XNOR2_X1 U445 ( .A(G134), .B(n376), .ZN(n378) );
  INV_X1 U446 ( .A(G107), .ZN(n377) );
  XOR2_X1 U447 ( .A(G116), .B(G122), .Z(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n683) );
  NOR2_X1 U449 ( .A1(n683), .A2(G902), .ZN(n385) );
  XNOR2_X1 U450 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n383) );
  XNOR2_X1 U451 ( .A(n435), .B(KEYINPUT10), .ZN(n410) );
  XOR2_X1 U452 ( .A(G131), .B(G140), .Z(n451) );
  XNOR2_X1 U453 ( .A(n410), .B(n451), .ZN(n710) );
  XOR2_X1 U454 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n388) );
  NAND2_X1 U455 ( .A1(G214), .A2(n386), .ZN(n387) );
  XNOR2_X1 U456 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U457 ( .A(G122), .B(G104), .Z(n390) );
  XNOR2_X1 U458 ( .A(G143), .B(G113), .ZN(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n710), .B(n393), .ZN(n609) );
  NOR2_X1 U462 ( .A1(G902), .A2(n609), .ZN(n395) );
  XNOR2_X1 U463 ( .A(KEYINPUT13), .B(KEYINPUT98), .ZN(n394) );
  XNOR2_X1 U464 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n396), .B(G475), .ZN(n499) );
  INV_X1 U466 ( .A(n499), .ZN(n470) );
  OR2_X1 U467 ( .A1(n500), .A2(n470), .ZN(n672) );
  XNOR2_X1 U468 ( .A(KEYINPUT15), .B(G902), .ZN(n582) );
  NAND2_X1 U469 ( .A1(n582), .A2(G234), .ZN(n397) );
  XNOR2_X1 U470 ( .A(n397), .B(KEYINPUT20), .ZN(n426) );
  AND2_X1 U471 ( .A1(n426), .A2(G217), .ZN(n400) );
  XNOR2_X1 U472 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n398) );
  XNOR2_X1 U473 ( .A(n398), .B(KEYINPUT25), .ZN(n399) );
  XNOR2_X1 U474 ( .A(n400), .B(n399), .ZN(n416) );
  NAND2_X1 U475 ( .A1(n401), .A2(G221), .ZN(n402) );
  XNOR2_X1 U476 ( .A(KEYINPUT67), .B(G137), .ZN(n449) );
  XNOR2_X1 U477 ( .A(n402), .B(n449), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n403), .B(G128), .ZN(n405) );
  XNOR2_X1 U479 ( .A(G110), .B(KEYINPUT24), .ZN(n404) );
  XNOR2_X1 U480 ( .A(n405), .B(n404), .ZN(n409) );
  XNOR2_X1 U481 ( .A(G140), .B(KEYINPUT89), .ZN(n407) );
  XNOR2_X1 U482 ( .A(KEYINPUT90), .B(KEYINPUT23), .ZN(n406) );
  XNOR2_X1 U483 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U484 ( .A(n409), .B(n408), .ZN(n411) );
  XNOR2_X1 U485 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U486 ( .A(n413), .B(n412), .ZN(n688) );
  XNOR2_X2 U487 ( .A(n416), .B(n415), .ZN(n617) );
  INV_X1 U488 ( .A(n617), .ZN(n558) );
  NAND2_X1 U489 ( .A1(G237), .A2(G234), .ZN(n418) );
  INV_X1 U490 ( .A(KEYINPUT14), .ZN(n417) );
  XNOR2_X1 U491 ( .A(n418), .B(n417), .ZN(n646) );
  NAND2_X1 U492 ( .A1(G953), .A2(G902), .ZN(n419) );
  NOR2_X1 U493 ( .A1(n646), .A2(n419), .ZN(n420) );
  XNOR2_X1 U494 ( .A(n420), .B(KEYINPUT105), .ZN(n421) );
  NOR2_X1 U495 ( .A1(G900), .A2(n421), .ZN(n423) );
  INV_X1 U496 ( .A(KEYINPUT106), .ZN(n422) );
  XNOR2_X1 U497 ( .A(n423), .B(n422), .ZN(n425) );
  NAND2_X1 U498 ( .A1(n712), .A2(G952), .ZN(n532) );
  OR2_X1 U499 ( .A1(n646), .A2(n532), .ZN(n424) );
  NAND2_X1 U500 ( .A1(n425), .A2(n424), .ZN(n472) );
  XOR2_X1 U501 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n428) );
  AND2_X1 U502 ( .A1(n426), .A2(G221), .ZN(n427) );
  XNOR2_X1 U503 ( .A(n428), .B(n427), .ZN(n616) );
  AND2_X1 U504 ( .A1(n472), .A2(n616), .ZN(n429) );
  NAND2_X1 U505 ( .A1(n558), .A2(n429), .ZN(n463) );
  NOR2_X1 U506 ( .A1(n672), .A2(n463), .ZN(n430) );
  NAND2_X1 U507 ( .A1(n634), .A2(n430), .ZN(n431) );
  NOR2_X1 U508 ( .A1(n572), .A2(n431), .ZN(n512) );
  NAND2_X1 U509 ( .A1(n432), .A2(G224), .ZN(n433) );
  XNOR2_X1 U510 ( .A(n434), .B(n433), .ZN(n436) );
  XNOR2_X1 U511 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U512 ( .A(n438), .B(n437), .ZN(n441) );
  XNOR2_X1 U513 ( .A(KEYINPUT72), .B(G110), .ZN(n439) );
  XNOR2_X1 U514 ( .A(n351), .B(n439), .ZN(n694) );
  INV_X1 U515 ( .A(KEYINPUT70), .ZN(n440) );
  XNOR2_X1 U516 ( .A(n694), .B(n440), .ZN(n453) );
  XNOR2_X1 U517 ( .A(n441), .B(n453), .ZN(n444) );
  XNOR2_X1 U518 ( .A(KEYINPUT16), .B(G122), .ZN(n442) );
  XNOR2_X1 U519 ( .A(n443), .B(n442), .ZN(n695) );
  XNOR2_X1 U520 ( .A(n444), .B(n695), .ZN(n601) );
  INV_X1 U521 ( .A(n582), .ZN(n586) );
  NAND2_X1 U522 ( .A1(n445), .A2(G210), .ZN(n446) );
  XNOR2_X2 U523 ( .A(n447), .B(n446), .ZN(n514) );
  INV_X1 U524 ( .A(n514), .ZN(n479) );
  NAND2_X1 U525 ( .A1(n512), .A2(n479), .ZN(n448) );
  XNOR2_X1 U526 ( .A(n448), .B(KEYINPUT36), .ZN(n461) );
  XOR2_X1 U527 ( .A(n450), .B(n449), .Z(n706) );
  NAND2_X1 U528 ( .A1(G227), .A2(n712), .ZN(n455) );
  XNOR2_X1 U529 ( .A(n706), .B(n458), .ZN(n679) );
  NOR2_X1 U530 ( .A1(n679), .A2(G902), .ZN(n460) );
  XNOR2_X1 U531 ( .A(KEYINPUT68), .B(G469), .ZN(n459) );
  XNOR2_X2 U532 ( .A(n460), .B(n459), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n474), .B(KEYINPUT1), .ZN(n621) );
  OR2_X1 U534 ( .A1(n461), .A2(n621), .ZN(n462) );
  XNOR2_X1 U535 ( .A(n462), .B(KEYINPUT113), .ZN(n719) );
  NOR2_X1 U536 ( .A1(n623), .A2(n463), .ZN(n466) );
  XNOR2_X1 U537 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n464) );
  XNOR2_X1 U538 ( .A(n466), .B(n465), .ZN(n467) );
  OR2_X2 U539 ( .A1(n474), .A2(n467), .ZN(n468) );
  XNOR2_X2 U540 ( .A(n468), .B(KEYINPUT111), .ZN(n504) );
  INV_X1 U541 ( .A(n634), .ZN(n476) );
  XNOR2_X1 U542 ( .A(n469), .B(n353), .ZN(n537) );
  AND2_X2 U543 ( .A1(n504), .A2(n537), .ZN(n668) );
  AND2_X1 U544 ( .A1(n500), .A2(n470), .ZN(n662) );
  XOR2_X1 U545 ( .A(KEYINPUT101), .B(n662), .Z(n522) );
  INV_X1 U546 ( .A(n672), .ZN(n667) );
  OR2_X1 U547 ( .A1(n522), .A2(n667), .ZN(n631) );
  NAND2_X1 U548 ( .A1(n668), .A2(n631), .ZN(n471) );
  NAND2_X1 U549 ( .A1(n471), .A2(KEYINPUT47), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n616), .B(KEYINPUT94), .ZN(n547) );
  AND2_X1 U551 ( .A1(n617), .A2(n547), .ZN(n528) );
  NAND2_X1 U552 ( .A1(n528), .A2(n472), .ZN(n473) );
  XNOR2_X1 U553 ( .A(n475), .B(KEYINPUT73), .ZN(n493) );
  OR2_X1 U554 ( .A1(n623), .A2(n476), .ZN(n478) );
  INV_X1 U555 ( .A(KEYINPUT30), .ZN(n477) );
  XNOR2_X1 U556 ( .A(n478), .B(n477), .ZN(n491) );
  AND2_X1 U557 ( .A1(n491), .A2(n479), .ZN(n480) );
  NAND2_X1 U558 ( .A1(n493), .A2(n480), .ZN(n481) );
  XOR2_X1 U559 ( .A(n481), .B(KEYINPUT108), .Z(n482) );
  AND2_X1 U560 ( .A1(n500), .A2(n499), .ZN(n542) );
  NAND2_X1 U561 ( .A1(n482), .A2(n542), .ZN(n666) );
  NAND2_X1 U562 ( .A1(n483), .A2(n666), .ZN(n485) );
  INV_X1 U563 ( .A(KEYINPUT78), .ZN(n484) );
  XNOR2_X1 U564 ( .A(n485), .B(n484), .ZN(n489) );
  XOR2_X1 U565 ( .A(KEYINPUT79), .B(n631), .Z(n569) );
  INV_X1 U566 ( .A(n569), .ZN(n486) );
  NOR2_X1 U567 ( .A1(n486), .A2(KEYINPUT47), .ZN(n487) );
  NAND2_X1 U568 ( .A1(n668), .A2(n487), .ZN(n488) );
  NAND2_X1 U569 ( .A1(n489), .A2(n488), .ZN(n490) );
  NOR2_X1 U570 ( .A1(n719), .A2(n490), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n514), .B(KEYINPUT38), .ZN(n636) );
  NAND2_X1 U572 ( .A1(n493), .A2(n492), .ZN(n496) );
  INV_X1 U573 ( .A(KEYINPUT83), .ZN(n494) );
  XNOR2_X1 U574 ( .A(n494), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U575 ( .A(n496), .B(n495), .ZN(n523) );
  NAND2_X1 U576 ( .A1(n523), .A2(n667), .ZN(n498) );
  XNOR2_X1 U577 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U578 ( .A(n498), .B(n497), .ZN(n597) );
  OR2_X1 U579 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U580 ( .A(n501), .B(KEYINPUT103), .ZN(n637) );
  AND2_X1 U581 ( .A1(n636), .A2(n634), .ZN(n502) );
  NAND2_X1 U582 ( .A1(n637), .A2(n502), .ZN(n503) );
  XNOR2_X1 U583 ( .A(n503), .B(KEYINPUT41), .ZN(n649) );
  NAND2_X1 U584 ( .A1(n504), .A2(n649), .ZN(n505) );
  NAND2_X1 U585 ( .A1(n597), .A2(n599), .ZN(n507) );
  XNOR2_X1 U586 ( .A(n507), .B(n506), .ZN(n508) );
  NAND2_X1 U587 ( .A1(n509), .A2(n508), .ZN(n511) );
  INV_X1 U588 ( .A(KEYINPUT48), .ZN(n510) );
  XNOR2_X1 U589 ( .A(n511), .B(n510), .ZN(n519) );
  NAND2_X1 U590 ( .A1(n512), .A2(n621), .ZN(n513) );
  XNOR2_X1 U591 ( .A(KEYINPUT43), .B(n513), .ZN(n515) );
  AND2_X1 U592 ( .A1(n515), .A2(n514), .ZN(n517) );
  INV_X1 U593 ( .A(KEYINPUT107), .ZN(n516) );
  XNOR2_X1 U594 ( .A(n517), .B(n516), .ZN(n723) );
  INV_X1 U595 ( .A(n723), .ZN(n518) );
  NAND2_X1 U596 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X1 U597 ( .A(n521), .B(n520), .ZN(n527) );
  NAND2_X1 U598 ( .A1(n523), .A2(n522), .ZN(n525) );
  INV_X1 U599 ( .A(KEYINPUT114), .ZN(n524) );
  XNOR2_X1 U600 ( .A(n525), .B(n524), .ZN(n724) );
  XNOR2_X1 U601 ( .A(n711), .B(KEYINPUT81), .ZN(n581) );
  INV_X1 U602 ( .A(n528), .ZN(n620) );
  OR2_X2 U603 ( .A1(n621), .A2(n620), .ZN(n563) );
  OR2_X2 U604 ( .A1(n563), .A2(n572), .ZN(n530) );
  XOR2_X1 U605 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n529) );
  XNOR2_X2 U606 ( .A(n530), .B(n529), .ZN(n648) );
  NOR2_X1 U607 ( .A1(G898), .A2(n712), .ZN(n531) );
  XOR2_X1 U608 ( .A(KEYINPUT87), .B(n531), .Z(n696) );
  NAND2_X1 U609 ( .A1(n696), .A2(G902), .ZN(n533) );
  NAND2_X1 U610 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U611 ( .A(n646), .ZN(n534) );
  AND2_X1 U612 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U613 ( .A1(n537), .A2(n536), .ZN(n539) );
  INV_X1 U614 ( .A(KEYINPUT0), .ZN(n538) );
  XNOR2_X2 U615 ( .A(n539), .B(n538), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n648), .A2(n549), .ZN(n541) );
  XNOR2_X1 U617 ( .A(KEYINPUT34), .B(KEYINPUT75), .ZN(n540) );
  XNOR2_X1 U618 ( .A(n541), .B(n540), .ZN(n543) );
  XNOR2_X1 U619 ( .A(n544), .B(KEYINPUT35), .ZN(n721) );
  NAND2_X1 U620 ( .A1(n572), .A2(n558), .ZN(n545) );
  OR2_X1 U621 ( .A1(n621), .A2(n545), .ZN(n546) );
  XNOR2_X1 U622 ( .A(n546), .B(KEYINPUT77), .ZN(n552) );
  AND2_X1 U623 ( .A1(n637), .A2(n547), .ZN(n548) );
  NAND2_X1 U624 ( .A1(n549), .A2(n548), .ZN(n551) );
  INV_X1 U625 ( .A(KEYINPUT22), .ZN(n550) );
  NAND2_X1 U626 ( .A1(n552), .A2(n555), .ZN(n554) );
  XNOR2_X1 U627 ( .A(KEYINPUT32), .B(KEYINPUT76), .ZN(n553) );
  XNOR2_X1 U628 ( .A(n554), .B(n553), .ZN(n722) );
  NAND2_X1 U629 ( .A1(n621), .A2(n555), .ZN(n574) );
  INV_X1 U630 ( .A(n574), .ZN(n556) );
  NAND2_X1 U631 ( .A1(n556), .A2(n623), .ZN(n557) );
  XNOR2_X1 U632 ( .A(n557), .B(KEYINPUT65), .ZN(n559) );
  NAND2_X1 U633 ( .A1(n559), .A2(n558), .ZN(n598) );
  AND2_X1 U634 ( .A1(n722), .A2(n598), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n721), .A2(n560), .ZN(n562) );
  NOR2_X1 U636 ( .A1(n563), .A2(n623), .ZN(n628) );
  NAND2_X1 U637 ( .A1(n628), .A2(n549), .ZN(n564) );
  XNOR2_X1 U638 ( .A(n564), .B(KEYINPUT31), .ZN(n565) );
  XNOR2_X1 U639 ( .A(KEYINPUT97), .B(n565), .ZN(n674) );
  NOR2_X1 U640 ( .A1(n474), .A2(n620), .ZN(n566) );
  NAND2_X1 U641 ( .A1(n566), .A2(n549), .ZN(n567) );
  XNOR2_X1 U642 ( .A(n567), .B(KEYINPUT95), .ZN(n568) );
  NAND2_X1 U643 ( .A1(n568), .A2(n623), .ZN(n658) );
  NAND2_X1 U644 ( .A1(n674), .A2(n658), .ZN(n570) );
  NAND2_X1 U645 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U646 ( .A(n571), .B(KEYINPUT102), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n572), .A2(n617), .ZN(n573) );
  OR2_X1 U648 ( .A1(n574), .A2(n573), .ZN(n576) );
  INV_X1 U649 ( .A(KEYINPUT104), .ZN(n575) );
  XNOR2_X1 U650 ( .A(n576), .B(n575), .ZN(n725) );
  INV_X1 U651 ( .A(n725), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n579), .A2(n354), .ZN(n580) );
  XNOR2_X2 U653 ( .A(n580), .B(KEYINPUT45), .ZN(n698) );
  XOR2_X1 U654 ( .A(KEYINPUT80), .B(n582), .Z(n583) );
  AND2_X1 U655 ( .A1(KEYINPUT2), .A2(n583), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n614), .A2(n584), .ZN(n589) );
  XOR2_X1 U657 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n585) );
  NOR2_X1 U658 ( .A1(n711), .A2(n585), .ZN(n615) );
  AND2_X2 U659 ( .A1(n698), .A2(n586), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n687), .A2(G472), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n592), .B(n591), .ZN(n594) );
  INV_X1 U663 ( .A(G952), .ZN(n593) );
  NOR2_X2 U664 ( .A1(n594), .A2(n691), .ZN(n596) );
  XNOR2_X1 U665 ( .A(KEYINPUT63), .B(KEYINPUT85), .ZN(n595) );
  XNOR2_X1 U666 ( .A(n596), .B(n595), .ZN(G57) );
  XNOR2_X1 U667 ( .A(n597), .B(G131), .ZN(G33) );
  XNOR2_X1 U668 ( .A(n598), .B(G110), .ZN(G12) );
  XNOR2_X1 U669 ( .A(n599), .B(G137), .ZN(G39) );
  NAND2_X1 U670 ( .A1(n687), .A2(G210), .ZN(n603) );
  XOR2_X1 U671 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n600) );
  XNOR2_X1 U672 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X1 U673 ( .A(n603), .B(n602), .ZN(n604) );
  NOR2_X2 U674 ( .A1(n604), .A2(n691), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n605), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U676 ( .A1(n687), .A2(G475), .ZN(n611) );
  XNOR2_X1 U677 ( .A(KEYINPUT84), .B(KEYINPUT121), .ZN(n607) );
  XNOR2_X1 U678 ( .A(KEYINPUT59), .B(KEYINPUT66), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n611), .B(n610), .ZN(n612) );
  NOR2_X2 U682 ( .A1(n612), .A2(n691), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n613), .B(KEYINPUT60), .ZN(G60) );
  AND2_X1 U684 ( .A1(n614), .A2(KEYINPUT2), .ZN(n655) );
  XOR2_X1 U685 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n619) );
  NOR2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U687 ( .A(n619), .B(n618), .Z(n626) );
  NAND2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U689 ( .A(n622), .B(KEYINPUT50), .ZN(n624) );
  NAND2_X1 U690 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U692 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U693 ( .A(KEYINPUT51), .B(n629), .ZN(n630) );
  NAND2_X1 U694 ( .A1(n630), .A2(n649), .ZN(n642) );
  NAND2_X1 U695 ( .A1(n631), .A2(n636), .ZN(n633) );
  INV_X1 U696 ( .A(n637), .ZN(n632) );
  NAND2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U698 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U699 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U700 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U701 ( .A1(n648), .A2(n640), .ZN(n641) );
  NAND2_X1 U702 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U703 ( .A(n643), .B(KEYINPUT52), .ZN(n644) );
  XNOR2_X1 U704 ( .A(n644), .B(KEYINPUT120), .ZN(n645) );
  NAND2_X1 U705 ( .A1(n645), .A2(G952), .ZN(n647) );
  NOR2_X1 U706 ( .A1(n647), .A2(n646), .ZN(n652) );
  NAND2_X1 U707 ( .A1(n648), .A2(n649), .ZN(n650) );
  NAND2_X1 U708 ( .A1(n650), .A2(n712), .ZN(n651) );
  NOR2_X1 U709 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U710 ( .A1(n352), .A2(n653), .ZN(n654) );
  NOR2_X1 U711 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U712 ( .A(n656), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U713 ( .A1(n672), .A2(n658), .ZN(n657) );
  XOR2_X1 U714 ( .A(G104), .B(n657), .Z(G6) );
  INV_X1 U715 ( .A(n662), .ZN(n675) );
  NOR2_X1 U716 ( .A1(n675), .A2(n658), .ZN(n660) );
  XNOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n659) );
  XNOR2_X1 U718 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U719 ( .A(G107), .B(n661), .ZN(G9) );
  XOR2_X1 U720 ( .A(G128), .B(KEYINPUT29), .Z(n664) );
  NAND2_X1 U721 ( .A1(n668), .A2(n662), .ZN(n663) );
  XNOR2_X1 U722 ( .A(n664), .B(n663), .ZN(G30) );
  XOR2_X1 U723 ( .A(G143), .B(KEYINPUT115), .Z(n665) );
  XNOR2_X1 U724 ( .A(n666), .B(n665), .ZN(G45) );
  XOR2_X1 U725 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n670) );
  NAND2_X1 U726 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U727 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U728 ( .A(G146), .B(n671), .ZN(G48) );
  NOR2_X1 U729 ( .A1(n672), .A2(n674), .ZN(n673) );
  XOR2_X1 U730 ( .A(G113), .B(n673), .Z(G15) );
  NOR2_X1 U731 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U732 ( .A(KEYINPUT118), .B(n676), .Z(n677) );
  XNOR2_X1 U733 ( .A(G116), .B(n677), .ZN(G18) );
  NAND2_X1 U734 ( .A1(n687), .A2(G469), .ZN(n681) );
  XOR2_X1 U735 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n678) );
  XNOR2_X1 U736 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U737 ( .A1(n691), .A2(n682), .ZN(G54) );
  NAND2_X1 U738 ( .A1(n687), .A2(G478), .ZN(n685) );
  XNOR2_X1 U739 ( .A(n683), .B(KEYINPUT122), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U741 ( .A1(n691), .A2(n686), .ZN(G63) );
  NAND2_X1 U742 ( .A1(n687), .A2(G217), .ZN(n690) );
  XNOR2_X1 U743 ( .A(n688), .B(KEYINPUT123), .ZN(n689) );
  XNOR2_X1 U744 ( .A(n690), .B(n689), .ZN(n692) );
  NOR2_X2 U745 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U746 ( .A(n693), .B(KEYINPUT124), .ZN(G66) );
  XNOR2_X1 U747 ( .A(n695), .B(n694), .ZN(n697) );
  NOR2_X1 U748 ( .A1(n697), .A2(n696), .ZN(n705) );
  NAND2_X1 U749 ( .A1(n698), .A2(n712), .ZN(n703) );
  XOR2_X1 U750 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n700) );
  NAND2_X1 U751 ( .A1(G224), .A2(G953), .ZN(n699) );
  XNOR2_X1 U752 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U753 ( .A1(n701), .A2(G898), .ZN(n702) );
  NAND2_X1 U754 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U755 ( .A(n705), .B(n704), .ZN(G69) );
  XOR2_X1 U756 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n708) );
  INV_X1 U757 ( .A(n706), .ZN(n707) );
  XNOR2_X1 U758 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X1 U759 ( .A(n710), .B(n709), .ZN(n714) );
  XOR2_X1 U760 ( .A(n711), .B(n714), .Z(n713) );
  NAND2_X1 U761 ( .A1(n713), .A2(n712), .ZN(n718) );
  XOR2_X1 U762 ( .A(G227), .B(n714), .Z(n715) );
  NAND2_X1 U763 ( .A1(n715), .A2(G900), .ZN(n716) );
  NAND2_X1 U764 ( .A1(n716), .A2(G953), .ZN(n717) );
  NAND2_X1 U765 ( .A1(n718), .A2(n717), .ZN(G72) );
  XNOR2_X1 U766 ( .A(G125), .B(n719), .ZN(n720) );
  XNOR2_X1 U767 ( .A(n720), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U768 ( .A(n721), .B(G122), .ZN(G24) );
  XNOR2_X1 U769 ( .A(G119), .B(n722), .ZN(G21) );
  XOR2_X1 U770 ( .A(G140), .B(n723), .Z(G42) );
  XOR2_X1 U771 ( .A(G134), .B(n724), .Z(G36) );
  XOR2_X1 U772 ( .A(G101), .B(n725), .Z(G3) );
endmodule

