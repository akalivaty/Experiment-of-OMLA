

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580;

  XNOR2_X1 U322 ( .A(KEYINPUT110), .B(KEYINPUT47), .ZN(n366) );
  XNOR2_X1 U323 ( .A(n352), .B(n351), .ZN(n353) );
  INV_X1 U324 ( .A(n526), .ZN(n456) );
  XNOR2_X1 U325 ( .A(n455), .B(KEYINPUT113), .ZN(n457) );
  XNOR2_X1 U326 ( .A(G15GAT), .B(G1GAT), .ZN(n292) );
  XNOR2_X1 U327 ( .A(n314), .B(G22GAT), .ZN(n315) );
  XNOR2_X1 U328 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U329 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U330 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U331 ( .A(n323), .B(n322), .ZN(n324) );
  AND2_X1 U332 ( .A1(n457), .A2(n456), .ZN(n458) );
  XOR2_X1 U333 ( .A(n361), .B(KEYINPUT41), .Z(n562) );
  XOR2_X1 U334 ( .A(n425), .B(n424), .Z(n524) );
  XNOR2_X1 U335 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U336 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U337 ( .A(n450), .B(n449), .ZN(G1352GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT124), .B(KEYINPUT122), .Z(n445) );
  XOR2_X1 U339 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n291) );
  XNOR2_X1 U340 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n290) );
  XOR2_X1 U341 ( .A(n291), .B(n290), .Z(n299) );
  XOR2_X1 U342 ( .A(G141GAT), .B(G22GAT), .Z(n429) );
  XNOR2_X1 U343 ( .A(n292), .B(KEYINPUT68), .ZN(n313) );
  XOR2_X1 U344 ( .A(n429), .B(n313), .Z(n294) );
  NAND2_X1 U345 ( .A1(G229GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U347 ( .A(G169GAT), .B(G8GAT), .Z(n376) );
  XOR2_X1 U348 ( .A(n295), .B(n376), .Z(n297) );
  XNOR2_X1 U349 ( .A(G113GAT), .B(G197GAT), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n304) );
  XOR2_X1 U352 ( .A(G29GAT), .B(KEYINPUT8), .Z(n301) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(G36GAT), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n303) );
  XOR2_X1 U355 ( .A(G50GAT), .B(KEYINPUT7), .Z(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n338) );
  XNOR2_X1 U357 ( .A(n304), .B(n338), .ZN(n504) );
  XOR2_X1 U358 ( .A(KEYINPUT70), .B(n504), .Z(n557) );
  XOR2_X1 U359 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n306) );
  XNOR2_X1 U360 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n305) );
  XOR2_X1 U361 ( .A(n306), .B(n305), .Z(n325) );
  XOR2_X1 U362 ( .A(G71GAT), .B(G127GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(G211GAT), .B(G78GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U365 ( .A(KEYINPUT76), .B(G64GAT), .Z(n310) );
  XNOR2_X1 U366 ( .A(G8GAT), .B(G183GAT), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U368 ( .A(n312), .B(n311), .Z(n318) );
  XOR2_X1 U369 ( .A(G155GAT), .B(n313), .Z(n316) );
  NAND2_X1 U370 ( .A1(G231GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n323) );
  XNOR2_X1 U372 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n319), .B(KEYINPUT71), .ZN(n351) );
  XNOR2_X1 U374 ( .A(n351), .B(KEYINPUT14), .ZN(n321) );
  INV_X1 U375 ( .A(KEYINPUT75), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n546) );
  XOR2_X1 U377 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n327) );
  XNOR2_X1 U378 ( .A(G92GAT), .B(KEYINPUT66), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n337) );
  XOR2_X1 U380 ( .A(KEYINPUT9), .B(G134GAT), .Z(n329) );
  XNOR2_X1 U381 ( .A(G162GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U383 ( .A(G99GAT), .B(G85GAT), .Z(n350) );
  XOR2_X1 U384 ( .A(KEYINPUT64), .B(n350), .Z(n331) );
  XNOR2_X1 U385 ( .A(G218GAT), .B(G190GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U387 ( .A(n333), .B(n332), .Z(n335) );
  NAND2_X1 U388 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n549) );
  XNOR2_X1 U392 ( .A(KEYINPUT36), .B(n549), .ZN(n578) );
  NOR2_X1 U393 ( .A1(n546), .A2(n578), .ZN(n340) );
  XNOR2_X1 U394 ( .A(KEYINPUT45), .B(n340), .ZN(n358) );
  XOR2_X1 U395 ( .A(KEYINPUT74), .B(G64GAT), .Z(n342) );
  XNOR2_X1 U396 ( .A(G204GAT), .B(G92GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U398 ( .A(G176GAT), .B(n343), .Z(n380) );
  XOR2_X1 U399 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n345) );
  XNOR2_X1 U400 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n380), .B(n346), .ZN(n356) );
  XNOR2_X1 U403 ( .A(G106GAT), .B(G78GAT), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n347), .B(G148GAT), .ZN(n436) );
  XNOR2_X1 U405 ( .A(n436), .B(KEYINPUT31), .ZN(n349) );
  AND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U408 ( .A(G120GAT), .B(G71GAT), .Z(n414) );
  XOR2_X1 U409 ( .A(n414), .B(n350), .Z(n352) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  INV_X1 U411 ( .A(n357), .ZN(n361) );
  NAND2_X1 U412 ( .A1(n358), .A2(n357), .ZN(n359) );
  NOR2_X1 U413 ( .A1(n557), .A2(n359), .ZN(n360) );
  XNOR2_X1 U414 ( .A(KEYINPUT111), .B(n360), .ZN(n369) );
  INV_X1 U415 ( .A(n549), .ZN(n566) );
  INV_X1 U416 ( .A(n562), .ZN(n543) );
  NOR2_X1 U417 ( .A1(n543), .A2(n504), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n362), .B(KEYINPUT46), .ZN(n363) );
  INV_X1 U419 ( .A(n546), .ZN(n573) );
  NOR2_X1 U420 ( .A1(n363), .A2(n573), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n364), .B(KEYINPUT109), .ZN(n365) );
  NOR2_X1 U422 ( .A1(n566), .A2(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n368) );
  NAND2_X1 U424 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n370), .B(KEYINPUT48), .ZN(n453) );
  XOR2_X1 U426 ( .A(G183GAT), .B(KEYINPUT84), .Z(n372) );
  XNOR2_X1 U427 ( .A(KEYINPUT85), .B(KEYINPUT18), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(n373), .B(KEYINPUT17), .Z(n375) );
  XNOR2_X1 U430 ( .A(KEYINPUT19), .B(G190GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n425) );
  XOR2_X1 U432 ( .A(n376), .B(KEYINPUT93), .Z(n378) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U435 ( .A(n379), .B(KEYINPUT92), .Z(n382) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(n380), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n425), .B(n383), .ZN(n387) );
  XOR2_X1 U439 ( .A(KEYINPUT88), .B(G218GAT), .Z(n385) );
  XNOR2_X1 U440 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(n386), .ZN(n441) );
  XNOR2_X1 U443 ( .A(n387), .B(n441), .ZN(n521) );
  NAND2_X1 U444 ( .A1(n453), .A2(n521), .ZN(n388) );
  XOR2_X1 U445 ( .A(KEYINPUT54), .B(n388), .Z(n410) );
  XOR2_X1 U446 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n390) );
  XNOR2_X1 U447 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n409) );
  XOR2_X1 U449 ( .A(G85GAT), .B(G148GAT), .Z(n392) );
  XNOR2_X1 U450 ( .A(G29GAT), .B(G141GAT), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U452 ( .A(KEYINPUT4), .B(G57GAT), .Z(n394) );
  XNOR2_X1 U453 ( .A(G1GAT), .B(G120GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U455 ( .A(n396), .B(n395), .Z(n407) );
  XNOR2_X1 U456 ( .A(G127GAT), .B(KEYINPUT81), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n397), .B(KEYINPUT0), .ZN(n398) );
  XOR2_X1 U458 ( .A(n398), .B(KEYINPUT80), .Z(n400) );
  XNOR2_X1 U459 ( .A(G113GAT), .B(G134GAT), .ZN(n399) );
  XNOR2_X1 U460 ( .A(n400), .B(n399), .ZN(n421) );
  XOR2_X1 U461 ( .A(G155GAT), .B(KEYINPUT3), .Z(n402) );
  XNOR2_X1 U462 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n401) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n437) );
  XOR2_X1 U464 ( .A(n437), .B(KEYINPUT1), .Z(n404) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n421), .B(n405), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U469 ( .A(n409), .B(n408), .Z(n519) );
  INV_X1 U470 ( .A(n519), .ZN(n474) );
  NAND2_X1 U471 ( .A1(n410), .A2(n474), .ZN(n552) );
  INV_X1 U472 ( .A(n552), .ZN(n443) );
  XOR2_X1 U473 ( .A(KEYINPUT82), .B(G176GAT), .Z(n412) );
  XNOR2_X1 U474 ( .A(G169GAT), .B(G15GAT), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U476 ( .A(n413), .B(G99GAT), .Z(n416) );
  XNOR2_X1 U477 ( .A(G43GAT), .B(n414), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U479 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n418) );
  NAND2_X1 U480 ( .A1(G227GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U482 ( .A(n420), .B(n419), .Z(n423) );
  XNOR2_X1 U483 ( .A(n421), .B(KEYINPUT65), .ZN(n422) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U485 ( .A(n524), .ZN(n556) );
  XOR2_X1 U486 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n427) );
  XNOR2_X1 U487 ( .A(G50GAT), .B(KEYINPUT24), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U489 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U492 ( .A(KEYINPUT86), .B(KEYINPUT23), .Z(n433) );
  XNOR2_X1 U493 ( .A(G204GAT), .B(KEYINPUT89), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U495 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U496 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U498 ( .A(n441), .B(n440), .Z(n553) );
  NAND2_X1 U499 ( .A1(n556), .A2(n553), .ZN(n442) );
  XOR2_X1 U500 ( .A(n442), .B(KEYINPUT26), .Z(n538) );
  NAND2_X1 U501 ( .A1(n443), .A2(n538), .ZN(n577) );
  OR2_X1 U502 ( .A1(n577), .A2(n504), .ZN(n444) );
  XNOR2_X1 U503 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U504 ( .A(n446), .B(KEYINPUT125), .Z(n450) );
  XOR2_X1 U505 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n448) );
  XNOR2_X1 U506 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n447) );
  XNOR2_X1 U507 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n451), .B(n521), .ZN(n471) );
  NAND2_X1 U509 ( .A1(n519), .A2(n471), .ZN(n452) );
  XNOR2_X1 U510 ( .A(KEYINPUT95), .B(n452), .ZN(n466) );
  NAND2_X1 U511 ( .A1(n466), .A2(n453), .ZN(n454) );
  XOR2_X1 U512 ( .A(KEYINPUT112), .B(n454), .Z(n539) );
  NAND2_X1 U513 ( .A1(n524), .A2(n539), .ZN(n455) );
  XNOR2_X1 U514 ( .A(KEYINPUT28), .B(n553), .ZN(n526) );
  XNOR2_X1 U515 ( .A(KEYINPUT114), .B(n458), .ZN(n533) );
  NAND2_X1 U516 ( .A1(n533), .A2(n562), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n460) );
  INV_X1 U518 ( .A(G120GAT), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n462), .B(n461), .ZN(G1341GAT) );
  NAND2_X1 U520 ( .A1(n573), .A2(n549), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT79), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT16), .B(n464), .ZN(n478) );
  NOR2_X1 U523 ( .A1(n526), .A2(n524), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT96), .ZN(n477) );
  AND2_X1 U526 ( .A1(n521), .A2(n524), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n553), .A2(n468), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n469) );
  XNOR2_X1 U529 ( .A(n470), .B(n469), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n471), .A2(n538), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n489) );
  NAND2_X1 U534 ( .A1(n478), .A2(n489), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n479), .B(KEYINPUT98), .ZN(n505) );
  NAND2_X1 U536 ( .A1(n557), .A2(n357), .ZN(n492) );
  NOR2_X1 U537 ( .A1(n505), .A2(n492), .ZN(n486) );
  NAND2_X1 U538 ( .A1(n486), .A2(n519), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT34), .ZN(n481) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  XOR2_X1 U541 ( .A(G8GAT), .B(KEYINPUT99), .Z(n483) );
  NAND2_X1 U542 ( .A1(n486), .A2(n521), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n524), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n486), .A2(n526), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT100), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(n488), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U551 ( .A1(n546), .A2(n489), .ZN(n490) );
  NOR2_X1 U552 ( .A1(n578), .A2(n490), .ZN(n491) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n491), .ZN(n518) );
  NOR2_X1 U554 ( .A1(n518), .A2(n492), .ZN(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(n493), .ZN(n502) );
  NAND2_X1 U556 ( .A1(n519), .A2(n502), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U558 ( .A(G29GAT), .B(n496), .Z(G1328GAT) );
  NAND2_X1 U559 ( .A1(n502), .A2(n521), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT102), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n500) );
  NAND2_X1 U563 ( .A1(n524), .A2(n502), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n502), .A2(n526), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n507) );
  NAND2_X1 U569 ( .A1(n504), .A2(n562), .ZN(n517) );
  NOR2_X1 U570 ( .A1(n505), .A2(n517), .ZN(n512) );
  NAND2_X1 U571 ( .A1(n512), .A2(n519), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  XOR2_X1 U574 ( .A(G64GAT), .B(KEYINPUT105), .Z(n510) );
  NAND2_X1 U575 ( .A1(n512), .A2(n521), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n524), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U580 ( .A1(n512), .A2(n526), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(n516) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT106), .Z(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n519), .A2(n527), .ZN(n520) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n527), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT108), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n524), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  NAND2_X1 U595 ( .A1(n533), .A2(n557), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n573), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(KEYINPUT50), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n532), .ZN(G1342GAT) );
  NAND2_X1 U600 ( .A1(n566), .A2(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT116), .Z(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1343GAT) );
  NAND2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n504), .A2(n548), .ZN(n540) );
  XOR2_X1 U607 ( .A(G141GAT), .B(n540), .Z(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n542) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n543), .A2(n548), .ZN(n544) );
  XOR2_X1 U612 ( .A(n545), .B(n544), .Z(G1345GAT) );
  NOR2_X1 U613 ( .A1(n546), .A2(n548), .ZN(n547) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n547), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1347GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n554), .B(KEYINPUT55), .ZN(n555) );
  NOR2_X1 U620 ( .A1(n556), .A2(n555), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n567), .A2(n557), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n560) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT120), .B(n561), .Z(n564) );
  NAND2_X1 U627 ( .A1(n567), .A2(n562), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n573), .A2(n567), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U632 ( .A(n568), .B(KEYINPUT58), .ZN(n569) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n571) );
  INV_X1 U635 ( .A(n577), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n574), .A2(n361), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n572), .ZN(G1353GAT) );
  XOR2_X1 U639 ( .A(G211GAT), .B(KEYINPUT127), .Z(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

