//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  INV_X1    g001(.A(G952), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(KEYINPUT96), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(KEYINPUT96), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n191), .B1(G234), .B2(G237), .ZN(new_n192));
  INV_X1    g006(.A(G902), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT70), .B(G953), .ZN(new_n194));
  AOI211_X1 g008(.A(new_n193), .B(new_n194), .C1(G234), .C2(G237), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT21), .B(G898), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G214), .B1(G237), .B2(G902), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT0), .B(G128), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n203), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n204), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT64), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n206), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G125), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n207), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(KEYINPUT1), .C1(new_n202), .C2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G128), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n220), .B(new_n211), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G128), .A3(new_n222), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n220), .B1(new_n229), .B2(new_n211), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n219), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n216), .B1(new_n231), .B2(G125), .ZN(new_n232));
  INV_X1    g046(.A(G224), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G953), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n232), .B(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT85), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n237));
  INV_X1    g051(.A(G107), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G104), .ZN(new_n239));
  INV_X1    g053(.A(G104), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G107), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n238), .A2(G104), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT80), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT80), .B(KEYINPUT3), .C1(new_n240), .C2(G107), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G101), .ZN(new_n249));
  INV_X1    g063(.A(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G116), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n255), .ZN(new_n257));
  INV_X1    g071(.A(G113), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT2), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G113), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G116), .B(G119), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n257), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n249), .A2(new_n256), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n239), .A2(new_n241), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT3), .B1(new_n240), .B2(G107), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n268), .B1(new_n271), .B2(new_n245), .ZN(new_n272));
  INV_X1    g086(.A(G101), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n272), .A2(KEYINPUT81), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n242), .B(new_n273), .C1(new_n244), .C2(new_n246), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT4), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT81), .B1(new_n272), .B2(new_n273), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n267), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n273), .B1(new_n243), .B2(new_n241), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n252), .A2(G119), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n258), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT5), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n284), .A2(new_n285), .B1(new_n263), .B2(new_n262), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n275), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n236), .B1(new_n279), .B2(new_n287), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n272), .A2(KEYINPUT4), .A3(new_n273), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n266), .A2(new_n256), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n248), .B1(new_n272), .B2(new_n273), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT81), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n247), .A2(new_n293), .A3(G101), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n278), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n287), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT85), .ZN(new_n297));
  XNOR2_X1  g111(.A(G110), .B(G122), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n288), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n296), .A2(new_n298), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(KEYINPUT6), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT86), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n291), .A2(new_n295), .ZN(new_n304));
  INV_X1    g118(.A(new_n287), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT85), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n236), .B(new_n287), .C1(new_n291), .C2(new_n295), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n298), .A2(KEYINPUT6), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n303), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND4_X1   g124(.A1(new_n303), .A2(new_n288), .A3(new_n297), .A4(new_n309), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n235), .B(new_n302), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT7), .B1(new_n233), .B2(G953), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n232), .B(new_n313), .Z(new_n314));
  NAND2_X1  g128(.A1(new_n275), .A2(new_n281), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n286), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n298), .B(KEYINPUT8), .Z(new_n317));
  INV_X1    g131(.A(new_n284), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT87), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n285), .B1(new_n284), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n264), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n280), .B1(new_n272), .B2(new_n273), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n296), .A2(new_n298), .B1(new_n316), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(G902), .B1(new_n314), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G210), .B1(G237), .B2(G902), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n312), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n312), .B2(new_n326), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n198), .B(new_n199), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n194), .A2(G227), .ZN(new_n332));
  XOR2_X1   g146(.A(G110), .B(G140), .Z(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT84), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n289), .A2(new_n215), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n275), .A2(KEYINPUT10), .A3(new_n281), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n336), .A2(new_n295), .B1(new_n231), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(G137), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(G137), .ZN(new_n342));
  INV_X1    g156(.A(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT11), .A3(G134), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G131), .ZN(new_n346));
  INV_X1    g160(.A(G131), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n341), .A2(new_n344), .A3(new_n347), .A4(new_n342), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n217), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n219), .B1(new_n352), .B2(new_n207), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n323), .B2(new_n353), .ZN(new_n354));
  AND4_X1   g168(.A1(new_n351), .A2(new_n275), .A3(new_n353), .A4(new_n281), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n338), .A2(new_n349), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n323), .A2(new_n351), .A3(new_n353), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n275), .A2(new_n353), .A3(new_n281), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT82), .ZN(new_n360));
  INV_X1    g174(.A(new_n219), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n211), .B1(new_n223), .B2(new_n224), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT67), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(new_n225), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n358), .A2(new_n360), .B1(new_n364), .B2(new_n315), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT12), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n365), .A2(new_n366), .A3(new_n349), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n315), .B(new_n219), .C1(new_n226), .C2(new_n230), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n354), .B2(new_n355), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n346), .A2(new_n348), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT12), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n335), .B(new_n357), .C1(new_n367), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n366), .B1(new_n365), .B2(new_n349), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n369), .A2(KEYINPUT12), .A3(new_n370), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n335), .B1(new_n376), .B2(new_n357), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n334), .B1(new_n373), .B2(new_n377), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n338), .A2(new_n349), .A3(new_n356), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n349), .B1(new_n338), .B2(new_n356), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n379), .A2(new_n380), .A3(new_n334), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(G469), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G469), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n193), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n334), .B1(new_n379), .B2(new_n380), .ZN(new_n386));
  INV_X1    g200(.A(new_n334), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n387), .B(new_n357), .C1(new_n367), .C2(new_n371), .ZN(new_n388));
  AOI21_X1  g202(.A(G902), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n385), .B1(new_n389), .B2(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G113), .B(G122), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(new_n240), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n187), .A2(KEYINPUT70), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G953), .ZN(new_n396));
  INV_X1    g210(.A(G237), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n394), .A2(new_n396), .A3(G214), .A4(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n202), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n194), .A2(G143), .A3(G214), .A4(new_n397), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n347), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT88), .A3(KEYINPUT18), .ZN(new_n402));
  INV_X1    g216(.A(G140), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G125), .ZN(new_n404));
  INV_X1    g218(.A(G125), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G140), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G125), .B(G140), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT78), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n411), .A3(new_n200), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n200), .B2(new_n410), .ZN(new_n413));
  NAND3_X1  g227(.A1(KEYINPUT88), .A2(KEYINPUT18), .A3(G131), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n399), .A2(new_n400), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n402), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n399), .A2(new_n400), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G131), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT17), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n399), .A2(new_n400), .A3(new_n347), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT16), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n403), .A3(G125), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n407), .B2(new_n423), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n200), .ZN(new_n426));
  OAI211_X1 g240(.A(G146), .B(new_n424), .C1(new_n407), .C2(new_n423), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(new_n418), .C2(new_n419), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n393), .B(new_n416), .C1(new_n422), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n427), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n431), .B1(KEYINPUT17), .B2(new_n401), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n421), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n393), .B1(new_n433), .B2(new_n416), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n193), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT89), .ZN(new_n436));
  OAI21_X1  g250(.A(G475), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n416), .B1(new_n422), .B2(new_n428), .ZN(new_n438));
  INV_X1    g252(.A(new_n393), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(G902), .B1(new_n440), .B2(new_n429), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT89), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT19), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n409), .A2(new_n411), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n407), .A2(KEYINPUT19), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n200), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n420), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n427), .B(new_n447), .C1(new_n448), .C2(new_n401), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n393), .B1(new_n416), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n429), .ZN(new_n452));
  NOR2_X1   g266(.A1(G475), .A2(G902), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n443), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  AOI211_X1 g269(.A(KEYINPUT20), .B(new_n455), .C1(new_n451), .C2(new_n429), .ZN(new_n456));
  OAI22_X1  g270(.A1(new_n437), .A2(new_n442), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n252), .A2(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT14), .ZN(new_n459));
  INV_X1    g273(.A(G122), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT90), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G122), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n252), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(G107), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT90), .B(G122), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n238), .B(new_n458), .C1(new_n466), .C2(new_n252), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n202), .A2(G128), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n217), .A2(G143), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n468), .A2(new_n469), .A3(new_n340), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n340), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n465), .B(new_n467), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT9), .B(G234), .ZN(new_n473));
  INV_X1    g287(.A(G217), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n473), .A2(new_n474), .A3(G953), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n217), .B2(G143), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT92), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT92), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n468), .A2(new_n479), .A3(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n202), .A2(KEYINPUT13), .A3(G128), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n478), .A2(new_n480), .A3(new_n469), .A4(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n470), .B1(new_n482), .B2(G134), .ZN(new_n483));
  INV_X1    g297(.A(new_n458), .ZN(new_n484));
  OAI21_X1  g298(.A(G107), .B1(new_n464), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT91), .A3(new_n467), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT91), .B1(new_n485), .B2(new_n467), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n472), .B(new_n475), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(new_n467), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n486), .A3(new_n483), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n475), .B1(new_n494), .B2(new_n472), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n193), .B1(new_n490), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G478), .ZN(new_n499));
  NOR2_X1   g313(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT93), .B(new_n193), .C1(new_n490), .C2(new_n495), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n496), .A2(new_n503), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT95), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n505), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n457), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(G221), .B1(new_n473), .B2(G902), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n391), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n331), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n512), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n383), .B2(new_n390), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n511), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT97), .B1(new_n518), .B2(new_n330), .ZN(new_n519));
  NOR2_X1   g333(.A1(G472), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT31), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT65), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n209), .B1(new_n207), .B2(new_n208), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n211), .A2(new_n213), .A3(KEYINPUT64), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND4_X1   g340(.A1(new_n523), .A2(new_n526), .A3(new_n370), .A4(new_n206), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n205), .B1(new_n524), .B2(new_n525), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n523), .B1(new_n528), .B2(new_n370), .ZN(new_n529));
  INV_X1    g343(.A(new_n342), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n340), .A2(G137), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n348), .ZN(new_n533));
  OAI22_X1  g347(.A1(new_n527), .A2(new_n529), .B1(new_n364), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n290), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT69), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n526), .A2(new_n370), .A3(new_n206), .ZN(new_n538));
  INV_X1    g352(.A(new_n533), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n231), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n540), .B2(KEYINPUT30), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n528), .A2(new_n370), .ZN(new_n542));
  OAI211_X1 g356(.A(KEYINPUT30), .B(new_n542), .C1(new_n364), .C2(new_n533), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(KEYINPUT69), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n536), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n290), .B(new_n542), .C1(new_n364), .C2(new_n533), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n194), .A2(G210), .A3(new_n397), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(G101), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n522), .B1(new_n545), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(KEYINPUT69), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n231), .A2(new_n539), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(new_n537), .A3(KEYINPUT30), .A4(new_n542), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI211_X1 g372(.A(KEYINPUT31), .B(new_n552), .C1(new_n558), .C2(new_n536), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n551), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT65), .B1(new_n215), .B2(new_n349), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n528), .A2(new_n523), .A3(new_n370), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n290), .B1(new_n565), .B2(new_n556), .ZN(new_n566));
  INV_X1    g380(.A(new_n546), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT28), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT28), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n546), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n562), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n290), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n534), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n569), .B1(new_n573), .B2(new_n546), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT72), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n561), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n521), .B1(new_n560), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n578));
  OAI21_X1  g392(.A(KEYINPUT74), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n545), .A2(new_n553), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT31), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n545), .A2(new_n522), .A3(new_n553), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n570), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT72), .B1(new_n574), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n568), .A2(new_n562), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n551), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n520), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n589));
  INV_X1    g403(.A(new_n578), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n579), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n551), .B1(new_n571), .B2(new_n575), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n567), .B1(new_n558), .B2(new_n536), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n561), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT29), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n540), .B(new_n290), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n584), .B1(new_n597), .B2(KEYINPUT28), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT29), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n561), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n596), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n560), .A2(new_n576), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT32), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n521), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n607), .ZN(new_n609));
  AOI211_X1 g423(.A(KEYINPUT75), .B(new_n609), .C1(new_n560), .C2(new_n576), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n592), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n474), .B1(G234), .B2(new_n193), .ZN(new_n613));
  INV_X1    g427(.A(new_n194), .ZN(new_n614));
  NAND2_X1  g428(.A1(G221), .A2(G234), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT79), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT79), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n194), .A2(new_n617), .A3(G221), .A4(G234), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT22), .B(G137), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n616), .B2(new_n618), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT76), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n250), .B2(G128), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n217), .A2(KEYINPUT76), .A3(G119), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n250), .A2(G128), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT24), .B(G110), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n250), .A2(G128), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n626), .B(new_n630), .C1(new_n631), .C2(KEYINPUT23), .ZN(new_n632));
  OAI22_X1  g446(.A1(new_n629), .A2(KEYINPUT77), .B1(G110), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n629), .A2(KEYINPUT77), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n427), .B(new_n412), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n632), .A2(G110), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n431), .B(new_n636), .C1(new_n628), .C2(new_n627), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n622), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n622), .B1(new_n635), .B2(new_n637), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n193), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT25), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n613), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n613), .A2(G902), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n515), .A2(new_n519), .A3(new_n612), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT98), .B(G101), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G3));
  NAND2_X1  g466(.A1(new_n605), .A2(new_n193), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(G472), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n588), .A2(new_n654), .A3(new_n517), .A4(new_n649), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n498), .A2(new_n504), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n499), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n472), .B1(new_n487), .B2(new_n488), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n475), .B(KEYINPUT99), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(KEYINPUT33), .A3(new_n489), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT33), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n490), .B2(new_n495), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n499), .A2(G902), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n657), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n457), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n330), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n655), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT34), .B(G104), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n454), .B2(new_n456), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n413), .A2(new_n415), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n432), .A2(new_n421), .B1(new_n677), .B2(new_n402), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n450), .B1(new_n678), .B2(new_n393), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT20), .B1(new_n679), .B2(new_n455), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n452), .A2(new_n443), .A3(new_n453), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(KEYINPUT101), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n435), .A2(new_n436), .ZN(new_n683));
  INV_X1    g497(.A(G475), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n441), .B2(KEYINPUT89), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n676), .A2(new_n682), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n510), .A3(new_n508), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n330), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n655), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT102), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  OR2_X1    g506(.A1(new_n622), .A2(KEYINPUT36), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n635), .A2(new_n637), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n693), .B(new_n694), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n646), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n644), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n654), .A2(new_n588), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n515), .A2(new_n519), .A3(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT37), .B(G110), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT103), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(G12));
  OAI21_X1  g517(.A(new_n199), .B1(new_n328), .B2(new_n329), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n685), .A2(new_n683), .ZN(new_n706));
  INV_X1    g520(.A(G900), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n192), .B1(new_n195), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n682), .ZN(new_n710));
  AOI21_X1  g524(.A(KEYINPUT101), .B1(new_n680), .B2(new_n681), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n706), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n508), .A2(new_n510), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n517), .A2(new_n697), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n612), .A2(new_n705), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  NAND2_X1  g532(.A1(new_n312), .A2(new_n326), .ZN(new_n719));
  INV_X1    g533(.A(new_n327), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n312), .A2(new_n326), .A3(new_n327), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT38), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n508), .A2(new_n457), .A3(new_n510), .ZN(new_n725));
  INV_X1    g539(.A(new_n199), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n725), .A2(new_n726), .A3(new_n697), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n708), .B(KEYINPUT39), .Z(new_n729));
  NAND2_X1  g543(.A1(new_n517), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n728), .B1(KEYINPUT40), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n594), .A2(new_n561), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n193), .B1(new_n597), .B2(new_n551), .ZN(new_n733));
  OAI21_X1  g547(.A(G472), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n592), .A2(new_n611), .A3(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n731), .B(new_n735), .C1(KEYINPUT40), .C2(new_n730), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G143), .ZN(G45));
  INV_X1    g551(.A(G472), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n561), .B1(new_n585), .B2(new_n586), .ZN(new_n739));
  INV_X1    g553(.A(new_n595), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n599), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n738), .B1(new_n741), .B2(new_n601), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n608), .A3(new_n610), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n715), .B1(new_n743), .B2(new_n592), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n669), .A2(new_n457), .A3(new_n709), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(new_n705), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G146), .ZN(G48));
  NOR2_X1   g562(.A1(new_n389), .A2(new_n384), .ZN(new_n749));
  AOI211_X1 g563(.A(G469), .B(G902), .C1(new_n386), .C2(new_n388), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n516), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n612), .A2(new_n649), .A3(new_n671), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT41), .B(G113), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G15));
  NAND4_X1  g568(.A1(new_n612), .A2(new_n649), .A3(new_n688), .A4(new_n751), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n648), .B1(new_n743), .B2(new_n592), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n758), .A3(new_n688), .A4(new_n751), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  NOR2_X1   g575(.A1(new_n749), .A2(new_n750), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n512), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n704), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n197), .B1(new_n644), .B2(new_n696), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n612), .A2(new_n511), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n598), .A2(new_n551), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n520), .B1(new_n583), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(G902), .B1(new_n560), .B2(new_n576), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n770), .B(new_n649), .C1(new_n771), .C2(new_n738), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n198), .A2(new_n508), .A3(new_n457), .A4(new_n510), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n764), .A2(new_n768), .A3(new_n773), .A4(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n723), .A2(new_n774), .A3(new_n751), .A4(new_n199), .ZN(new_n776));
  OAI21_X1  g590(.A(KEYINPUT105), .B1(new_n776), .B2(new_n772), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  NAND3_X1  g593(.A1(new_n654), .A2(new_n697), .A3(new_n770), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n745), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n764), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G125), .ZN(G27));
  AND2_X1   g597(.A1(new_n579), .A2(new_n591), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n605), .A2(new_n607), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT75), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n605), .A2(new_n604), .A3(new_n607), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n603), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n649), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n357), .B1(new_n367), .B2(new_n371), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT84), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n387), .B1(new_n791), .B2(new_n372), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n384), .A3(new_n381), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n389), .A2(new_n384), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n385), .B(KEYINPUT106), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n512), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT107), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n721), .A2(new_n199), .A3(new_n722), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g615(.A(KEYINPUT107), .B(new_n512), .C1(new_n793), .C2(new_n796), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n789), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT42), .B1(new_n804), .B2(new_n746), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT42), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n745), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n785), .B1(new_n577), .B2(KEYINPUT32), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n807), .B(new_n649), .C1(new_n808), .C2(new_n742), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT108), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n803), .B2(new_n809), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n805), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(new_n347), .ZN(G33));
  XNOR2_X1  g631(.A(new_n714), .B(KEYINPUT109), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n811), .A2(new_n757), .A3(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G134), .ZN(G36));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n792), .B2(new_n381), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n378), .A2(KEYINPUT45), .A3(new_n382), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(G469), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n795), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(KEYINPUT46), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(KEYINPUT46), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n794), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n512), .ZN(new_n830));
  INV_X1    g644(.A(new_n729), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n821), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(KEYINPUT110), .A3(new_n512), .A4(new_n729), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n457), .A2(KEYINPUT111), .ZN(new_n834));
  INV_X1    g648(.A(new_n457), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n837), .A3(new_n669), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT43), .ZN(new_n839));
  INV_X1    g653(.A(new_n669), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n840), .A2(KEYINPUT43), .A3(new_n457), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n654), .A2(new_n588), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n843), .A3(new_n697), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT44), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n800), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n832), .A2(new_n833), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(G137), .ZN(G39));
  NOR4_X1   g663(.A1(new_n612), .A2(new_n649), .A3(new_n745), .A4(new_n800), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n829), .A2(KEYINPUT47), .A3(new_n512), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT47), .B1(new_n829), .B2(new_n512), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G140), .ZN(G42));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n192), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n855), .A2(new_n772), .ZN(new_n856));
  INV_X1    g670(.A(new_n724), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n763), .A2(new_n199), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT50), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n801), .A2(new_n751), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n780), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT119), .ZN(new_n864));
  INV_X1    g678(.A(new_n192), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n861), .A2(new_n648), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n735), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n835), .A3(new_n840), .A4(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n860), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n851), .A2(new_n852), .ZN(new_n870));
  INV_X1    g684(.A(new_n762), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n512), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n801), .A3(new_n856), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT51), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n649), .B1(new_n808), .B2(new_n742), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n862), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT48), .Z(new_n877));
  AOI21_X1  g691(.A(new_n191), .B1(new_n856), .B2(new_n764), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n866), .A2(new_n867), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n877), .B(new_n878), .C1(new_n670), .C2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n869), .A2(KEYINPUT51), .A3(new_n873), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n507), .A2(KEYINPUT113), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT113), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n505), .A2(new_n885), .A3(new_n506), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n835), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n670), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n655), .A2(new_n331), .A3(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n650), .A2(new_n890), .A3(new_n700), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n891), .B1(new_n805), .B2(new_n815), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n686), .A2(new_n709), .A3(new_n886), .A4(new_n884), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT114), .B1(new_n800), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n712), .A2(new_n887), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n328), .A2(new_n329), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n199), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n744), .A2(KEYINPUT115), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT115), .B1(new_n744), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n811), .A2(new_n781), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n819), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT116), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n744), .A2(new_n899), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n744), .A2(KEYINPUT115), .A3(new_n899), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n819), .A2(new_n903), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n892), .B1(new_n905), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n778), .A2(new_n752), .A3(new_n766), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT112), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n915), .A2(new_n760), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n915), .B2(new_n760), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n697), .A2(new_n708), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT118), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n797), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n704), .A2(new_n725), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n735), .A3(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n747), .A2(new_n924), .A3(new_n717), .A4(new_n782), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n925), .A2(KEYINPUT52), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(KEYINPUT52), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n914), .A2(new_n919), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT53), .ZN(new_n930));
  INV_X1    g744(.A(new_n747), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n717), .A2(new_n782), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(KEYINPUT117), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n932), .A2(KEYINPUT117), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n934), .A3(new_n924), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n927), .B1(new_n935), .B2(KEYINPUT52), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT53), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n936), .A2(new_n914), .A3(new_n919), .A4(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n930), .A2(KEYINPUT54), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n929), .A2(new_n937), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n915), .A2(new_n760), .A3(KEYINPUT53), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n936), .A2(new_n914), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n883), .A2(new_n945), .B1(G952), .B2(G953), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n871), .A2(KEYINPUT49), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n871), .A2(KEYINPUT49), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n649), .A2(new_n199), .A3(new_n512), .ZN(new_n949));
  NOR4_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n838), .A4(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n857), .A3(new_n867), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G75));
  AOI21_X1  g766(.A(new_n193), .B1(new_n940), .B2(new_n943), .ZN(new_n953));
  AOI21_X1  g767(.A(KEYINPUT56), .B1(new_n953), .B2(G210), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n302), .B1(new_n310), .B2(new_n311), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT120), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n235), .B(KEYINPUT55), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n954), .A2(new_n958), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n194), .A2(G952), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G51));
  XOR2_X1   g776(.A(new_n795), .B(KEYINPUT57), .Z(new_n963));
  AND3_X1   g777(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n941), .B1(new_n940), .B2(new_n943), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT121), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n386), .A2(new_n388), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT121), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n969), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n953), .A2(G469), .A3(new_n824), .A4(new_n823), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n961), .B1(new_n971), .B2(new_n972), .ZN(G54));
  AND2_X1   g787(.A1(KEYINPUT58), .A2(G475), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n953), .A2(new_n452), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n452), .B1(new_n953), .B2(new_n974), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n975), .A2(new_n976), .A3(new_n961), .ZN(G60));
  NOR2_X1   g791(.A1(new_n964), .A2(new_n965), .ZN(new_n978));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT59), .Z(new_n980));
  OR2_X1    g794(.A1(new_n666), .A2(new_n980), .ZN(new_n981));
  OAI22_X1  g795(.A1(new_n978), .A2(new_n981), .B1(G952), .B2(new_n194), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n939), .B2(new_n944), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT122), .ZN(new_n984));
  INV_X1    g798(.A(new_n666), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n983), .B2(new_n985), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n982), .B1(new_n986), .B2(new_n987), .ZN(G63));
  NAND2_X1  g802(.A1(new_n940), .A2(new_n943), .ZN(new_n989));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT60), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n645), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n961), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n991), .B1(new_n940), .B2(new_n943), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT123), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n996), .A2(new_n997), .A3(new_n695), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n996), .B2(new_n695), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n995), .B(KEYINPUT61), .C1(new_n998), .C2(new_n999), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(G66));
  OAI21_X1  g818(.A(G953), .B1(new_n196), .B2(new_n233), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT124), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n919), .A2(new_n891), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n1008), .B2(new_n614), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n956), .B1(G898), .B2(new_n194), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G69));
  NAND2_X1  g825(.A1(new_n534), .A2(new_n535), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n558), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n445), .A2(new_n446), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n614), .A2(G900), .ZN(new_n1016));
  INV_X1    g830(.A(new_n816), .ZN(new_n1017));
  AND4_X1   g831(.A1(new_n1017), .A2(new_n819), .A3(new_n934), .A4(new_n933), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n875), .A2(new_n704), .A3(new_n725), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n832), .A2(new_n833), .A3(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1018), .A2(new_n848), .A3(new_n853), .A4(new_n1020), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1015), .B(new_n1016), .C1(new_n1021), .C2(new_n614), .ZN(new_n1022));
  INV_X1    g836(.A(new_n730), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n757), .A2(new_n1023), .A3(new_n801), .A4(new_n889), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n848), .A2(new_n853), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n736), .A2(new_n933), .A3(new_n934), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1026), .A2(KEYINPUT62), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT125), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1025), .A2(new_n1028), .A3(KEYINPUT125), .A4(new_n1027), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n614), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1022), .B1(new_n1033), .B2(new_n1015), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1034), .B(new_n1035), .ZN(G72));
  NAND3_X1  g850(.A1(new_n1031), .A2(new_n1008), .A3(new_n1032), .ZN(new_n1037));
  NAND2_X1  g851(.A1(G472), .A2(G902), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT63), .Z(new_n1039));
  NAND2_X1  g853(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n732), .ZN(new_n1041));
  INV_X1    g855(.A(KEYINPUT127), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1039), .B1(new_n1021), .B2(new_n1007), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n740), .ZN(new_n1044));
  AND2_X1   g858(.A1(new_n930), .A2(new_n938), .ZN(new_n1045));
  INV_X1    g859(.A(new_n732), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1046), .A2(new_n595), .A3(new_n1039), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT126), .Z(new_n1048));
  AOI21_X1  g862(.A(new_n961), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g863(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(new_n1044), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1046), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1052));
  OAI21_X1  g866(.A(KEYINPUT127), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1050), .A2(new_n1053), .ZN(G57));
endmodule


