//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI21_X1  g031(.A(KEYINPUT66), .B1(new_n452), .B2(G2106), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n454), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n452), .A2(KEYINPUT66), .A3(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G101), .A3(G2104), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT69), .Z(new_n476));
  OAI21_X1  g051(.A(KEYINPUT68), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n464), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n463), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT67), .B(G2105), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n478), .A2(G137), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n473), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  AND2_X1   g058(.A1(new_n478), .A2(new_n479), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n474), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n480), .C2(G112), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n478), .A2(new_n479), .A3(new_n472), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT70), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n465), .B2(G2104), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n465), .A2(G2104), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n479), .B(new_n495), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n474), .B2(G114), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(G2104), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT4), .A2(G138), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n478), .A2(new_n479), .A3(new_n480), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  OAI21_X1  g084(.A(G138), .B1(new_n470), .B2(new_n471), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(new_n467), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT72), .B1(new_n499), .B2(new_n505), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n506), .A2(new_n512), .A3(new_n513), .ZN(G164));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n517), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT73), .A3(G50), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n523), .B2(KEYINPUT5), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT74), .A3(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n516), .ZN(new_n530));
  INV_X1    g105(.A(G88), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n519), .B(new_n521), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n529), .A2(G62), .ZN(new_n534));
  NAND2_X1  g109(.A1(G75), .A2(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G166));
  AND2_X1   g112(.A1(new_n529), .A2(new_n516), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G89), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n529), .A2(G63), .A3(G651), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n520), .A2(G51), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  AOI22_X1  g120(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n533), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n520), .A2(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n530), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n529), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n533), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n520), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n530), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  AOI22_X1  g138(.A1(new_n529), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n533), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n538), .A2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n520), .A2(G53), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND3_X1  g147(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT75), .Z(new_n574));
  NAND3_X1  g149(.A1(new_n529), .A2(G87), .A3(new_n516), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND4_X1  g152(.A1(new_n527), .A2(G86), .A3(new_n528), .A4(new_n516), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n517), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n527), .A2(G61), .A3(new_n528), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(KEYINPUT76), .B1(G73), .B2(G543), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n529), .A2(new_n583), .A3(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n580), .B1(new_n585), .B2(G651), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n520), .A2(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI221_X1 g165(.A(new_n588), .B1(new_n530), .B2(new_n589), .C1(new_n590), .C2(new_n533), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n538), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n529), .A2(G66), .ZN(new_n596));
  INV_X1    g171(.A(G79), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n523), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G284));
  XNOR2_X1  g177(.A(G284), .B(KEYINPUT77), .ZN(G321));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT78), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n610), .ZN(G297));
  XNOR2_X1  g186(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n601), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n601), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n490), .A2(G123), .ZN(new_n619));
  OAI221_X1 g194(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n480), .C2(G111), .ZN(new_n620));
  INV_X1    g195(.A(G135), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n619), .B(new_n620), .C1(new_n485), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT82), .B(G2096), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NOR2_X1   g199(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  AND2_X1   g203(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n624), .B(new_n630), .C1(new_n629), .C2(new_n628), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  INV_X1    g207(.A(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  OAI21_X1  g210(.A(KEYINPUT14), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT84), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n639), .B(new_n642), .Z(new_n643));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n643), .A2(new_n645), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n643), .A2(new_n645), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(G14), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT85), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2067), .B(G2678), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(new_n660), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n661), .B1(new_n657), .B2(new_n665), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n663), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2096), .B(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n672), .A2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n679), .ZN(new_n682));
  INV_X1    g257(.A(G1991), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(G1996), .ZN(new_n688));
  INV_X1    g263(.A(G1986), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT86), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1981), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n687), .A2(new_n690), .A3(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(G229));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(G4), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n600), .B2(G16), .ZN(new_n701));
  INV_X1    g276(.A(G1348), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n557), .A2(new_n699), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n699), .A2(G19), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT90), .B(G1341), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OR3_X1    g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT28), .ZN(new_n709));
  INV_X1    g284(.A(G26), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G29), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n490), .A2(G128), .ZN(new_n713));
  OAI221_X1 g288(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n480), .C2(G116), .ZN(new_n714));
  INV_X1    g289(.A(G140), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n713), .B(new_n714), .C1(new_n485), .C2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n712), .B1(new_n716), .B2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n717), .B2(new_n709), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G2067), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n707), .B1(new_n704), .B2(new_n705), .ZN(new_n720));
  NOR2_X1   g295(.A1(G5), .A2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G171), .B2(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G1961), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n708), .A2(new_n719), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n718), .A2(G2067), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n703), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n699), .A2(G20), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G299), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1956), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n699), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G168), .B2(new_n699), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT99), .B(G1966), .Z(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G28), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT30), .ZN(new_n738));
  AOI21_X1  g313(.A(G29), .B1(new_n737), .B2(KEYINPUT30), .ZN(new_n739));
  OR2_X1    g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT31), .A2(G11), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n738), .A2(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n622), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n734), .B2(new_n735), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n743), .ZN(new_n747));
  INV_X1    g322(.A(G2078), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AND4_X1   g324(.A1(new_n732), .A2(new_n736), .A3(new_n745), .A4(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n751), .A2(G2072), .B1(new_n743), .B2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT91), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n755));
  INV_X1    g330(.A(G139), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n754), .A2(new_n755), .B1(new_n756), .B2(new_n485), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n755), .B2(new_n754), .ZN(new_n758));
  NAND2_X1  g333(.A1(G115), .A2(G2104), .ZN(new_n759));
  INV_X1    g334(.A(G127), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n467), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n480), .B1(new_n761), .B2(KEYINPUT92), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT92), .B2(new_n761), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n752), .B1(new_n765), .B2(new_n743), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n751), .A2(G2072), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n743), .A2(G35), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT101), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n493), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n490), .A2(G129), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT26), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n463), .A2(G2105), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n778), .A2(new_n779), .B1(G105), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G141), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n775), .B(new_n781), .C1(new_n485), .C2(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G32), .B(new_n783), .S(G29), .Z(new_n784));
  AND2_X1   g359(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(KEYINPUT97), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT98), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n769), .A2(new_n774), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n727), .A2(new_n750), .A3(new_n768), .A4(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n788), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n785), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT24), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G34), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G34), .ZN(new_n797));
  AOI21_X1  g372(.A(G29), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n482), .B2(G29), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT95), .Z(new_n800));
  OAI22_X1  g375(.A1(new_n800), .A2(G2084), .B1(new_n722), .B2(G1961), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n794), .A2(new_n801), .A3(KEYINPUT100), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT100), .B1(new_n794), .B2(new_n801), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n800), .A2(G2084), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT98), .B1(new_n787), .B2(new_n788), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n774), .A2(new_n769), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n804), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n792), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G22), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G166), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT89), .B(G1971), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n699), .A2(G6), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n586), .B2(new_n699), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT32), .B(G1981), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(G16), .A2(G23), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G288), .B2(new_n699), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT33), .B(G1976), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n817), .A2(new_n818), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n815), .A2(new_n819), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT34), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n743), .A2(G25), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT87), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n486), .A2(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n490), .A2(G119), .ZN(new_n831));
  OAI221_X1 g406(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n480), .C2(G107), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n829), .B1(new_n834), .B2(new_n743), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT35), .B(G1991), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT88), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n835), .B(new_n837), .Z(new_n838));
  MUX2_X1   g413(.A(G24), .B(G290), .S(G16), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G1986), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n811), .B1(new_n827), .B2(new_n841), .ZN(new_n842));
  NOR4_X1   g417(.A1(new_n826), .A2(KEYINPUT36), .A3(new_n838), .A4(new_n840), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n810), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(G311));
  NAND2_X1  g420(.A1(new_n844), .A2(KEYINPUT104), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n810), .B(new_n847), .C1(new_n842), .C2(new_n843), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G150));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n601), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n520), .A2(G55), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n530), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n529), .A2(G67), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n533), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n557), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n553), .A2(new_n556), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n852), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n850), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n865), .B2(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n865), .A2(new_n850), .A3(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n860), .A2(KEYINPUT37), .A3(G860), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT37), .B1(new_n860), .B2(G860), .ZN(new_n872));
  OAI22_X1  g447(.A1(new_n868), .A2(new_n869), .B1(new_n871), .B2(new_n872), .ZN(G145));
  XOR2_X1   g448(.A(new_n493), .B(new_n622), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n490), .A2(G130), .ZN(new_n875));
  OAI221_X1 g450(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n480), .C2(G118), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n875), .B(new_n876), .C1(new_n485), .C2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n482), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n874), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n833), .B(new_n783), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n508), .A2(new_n511), .A3(new_n499), .A4(new_n505), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n881), .B(new_n883), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n765), .A2(KEYINPUT106), .A3(KEYINPUT107), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT106), .B1(new_n765), .B2(KEYINPUT107), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n884), .B1(new_n886), .B2(new_n885), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n880), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n879), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n874), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n885), .A2(new_n886), .ZN(new_n893));
  INV_X1    g468(.A(new_n884), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n895), .A3(new_n887), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n716), .B(new_n627), .Z(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n890), .A2(new_n898), .A3(new_n896), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(G395));
  INV_X1    g483(.A(new_n864), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n615), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n600), .A2(new_n604), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n595), .A2(G299), .A3(new_n599), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n914), .B1(new_n918), .B2(new_n910), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(G288), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n921), .A2(G166), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(G166), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n922), .A2(new_n923), .A3(G305), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(G305), .B1(new_n922), .B2(new_n923), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(KEYINPUT42), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n928), .B1(new_n929), .B2(new_n924), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n919), .A2(new_n920), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n930), .A2(new_n927), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n931), .B1(new_n932), .B2(new_n919), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n920), .B1(new_n932), .B2(new_n919), .ZN(new_n934));
  OAI21_X1  g509(.A(G868), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n860), .A2(new_n606), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(G295));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(G331));
  INV_X1    g513(.A(new_n917), .ZN(new_n939));
  XNOR2_X1  g514(.A(G171), .B(G286), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n940), .A2(new_n864), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n864), .ZN(new_n942));
  AOI22_X1  g517(.A1(new_n939), .A2(new_n915), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n913), .A3(new_n942), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n943), .A2(new_n945), .B1(new_n929), .B2(new_n924), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n941), .A2(new_n942), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n916), .B2(new_n917), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(new_n925), .A3(new_n926), .A4(new_n944), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n946), .A2(new_n949), .A3(new_n950), .A4(new_n902), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT110), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT44), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n946), .A2(new_n949), .A3(new_n902), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n951), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n952), .A2(new_n955), .A3(KEYINPUT44), .A4(new_n951), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(G397));
  NOR2_X1   g534(.A1(G290), .A2(G1986), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT112), .Z(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n882), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(KEYINPUT111), .B(G40), .Z(new_n966));
  NAND4_X1  g541(.A1(new_n473), .A2(new_n476), .A3(new_n481), .A4(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(G1986), .A3(G290), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT113), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n716), .B(G2067), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n783), .B(G1996), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n968), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n975), .B(KEYINPUT114), .Z(new_n976));
  INV_X1    g551(.A(new_n968), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n834), .A2(new_n837), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n834), .A2(new_n837), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n972), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1971), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n499), .A2(new_n505), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT72), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n505), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n508), .A4(new_n511), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n988), .B2(new_n962), .ZN(new_n989));
  INV_X1    g564(.A(new_n967), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n882), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n983), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n512), .A2(new_n513), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n997), .B2(new_n987), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n988), .A2(new_n962), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n882), .A2(new_n962), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n967), .B1(new_n1003), .B2(new_n999), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1000), .A2(new_n1002), .A3(new_n769), .A4(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT115), .B(new_n983), .C1(new_n989), .C2(new_n992), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n995), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(G166), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT55), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1009), .B(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(KEYINPUT119), .B(new_n990), .C1(new_n1003), .C2(new_n999), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n999), .B1(new_n882), .B2(new_n962), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n967), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n988), .A2(new_n999), .A3(new_n962), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1014), .A2(new_n769), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1019), .A2(new_n993), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1013), .B1(new_n1020), .B2(new_n1008), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1008), .B1(new_n1003), .B2(new_n990), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n585), .A2(G651), .ZN(new_n1025));
  INV_X1    g600(.A(new_n580), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g602(.A(KEYINPUT49), .B(new_n580), .C1(new_n585), .C2(G651), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1023), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1032), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AND3_X1   g612(.A1(G288), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1003), .A2(new_n990), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(G8), .C1(new_n1037), .C2(G288), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1036), .A2(KEYINPUT117), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1022), .B(new_n1041), .C1(new_n1037), .C2(G288), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1033), .A2(new_n1035), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1011), .A2(new_n1021), .A3(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT125), .ZN(new_n1047));
  INV_X1    g622(.A(new_n735), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n998), .A2(KEYINPUT45), .B1(new_n965), .B2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n988), .A2(new_n1049), .A3(KEYINPUT45), .A4(new_n962), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n990), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1048), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G2084), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1000), .A2(new_n1002), .A3(new_n1054), .A4(new_n1004), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G8), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G286), .A2(G8), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT51), .A3(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1056), .A2(G8), .A3(G286), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(G8), .C1(new_n1056), .C2(G286), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  OR3_X1    g638(.A1(new_n547), .A2(new_n550), .A3(KEYINPUT54), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT54), .B1(new_n547), .B2(new_n550), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT124), .B(G2078), .ZN(new_n1067));
  AND2_X1   g642(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1068));
  AND4_X1   g643(.A1(G160), .A2(new_n991), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n965), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n989), .A2(new_n992), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n748), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1075));
  INV_X1    g650(.A(G1961), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1070), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g653(.A1(new_n1073), .A2(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1051), .A2(new_n990), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT45), .B1(new_n882), .B2(new_n962), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1001), .A2(new_n964), .B1(KEYINPUT120), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1080), .A2(KEYINPUT123), .A3(new_n748), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT53), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT123), .B1(new_n1085), .B2(new_n748), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1079), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1078), .B1(new_n1087), .B2(new_n1066), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1063), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1014), .A2(new_n1018), .A3(new_n1017), .ZN(new_n1090));
  INV_X1    g665(.A(G1956), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1091), .B1(new_n1071), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g669(.A1(G299), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n566), .A2(KEYINPUT57), .A3(new_n569), .A4(new_n567), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n990), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n996), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n1103), .B2(new_n1002), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1039), .A2(G2067), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n601), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1093), .A2(new_n1099), .A3(new_n1097), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1098), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n999), .B1(new_n988), .B2(new_n962), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1004), .B1(new_n1112), .B2(KEYINPUT116), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1102), .A2(new_n996), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n702), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1105), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1111), .A2(new_n601), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1093), .A2(new_n1119), .A3(new_n1097), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1071), .A2(new_n1092), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1097), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1098), .B1(new_n1123), .B2(KEYINPUT61), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1118), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  AOI22_X1  g701(.A1(new_n1071), .A2(new_n685), .B1(new_n1039), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n1128));
  OR3_X1    g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n862), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n600), .A4(new_n1116), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1127), .B2(new_n862), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1109), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1089), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1063), .A2(KEYINPUT62), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1087), .A2(G171), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1059), .A2(new_n1137), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1047), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1008), .B(G286), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1011), .A2(new_n1141), .A3(new_n1021), .A4(new_n1045), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(KEYINPUT121), .A3(new_n1143), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1057), .A2(new_n1143), .A3(G286), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1007), .A2(G8), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1013), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1148), .A2(new_n1011), .A3(new_n1045), .A4(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1146), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1153));
  INV_X1    g728(.A(G288), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1037), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n586), .A2(new_n1030), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1023), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1011), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n1045), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1152), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n982), .B1(new_n1140), .B2(new_n1160), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n969), .B(KEYINPUT48), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  OAI22_X1  g740(.A1(new_n976), .A2(new_n979), .B1(G2067), .B2(new_n716), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n968), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT46), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n977), .B2(G1996), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n968), .B1(new_n973), .B2(new_n783), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n968), .A2(KEYINPUT46), .A3(new_n685), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT47), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1165), .A2(new_n1167), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1161), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g750(.A1(G227), .A2(new_n460), .ZN(new_n1177));
  AND4_X1   g751(.A1(new_n653), .A2(new_n696), .A3(new_n697), .A4(new_n1177), .ZN(new_n1178));
  AND3_X1   g752(.A1(new_n1178), .A2(new_n903), .A3(new_n956), .ZN(G308));
  NAND3_X1  g753(.A1(new_n1178), .A2(new_n903), .A3(new_n956), .ZN(G225));
endmodule


