

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(n971), .ZN(n751) );
  AND2_X1 U556 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U557 ( .A1(n689), .A2(n776), .ZN(n714) );
  NOR2_X1 U558 ( .A1(G651), .A2(n649), .ZN(n648) );
  AND2_X1 U559 ( .A1(n529), .A2(n528), .ZN(G160) );
  INV_X1 U560 ( .A(G2105), .ZN(n524) );
  NOR2_X1 U561 ( .A1(G2104), .A2(n524), .ZN(n863) );
  NAND2_X1 U562 ( .A1(G125), .A2(n863), .ZN(n521) );
  AND2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n864) );
  NAND2_X1 U564 ( .A1(G113), .A2(n864), .ZN(n520) );
  AND2_X1 U565 ( .A1(n521), .A2(n520), .ZN(n529) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U567 ( .A(KEYINPUT17), .B(n522), .Z(n868) );
  NAND2_X1 U568 ( .A1(G137), .A2(n868), .ZN(n523) );
  XNOR2_X1 U569 ( .A(n523), .B(KEYINPUT64), .ZN(n527) );
  AND2_X1 U570 ( .A1(n524), .A2(G2104), .ZN(n867) );
  NAND2_X1 U571 ( .A1(G101), .A2(n867), .ZN(n525) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n525), .Z(n526) );
  AND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n637) );
  NAND2_X1 U575 ( .A1(G85), .A2(n637), .ZN(n531) );
  XOR2_X1 U576 ( .A(G543), .B(KEYINPUT0), .Z(n649) );
  INV_X1 U577 ( .A(G651), .ZN(n532) );
  NOR2_X1 U578 ( .A1(n649), .A2(n532), .ZN(n640) );
  NAND2_X1 U579 ( .A1(G72), .A2(n640), .ZN(n530) );
  NAND2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n537) );
  NOR2_X1 U581 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n533), .Z(n653) );
  NAND2_X1 U583 ( .A1(G60), .A2(n653), .ZN(n535) );
  NAND2_X1 U584 ( .A1(G47), .A2(n648), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n536) );
  OR2_X1 U586 ( .A1(n537), .A2(n536), .ZN(G290) );
  XOR2_X1 U587 ( .A(G2438), .B(G2454), .Z(n539) );
  XNOR2_X1 U588 ( .A(G2435), .B(G2430), .ZN(n538) );
  XNOR2_X1 U589 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U590 ( .A(n540), .B(G2427), .Z(n542) );
  XNOR2_X1 U591 ( .A(G1341), .B(G1348), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n542), .B(n541), .ZN(n546) );
  XOR2_X1 U593 ( .A(G2443), .B(G2446), .Z(n544) );
  XNOR2_X1 U594 ( .A(KEYINPUT100), .B(G2451), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U596 ( .A(n546), .B(n545), .Z(n547) );
  AND2_X1 U597 ( .A1(G14), .A2(n547), .ZN(G401) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  NAND2_X1 U602 ( .A1(G88), .A2(n637), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G75), .A2(n640), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U605 ( .A1(n648), .A2(G50), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT80), .ZN(n552) );
  NAND2_X1 U607 ( .A1(G62), .A2(n653), .ZN(n551) );
  NAND2_X1 U608 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U609 ( .A(KEYINPUT81), .B(n553), .Z(n554) );
  NOR2_X1 U610 ( .A1(n555), .A2(n554), .ZN(G166) );
  NAND2_X1 U611 ( .A1(n637), .A2(G89), .ZN(n556) );
  XNOR2_X1 U612 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G76), .A2(n640), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U615 ( .A(n559), .B(KEYINPUT5), .ZN(n566) );
  XNOR2_X1 U616 ( .A(KEYINPUT6), .B(KEYINPUT71), .ZN(n564) );
  NAND2_X1 U617 ( .A1(n648), .A2(G51), .ZN(n560) );
  XNOR2_X1 U618 ( .A(n560), .B(KEYINPUT70), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G63), .A2(n653), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U621 ( .A(n564), .B(n563), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U623 ( .A(KEYINPUT7), .B(n567), .ZN(G168) );
  XOR2_X1 U624 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U626 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n828) );
  NAND2_X1 U628 ( .A1(n828), .A2(G567), .ZN(n569) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  INV_X1 U630 ( .A(G860), .ZN(n608) );
  NAND2_X1 U631 ( .A1(G43), .A2(n648), .ZN(n579) );
  NAND2_X1 U632 ( .A1(n653), .A2(G56), .ZN(n570) );
  XNOR2_X1 U633 ( .A(KEYINPUT14), .B(n570), .ZN(n576) );
  NAND2_X1 U634 ( .A1(n637), .A2(G81), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G68), .A2(n640), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT13), .B(n574), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT67), .B(n577), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U642 ( .A(n580), .B(KEYINPUT68), .ZN(n969) );
  OR2_X1 U643 ( .A1(n608), .A2(n969), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G64), .A2(n653), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G52), .A2(n648), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n640), .A2(G77), .ZN(n583) );
  XOR2_X1 U648 ( .A(KEYINPUT65), .B(n583), .Z(n585) );
  NAND2_X1 U649 ( .A1(n637), .A2(G90), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT9), .B(n586), .Z(n587) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(KEYINPUT66), .B(n589), .ZN(G171) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G301), .A2(G868), .ZN(n599) );
  NAND2_X1 U656 ( .A1(G66), .A2(n653), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G92), .A2(n637), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G79), .A2(n640), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G54), .A2(n648), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n595), .A2(n594), .ZN(n597) );
  XNOR2_X1 U663 ( .A(KEYINPUT69), .B(KEYINPUT15), .ZN(n596) );
  XNOR2_X1 U664 ( .A(n597), .B(n596), .ZN(n881) );
  INV_X1 U665 ( .A(n881), .ZN(n973) );
  INV_X1 U666 ( .A(G868), .ZN(n611) );
  NAND2_X1 U667 ( .A1(n973), .A2(n611), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U669 ( .A1(G65), .A2(n653), .ZN(n601) );
  NAND2_X1 U670 ( .A1(G53), .A2(n648), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G91), .A2(n637), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G78), .A2(n640), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n970) );
  INV_X1 U676 ( .A(n970), .ZN(G299) );
  NOR2_X1 U677 ( .A1(G286), .A2(n611), .ZN(n607) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n606) );
  NOR2_X1 U679 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n608), .A2(G559), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n609), .A2(n881), .ZN(n610) );
  XNOR2_X1 U682 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(n973), .A2(n611), .ZN(n612) );
  XOR2_X1 U684 ( .A(KEYINPUT72), .B(n612), .Z(n613) );
  NOR2_X1 U685 ( .A1(G559), .A2(n613), .ZN(n615) );
  NOR2_X1 U686 ( .A1(n969), .A2(G868), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U688 ( .A1(G123), .A2(n863), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(KEYINPUT18), .ZN(n624) );
  NAND2_X1 U690 ( .A1(G111), .A2(n864), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G99), .A2(n867), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U693 ( .A(KEYINPUT74), .B(n619), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G135), .A2(n868), .ZN(n620) );
  XNOR2_X1 U695 ( .A(KEYINPUT73), .B(n620), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n929) );
  XOR2_X1 U698 ( .A(n929), .B(G2096), .Z(n626) );
  XNOR2_X1 U699 ( .A(G2100), .B(KEYINPUT75), .ZN(n625) );
  NAND2_X1 U700 ( .A1(n626), .A2(n625), .ZN(G156) );
  NAND2_X1 U701 ( .A1(G67), .A2(n653), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G55), .A2(n648), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n633) );
  NAND2_X1 U704 ( .A1(G93), .A2(n637), .ZN(n630) );
  NAND2_X1 U705 ( .A1(G80), .A2(n640), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U707 ( .A(KEYINPUT77), .B(n631), .Z(n632) );
  NOR2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n664) );
  NAND2_X1 U709 ( .A1(G559), .A2(n881), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n634), .B(n969), .ZN(n662) );
  XNOR2_X1 U711 ( .A(KEYINPUT76), .B(n662), .ZN(n635) );
  NOR2_X1 U712 ( .A1(G860), .A2(n635), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n664), .B(n636), .ZN(G145) );
  NAND2_X1 U714 ( .A1(G61), .A2(n653), .ZN(n639) );
  NAND2_X1 U715 ( .A1(G86), .A2(n637), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n644) );
  NAND2_X1 U717 ( .A1(G73), .A2(n640), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n641), .B(KEYINPUT2), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n642), .B(KEYINPUT79), .ZN(n643) );
  NOR2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n648), .A2(G48), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n647), .B(KEYINPUT78), .ZN(n655) );
  NAND2_X1 U725 ( .A1(G49), .A2(n648), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G87), .A2(n649), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(G288) );
  XNOR2_X1 U730 ( .A(G166), .B(n664), .ZN(n661) );
  XNOR2_X1 U731 ( .A(KEYINPUT82), .B(G305), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n656), .B(G288), .ZN(n657) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(n657), .ZN(n659) );
  XNOR2_X1 U734 ( .A(G290), .B(n970), .ZN(n658) );
  XNOR2_X1 U735 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n880) );
  XNOR2_X1 U737 ( .A(n880), .B(n662), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n663), .A2(G868), .ZN(n666) );
  OR2_X1 U739 ( .A1(G868), .A2(n664), .ZN(n665) );
  NAND2_X1 U740 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U745 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XOR2_X1 U746 ( .A(KEYINPUT83), .B(G44), .Z(n671) );
  XNOR2_X1 U747 ( .A(KEYINPUT3), .B(n671), .ZN(G218) );
  NAND2_X1 U748 ( .A1(G120), .A2(G69), .ZN(n672) );
  NOR2_X1 U749 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(G108), .A2(n673), .ZN(n834) );
  NAND2_X1 U751 ( .A1(n834), .A2(G567), .ZN(n679) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U754 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G96), .A2(n676), .ZN(n833) );
  NAND2_X1 U756 ( .A1(G2106), .A2(n833), .ZN(n677) );
  XNOR2_X1 U757 ( .A(KEYINPUT84), .B(n677), .ZN(n678) );
  NAND2_X1 U758 ( .A1(n679), .A2(n678), .ZN(n913) );
  NAND2_X1 U759 ( .A1(G483), .A2(G661), .ZN(n680) );
  NOR2_X1 U760 ( .A1(n913), .A2(n680), .ZN(n830) );
  NAND2_X1 U761 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U762 ( .A1(n867), .A2(G102), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G114), .A2(n864), .ZN(n681) );
  XOR2_X1 U764 ( .A(KEYINPUT85), .B(n681), .Z(n682) );
  NAND2_X1 U765 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U766 ( .A1(G126), .A2(n863), .ZN(n685) );
  NAND2_X1 U767 ( .A1(G138), .A2(n868), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U769 ( .A1(n687), .A2(n686), .ZN(G164) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NAND2_X1 U771 ( .A1(G40), .A2(G160), .ZN(n688) );
  XNOR2_X1 U772 ( .A(n688), .B(KEYINPUT86), .ZN(n777) );
  INV_X1 U773 ( .A(n777), .ZN(n689) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n776) );
  NAND2_X1 U775 ( .A1(G8), .A2(n714), .ZN(n771) );
  NOR2_X1 U776 ( .A1(G1966), .A2(n771), .ZN(n748) );
  NOR2_X1 U777 ( .A1(G2084), .A2(n714), .ZN(n744) );
  NOR2_X1 U778 ( .A1(n748), .A2(n744), .ZN(n690) );
  NAND2_X1 U779 ( .A1(G8), .A2(n690), .ZN(n691) );
  XNOR2_X1 U780 ( .A(n691), .B(KEYINPUT30), .ZN(n692) );
  NOR2_X1 U781 ( .A1(G168), .A2(n692), .ZN(n696) );
  INV_X1 U782 ( .A(G1961), .ZN(n1004) );
  NAND2_X1 U783 ( .A1(n714), .A2(n1004), .ZN(n694) );
  INV_X1 U784 ( .A(n714), .ZN(n717) );
  XNOR2_X1 U785 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NAND2_X1 U786 ( .A1(n717), .A2(n943), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n704) );
  NOR2_X1 U788 ( .A1(n704), .A2(G171), .ZN(n695) );
  NOR2_X1 U789 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U790 ( .A(KEYINPUT31), .B(n697), .Z(n742) );
  INV_X1 U791 ( .A(G8), .ZN(n703) );
  NOR2_X1 U792 ( .A1(G2090), .A2(n714), .ZN(n698) );
  XNOR2_X1 U793 ( .A(KEYINPUT95), .B(n698), .ZN(n701) );
  NOR2_X1 U794 ( .A1(G1971), .A2(n771), .ZN(n699) );
  NOR2_X1 U795 ( .A1(G166), .A2(n699), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n702) );
  OR2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n737) );
  AND2_X1 U798 ( .A1(n742), .A2(n737), .ZN(n736) );
  AND2_X1 U799 ( .A1(G171), .A2(n704), .ZN(n705) );
  XNOR2_X1 U800 ( .A(n705), .B(KEYINPUT93), .ZN(n735) );
  NAND2_X1 U801 ( .A1(n717), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U802 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  AND2_X1 U803 ( .A1(G1956), .A2(n714), .ZN(n707) );
  NOR2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n710) );
  NOR2_X1 U805 ( .A1(n710), .A2(n970), .ZN(n709) );
  XOR2_X1 U806 ( .A(n709), .B(KEYINPUT28), .Z(n732) );
  NAND2_X1 U807 ( .A1(n970), .A2(n710), .ZN(n730) );
  NAND2_X1 U808 ( .A1(G1348), .A2(n714), .ZN(n712) );
  NAND2_X1 U809 ( .A1(G2067), .A2(n717), .ZN(n711) );
  NAND2_X1 U810 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U811 ( .A1(n713), .A2(n973), .ZN(n728) );
  OR2_X1 U812 ( .A1(n713), .A2(n973), .ZN(n726) );
  AND2_X1 U813 ( .A1(n714), .A2(G1341), .ZN(n719) );
  AND2_X1 U814 ( .A1(KEYINPUT26), .A2(n719), .ZN(n715) );
  NOR2_X1 U815 ( .A1(KEYINPUT94), .A2(n715), .ZN(n716) );
  NOR2_X1 U816 ( .A1(n969), .A2(n716), .ZN(n724) );
  NAND2_X1 U817 ( .A1(G1996), .A2(n717), .ZN(n718) );
  XNOR2_X1 U818 ( .A(KEYINPUT26), .B(n718), .ZN(n721) );
  INV_X1 U819 ( .A(n719), .ZN(n720) );
  NAND2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U821 ( .A1(KEYINPUT94), .A2(n722), .ZN(n723) );
  NAND2_X1 U822 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U823 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U825 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U827 ( .A(n733), .B(KEYINPUT29), .Z(n734) );
  NAND2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n743) );
  NAND2_X1 U829 ( .A1(n736), .A2(n743), .ZN(n740) );
  INV_X1 U830 ( .A(n737), .ZN(n738) );
  OR2_X1 U831 ( .A1(n738), .A2(G286), .ZN(n739) );
  NAND2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U833 ( .A(n741), .B(KEYINPUT32), .ZN(n766) );
  NAND2_X1 U834 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U835 ( .A1(G8), .A2(n744), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  OR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n765) );
  NAND2_X1 U838 ( .A1(n766), .A2(n765), .ZN(n750) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n756), .A2(n749), .ZN(n986) );
  NAND2_X1 U842 ( .A1(n750), .A2(n986), .ZN(n753) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NOR2_X1 U844 ( .A1(n771), .A2(n751), .ZN(n752) );
  NOR2_X1 U845 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  XNOR2_X1 U846 ( .A(n755), .B(KEYINPUT96), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  OR2_X1 U848 ( .A1(n771), .A2(n757), .ZN(n758) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n966) );
  NAND2_X1 U850 ( .A1(n758), .A2(n966), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n764) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n761) );
  XOR2_X1 U853 ( .A(n761), .B(KEYINPUT24), .Z(n762) );
  NOR2_X1 U854 ( .A1(n771), .A2(n762), .ZN(n763) );
  NOR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n775) );
  AND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n769) );
  NAND2_X1 U857 ( .A1(G166), .A2(G8), .ZN(n767) );
  NOR2_X1 U858 ( .A1(G2090), .A2(n767), .ZN(n768) );
  NOR2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n770), .B(KEYINPUT97), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U862 ( .A(n773), .B(KEYINPUT98), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n811) );
  XNOR2_X1 U864 ( .A(G1986), .B(G290), .ZN(n979) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n823) );
  AND2_X1 U866 ( .A1(n979), .A2(n823), .ZN(n809) );
  NAND2_X1 U867 ( .A1(n867), .A2(G104), .ZN(n778) );
  XOR2_X1 U868 ( .A(KEYINPUT87), .B(n778), .Z(n780) );
  NAND2_X1 U869 ( .A1(n868), .A2(G140), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n781), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G128), .A2(n863), .ZN(n783) );
  NAND2_X1 U873 ( .A1(G116), .A2(n864), .ZN(n782) );
  NAND2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U875 ( .A(KEYINPUT88), .B(n784), .Z(n785) );
  XNOR2_X1 U876 ( .A(KEYINPUT35), .B(n785), .ZN(n786) );
  NOR2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U878 ( .A(KEYINPUT36), .B(n788), .Z(n860) );
  XOR2_X1 U879 ( .A(KEYINPUT37), .B(G2067), .Z(n820) );
  NAND2_X1 U880 ( .A1(n860), .A2(n820), .ZN(n789) );
  XNOR2_X1 U881 ( .A(KEYINPUT89), .B(n789), .ZN(n936) );
  NAND2_X1 U882 ( .A1(n823), .A2(n936), .ZN(n818) );
  NAND2_X1 U883 ( .A1(G119), .A2(n863), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G107), .A2(n864), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G95), .A2(n867), .ZN(n793) );
  NAND2_X1 U887 ( .A1(G131), .A2(n868), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U890 ( .A(KEYINPUT90), .B(n796), .ZN(n859) );
  XNOR2_X1 U891 ( .A(KEYINPUT91), .B(G1991), .ZN(n941) );
  NOR2_X1 U892 ( .A1(n859), .A2(n941), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G141), .A2(n868), .ZN(n797) );
  XNOR2_X1 U894 ( .A(n797), .B(KEYINPUT92), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G129), .A2(n863), .ZN(n799) );
  NAND2_X1 U896 ( .A1(G117), .A2(n864), .ZN(n798) );
  NAND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n867), .A2(G105), .ZN(n800) );
  XOR2_X1 U899 ( .A(KEYINPUT38), .B(n800), .Z(n801) );
  NOR2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n874) );
  AND2_X1 U902 ( .A1(n874), .A2(G1996), .ZN(n805) );
  NOR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n925) );
  INV_X1 U904 ( .A(n925), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n807), .A2(n823), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n818), .A2(n812), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n826) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n874), .ZN(n921) );
  INV_X1 U910 ( .A(n812), .ZN(n815) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n813) );
  AND2_X1 U912 ( .A1(n859), .A2(n941), .ZN(n928) );
  NOR2_X1 U913 ( .A1(n813), .A2(n928), .ZN(n814) );
  NOR2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n921), .A2(n816), .ZN(n817) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n817), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n821) );
  OR2_X1 U918 ( .A1(n860), .A2(n820), .ZN(n933) );
  NAND2_X1 U919 ( .A1(n821), .A2(n933), .ZN(n822) );
  XOR2_X1 U920 ( .A(KEYINPUT99), .B(n822), .Z(n824) );
  NAND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U929 ( .A(KEYINPUT101), .B(n832), .Z(G188) );
  XOR2_X1 U930 ( .A(G69), .B(KEYINPUT102), .Z(G235) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G325) );
  XNOR2_X1 U932 ( .A(KEYINPUT103), .B(G325), .ZN(G261) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  NAND2_X1 U936 ( .A1(G124), .A2(n863), .ZN(n835) );
  XNOR2_X1 U937 ( .A(n835), .B(KEYINPUT44), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n836), .B(KEYINPUT106), .ZN(n838) );
  NAND2_X1 U939 ( .A1(G112), .A2(n864), .ZN(n837) );
  NAND2_X1 U940 ( .A1(n838), .A2(n837), .ZN(n842) );
  NAND2_X1 U941 ( .A1(G100), .A2(n867), .ZN(n840) );
  NAND2_X1 U942 ( .A1(G136), .A2(n868), .ZN(n839) );
  NAND2_X1 U943 ( .A1(n840), .A2(n839), .ZN(n841) );
  NOR2_X1 U944 ( .A1(n842), .A2(n841), .ZN(G162) );
  XNOR2_X1 U945 ( .A(G164), .B(G162), .ZN(n857) );
  XOR2_X1 U946 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n844) );
  XNOR2_X1 U947 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U949 ( .A(n845), .B(KEYINPUT111), .Z(n855) );
  NAND2_X1 U950 ( .A1(G103), .A2(n867), .ZN(n847) );
  NAND2_X1 U951 ( .A1(G139), .A2(n868), .ZN(n846) );
  NAND2_X1 U952 ( .A1(n847), .A2(n846), .ZN(n853) );
  NAND2_X1 U953 ( .A1(G127), .A2(n863), .ZN(n849) );
  NAND2_X1 U954 ( .A1(G115), .A2(n864), .ZN(n848) );
  NAND2_X1 U955 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U956 ( .A(KEYINPUT109), .B(n850), .ZN(n851) );
  XNOR2_X1 U957 ( .A(KEYINPUT47), .B(n851), .ZN(n852) );
  NOR2_X1 U958 ( .A1(n853), .A2(n852), .ZN(n914) );
  XNOR2_X1 U959 ( .A(n914), .B(KEYINPUT48), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U961 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U962 ( .A(n929), .B(n858), .ZN(n862) );
  XOR2_X1 U963 ( .A(n860), .B(n859), .Z(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n878) );
  NAND2_X1 U965 ( .A1(G130), .A2(n863), .ZN(n866) );
  NAND2_X1 U966 ( .A1(G118), .A2(n864), .ZN(n865) );
  NAND2_X1 U967 ( .A1(n866), .A2(n865), .ZN(n873) );
  NAND2_X1 U968 ( .A1(G106), .A2(n867), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G142), .A2(n868), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(n871), .B(KEYINPUT45), .Z(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(G160), .B(n876), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n879) );
  NOR2_X1 U976 ( .A1(G37), .A2(n879), .ZN(G395) );
  XOR2_X1 U977 ( .A(KEYINPUT112), .B(n880), .Z(n883) );
  XNOR2_X1 U978 ( .A(n881), .B(G301), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n885) );
  XOR2_X1 U980 ( .A(G286), .B(n969), .Z(n884) );
  XNOR2_X1 U981 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U982 ( .A1(G37), .A2(n886), .ZN(G397) );
  XOR2_X1 U983 ( .A(G1961), .B(G1956), .Z(n888) );
  XNOR2_X1 U984 ( .A(G1991), .B(G1986), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U986 ( .A(G1966), .B(G1971), .Z(n890) );
  XNOR2_X1 U987 ( .A(G1981), .B(G1976), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U989 ( .A(n892), .B(n891), .Z(n894) );
  XNOR2_X1 U990 ( .A(KEYINPUT41), .B(G2474), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U992 ( .A(KEYINPUT105), .B(n895), .ZN(n896) );
  XOR2_X1 U993 ( .A(n896), .B(G1996), .Z(G229) );
  XOR2_X1 U994 ( .A(G2096), .B(KEYINPUT43), .Z(n898) );
  XNOR2_X1 U995 ( .A(G2072), .B(KEYINPUT104), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(n899), .B(G2678), .Z(n901) );
  XNOR2_X1 U998 ( .A(G2067), .B(G2090), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U1000 ( .A(KEYINPUT42), .B(G2100), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G2078), .B(G2084), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(G227) );
  NOR2_X1 U1004 ( .A1(G395), .A2(G397), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(KEYINPUT114), .B(n906), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(n913), .A2(G401), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n907), .B(KEYINPUT113), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n908), .ZN(n909) );
  NOR2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n913), .ZN(G319) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1015 ( .A(G2072), .B(n914), .Z(n916) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(KEYINPUT116), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT50), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G2090), .B(G162), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(n919), .B(KEYINPUT115), .ZN(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n922), .Z(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n932) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n937), .ZN(n939) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(G29), .ZN(n1025) );
  XNOR2_X1 U1036 ( .A(KEYINPUT121), .B(G29), .ZN(n964) );
  XNOR2_X1 U1037 ( .A(G25), .B(n941), .ZN(n953) );
  XNOR2_X1 U1038 ( .A(KEYINPUT117), .B(G2072), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(n942), .B(G33), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G27), .B(n943), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(G28), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G26), .B(G2067), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT118), .B(G1996), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(G32), .B(n949), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT53), .B(n954), .ZN(n961) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G35), .ZN(n959) );
  XOR2_X1 U1051 ( .A(G34), .B(KEYINPUT120), .Z(n956) );
  XNOR2_X1 U1052 ( .A(G2084), .B(KEYINPUT54), .ZN(n955) );
  XNOR2_X1 U1053 ( .A(n956), .B(n955), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n957), .B(KEYINPUT119), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1057 ( .A(KEYINPUT55), .B(n962), .Z(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n965), .A2(G11), .ZN(n1023) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n991) );
  XNOR2_X1 U1061 ( .A(G1966), .B(G168), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(KEYINPUT57), .B(n968), .ZN(n989) );
  INV_X1 U1064 ( .A(G1341), .ZN(n992) );
  XNOR2_X1 U1065 ( .A(n969), .B(n992), .ZN(n981) );
  XNOR2_X1 U1066 ( .A(G1956), .B(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G1348), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1074 ( .A(G1961), .B(G171), .Z(n982) );
  XNOR2_X1 U1075 ( .A(KEYINPUT122), .B(n982), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT123), .B(n987), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n1021) );
  INV_X1 U1081 ( .A(G16), .ZN(n1019) );
  XNOR2_X1 U1082 ( .A(G19), .B(n992), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1956), .B(G20), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n999) );
  XOR2_X1 U1087 ( .A(KEYINPUT59), .B(G1348), .Z(n997) );
  XNOR2_X1 U1088 ( .A(G4), .B(n997), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1000), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT124), .B(n1003), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(n1004), .B(G5), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1016) );
  XNOR2_X1 U1096 ( .A(KEYINPUT125), .B(G1971), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(G1986), .B(KEYINPUT126), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(n1008), .B(G24), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1017), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1026), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

