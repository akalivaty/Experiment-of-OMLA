//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n570, new_n571, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n461), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OR3_X1    g047(.A1(new_n467), .A2(KEYINPUT65), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT65), .B1(new_n467), .B2(new_n472), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n471), .B1(new_n476), .B2(G2105), .ZN(G160));
  NOR2_X1   g052(.A1(new_n467), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(new_n461), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n461), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n479), .B(new_n481), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT66), .Z(G162));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n469), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n478), .A2(KEYINPUT4), .A3(G138), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n480), .A2(G126), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  NAND2_X1  g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT5), .A2(G543), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  OR2_X1    g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OR2_X1    g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n503), .A2(new_n495), .B1(new_n504), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n507), .B1(new_n504), .B2(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n501), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n506), .B1(new_n505), .B2(new_n510), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT69), .B(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(new_n508), .B2(new_n509), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(G50), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n502), .B1(new_n519), .B2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  XOR2_X1   g097(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n516), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n499), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(G89), .B2(new_n513), .ZN(G168));
  NAND2_X1  g104(.A1(G77), .A2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n498), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n513), .B2(G90), .ZN(G171));
  NAND2_X1  g111(.A1(new_n513), .A2(G81), .ZN(new_n537));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n498), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT72), .B(G43), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(G651), .B1(new_n516), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(new_n515), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n510), .A2(G53), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n516), .A2(KEYINPUT73), .A3(G53), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n501), .A2(KEYINPUT67), .A3(KEYINPUT6), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT67), .B1(new_n501), .B2(KEYINPUT6), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n496), .A2(new_n497), .B1(KEYINPUT6), .B2(new_n501), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT68), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n505), .A2(new_n506), .A3(new_n510), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G91), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n551), .A2(new_n552), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n498), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n555), .A2(new_n562), .A3(new_n564), .A4(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n560), .A2(new_n561), .ZN(new_n570));
  INV_X1    g145(.A(G90), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n533), .B(new_n534), .C1(new_n570), .C2(new_n571), .ZN(G301));
  NAND2_X1  g147(.A1(new_n513), .A2(G89), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n573), .A2(new_n526), .A3(new_n525), .A4(new_n527), .ZN(G286));
  NAND2_X1  g149(.A1(new_n513), .A2(G87), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n499), .A2(G74), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G49), .B2(new_n516), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n516), .A2(G48), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI221_X1 g156(.A(new_n579), .B1(new_n501), .B2(new_n580), .C1(new_n570), .C2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n501), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n513), .A2(G85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n516), .A2(G47), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G66), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n498), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n594));
  OAI21_X1  g169(.A(G54), .B1(new_n516), .B2(new_n594), .ZN(new_n595));
  NOR3_X1   g170(.A1(new_n558), .A2(KEYINPUT75), .A3(new_n515), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n560), .A2(G92), .A3(new_n561), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n560), .A2(KEYINPUT10), .A3(G92), .A4(new_n561), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n589), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NAND2_X1  g180(.A1(G299), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n605), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n543), .A2(new_n605), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n600), .A2(new_n601), .ZN(new_n612));
  INV_X1    g187(.A(new_n597), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n611), .B1(new_n615), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n468), .A2(new_n463), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G2100), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n478), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n480), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n461), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(G2096), .Z(new_n630));
  NAND3_X1  g205(.A1(new_n623), .A2(new_n624), .A3(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT78), .Z(new_n647));
  OAI21_X1  g222(.A(G14), .B1(new_n643), .B2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT79), .ZN(G401));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT17), .Z(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(new_n653), .B2(new_n651), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT80), .Z(new_n660));
  NAND3_X1  g235(.A1(new_n656), .A2(new_n653), .A3(new_n651), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT18), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n653), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n652), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G229));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G35), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G162), .B2(new_n686), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT29), .Z(new_n689));
  INV_X1    g264(.A(G2090), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT97), .ZN(new_n692));
  NAND2_X1  g267(.A1(G115), .A2(G2104), .ZN(new_n693));
  INV_X1    g268(.A(G127), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n467), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n461), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n697), .B1(new_n696), .B2(new_n695), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT25), .Z(new_n700));
  AOI21_X1  g275(.A(KEYINPUT88), .B1(new_n478), .B2(G139), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n478), .A2(KEYINPUT88), .A3(G139), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n698), .B(new_n700), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G33), .B(new_n705), .S(G29), .Z(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G2072), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT91), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n692), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n689), .A2(new_n690), .ZN(new_n710));
  INV_X1    g285(.A(G1348), .ZN(new_n711));
  NOR2_X1   g286(.A1(G4), .A2(G16), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n602), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n710), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n706), .A2(G2072), .B1(G1348), .B2(new_n713), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n686), .A2(G26), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT28), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n480), .A2(G128), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n461), .A2(G116), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G140), .B2(new_n478), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT87), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(G29), .ZN(new_n725));
  INV_X1    g300(.A(G2067), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(G19), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n543), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G1341), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n686), .A2(G27), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G164), .B2(new_n686), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G171), .A2(new_n728), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G5), .B2(new_n728), .ZN(new_n738));
  INV_X1    g313(.A(G1961), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n731), .A2(G1341), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n732), .A2(new_n736), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n686), .A2(G32), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n480), .A2(G129), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT93), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT26), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n745), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(new_n686), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n727), .A2(new_n742), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n686), .B1(new_n756), .B2(G34), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n756), .B2(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G160), .B2(G29), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2084), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT92), .Z(new_n761));
  NOR2_X1   g336(.A1(new_n759), .A2(G2084), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n715), .A2(new_n716), .A3(new_n755), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT30), .B(G28), .ZN(new_n766));
  OR2_X1    g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n766), .A2(new_n686), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI221_X1 g344(.A(new_n769), .B1(new_n686), .B2(new_n629), .C1(new_n738), .C2(new_n739), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n728), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n728), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1966), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n770), .A2(KEYINPUT95), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(KEYINPUT95), .B1(new_n770), .B2(new_n773), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n728), .A2(G20), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT23), .ZN(new_n777));
  AND4_X1   g352(.A1(new_n555), .A2(new_n562), .A3(new_n564), .A4(new_n568), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n728), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n775), .A2(new_n781), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n709), .A2(new_n765), .A3(new_n774), .A4(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G6), .B(G305), .S(G16), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  INV_X1    g360(.A(G1981), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n728), .A2(G22), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT85), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n728), .ZN(new_n790));
  INV_X1    g365(.A(G1971), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n728), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n728), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT83), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT33), .B(G1976), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT84), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n787), .A2(new_n792), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT82), .B(KEYINPUT34), .Z(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n802), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G24), .ZN(new_n805));
  INV_X1    g380(.A(G290), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G16), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G1986), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n686), .A2(G25), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT81), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n478), .A2(G131), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n480), .A2(G119), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n461), .A2(G107), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n811), .B(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n810), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n808), .A2(KEYINPUT86), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G1986), .B2(new_n807), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n803), .A2(KEYINPUT36), .A3(new_n804), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n803), .A2(new_n804), .A3(new_n821), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT36), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n783), .A2(new_n822), .A3(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  AOI22_X1  g402(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(new_n501), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT98), .B(G93), .Z(new_n831));
  NAND3_X1  g406(.A1(new_n560), .A2(new_n561), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n516), .A2(G55), .ZN(new_n833));
  AND3_X1   g408(.A1(new_n832), .A2(KEYINPUT99), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT99), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(KEYINPUT100), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n838), .B(new_n830), .C1(new_n834), .C2(new_n835), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n544), .B1(new_n837), .B2(new_n839), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n836), .A2(new_n543), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n614), .A2(new_n609), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n846), .A2(new_n847), .ZN(new_n852));
  OR3_X1    g427(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n849), .B2(new_n852), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n853), .A2(KEYINPUT39), .A3(new_n854), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n857), .A2(KEYINPUT101), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT101), .B1(new_n857), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n843), .B1(new_n859), .B2(new_n860), .ZN(G145));
  XNOR2_X1  g436(.A(new_n705), .B(new_n750), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n724), .B(new_n493), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n815), .B(KEYINPUT103), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n619), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n478), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n480), .A2(G130), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n872), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n864), .A2(KEYINPUT104), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(KEYINPUT104), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n878), .A3(new_n874), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n876), .B1(new_n864), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G160), .B(new_n629), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G162), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n876), .B(new_n883), .C1(new_n864), .C2(new_n880), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n889), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G395));
  XNOR2_X1  g468(.A(G303), .B(new_n794), .ZN(new_n894));
  XNOR2_X1  g469(.A(G305), .B(KEYINPUT107), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(G290), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(new_n896), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT108), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n897), .A2(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n901), .ZN(new_n904));
  NAND2_X1  g479(.A1(KEYINPUT108), .A2(KEYINPUT42), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n846), .B(new_n615), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n602), .A2(new_n778), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n602), .A2(new_n778), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT41), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n614), .A2(G299), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n602), .A2(new_n778), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n909), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n910), .A2(new_n911), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT106), .B1(new_n918), .B2(new_n913), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n908), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n908), .B1(new_n911), .B2(new_n910), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n907), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n907), .B1(new_n921), .B2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(G868), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n840), .A2(new_n605), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(G295));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n926), .ZN(G331));
  XOR2_X1   g503(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n832), .A2(new_n833), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT99), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n832), .A2(KEYINPUT99), .A3(new_n833), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n838), .B1(new_n935), .B2(new_n830), .ZN(new_n936));
  INV_X1    g511(.A(new_n839), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n543), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n845), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n940));
  NAND2_X1  g515(.A1(G171), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G301), .A2(KEYINPUT110), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n941), .A2(new_n942), .A3(G168), .ZN(new_n943));
  NAND3_X1  g518(.A1(G286), .A2(KEYINPUT110), .A3(G301), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n938), .A2(new_n939), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n844), .B2(new_n845), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n918), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT112), .A4(new_n918), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n948), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n953), .A2(KEYINPUT111), .A3(new_n920), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT111), .B1(new_n953), .B2(new_n920), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n951), .B(new_n952), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(new_n903), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n951), .A2(new_n952), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n899), .C1(new_n955), .C2(new_n954), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n930), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n953), .B1(new_n916), .B2(new_n912), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n949), .ZN(new_n962));
  AOI21_X1  g537(.A(G37), .B1(new_n962), .B2(new_n903), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n963), .B(new_n930), .C1(new_n956), .C2(new_n903), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n929), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n959), .A2(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n957), .A2(new_n930), .A3(new_n959), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(G397));
  INV_X1    g546(.A(G1384), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n493), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G160), .A2(G40), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n977), .A2(KEYINPUT114), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(KEYINPUT114), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n724), .B(new_n726), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n750), .B(G1996), .Z(new_n982));
  AOI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n980), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n815), .A2(new_n818), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n815), .A2(new_n818), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  AND2_X1   g566(.A1(G290), .A2(G1986), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT115), .Z(new_n994));
  AND2_X1   g569(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT118), .B(KEYINPUT50), .Z(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(G40), .B(G160), .C1(new_n973), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT119), .B(new_n999), .C1(new_n493), .C2(new_n972), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT119), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1348), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT124), .ZN(new_n1006));
  AND2_X1   g581(.A1(G160), .A2(G40), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n493), .A2(new_n972), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2067), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1005), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n976), .B1(new_n1008), .B2(new_n996), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n973), .A2(new_n1002), .A3(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1004), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n711), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1010), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT124), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT60), .B(new_n614), .C1(new_n1011), .C2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1007), .B1(new_n1008), .B2(new_n996), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n780), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n976), .B1(new_n973), .B2(new_n974), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n493), .A2(new_n1023), .A3(KEYINPUT45), .A4(new_n972), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT117), .B1(new_n973), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT56), .B(G2072), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1022), .A2(new_n1024), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1021), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT123), .B(KEYINPUT57), .ZN(new_n1030));
  XNOR2_X1  g605(.A(G299), .B(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1021), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(KEYINPUT61), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT61), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1026), .A2(new_n1007), .A3(new_n1024), .A4(new_n975), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n976), .A2(new_n973), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT58), .B(G1341), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1039), .A2(G1996), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n544), .A2(KEYINPUT126), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1042), .A2(KEYINPUT59), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT59), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND4_X1   g621(.A1(new_n1018), .A2(new_n1035), .A3(new_n1038), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT60), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1006), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1015), .A2(KEYINPUT124), .A3(new_n1016), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1048), .A2(new_n602), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1050), .A3(new_n602), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT125), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1049), .A2(new_n1050), .A3(new_n1056), .A4(new_n602), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1057), .A3(new_n1033), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1047), .A2(new_n1053), .B1(new_n1058), .B2(new_n1034), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1022), .A2(new_n735), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT127), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT127), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1065), .A3(new_n1062), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1064), .A2(new_n1066), .B1(new_n739), .B2(new_n1014), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1007), .B(KEYINPUT122), .C1(new_n1008), .C2(KEYINPUT45), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT45), .B1(new_n493), .B2(new_n972), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(new_n976), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n973), .A2(new_n974), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  OR3_X1    g648(.A1(new_n1073), .A2(new_n1062), .A3(G2078), .ZN(new_n1074));
  AOI21_X1  g649(.A(G301), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1014), .A2(new_n739), .ZN(new_n1076));
  OR3_X1    g651(.A1(new_n1039), .A2(new_n1062), .A3(G2078), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1061), .A2(new_n1065), .A3(new_n1062), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1065), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1076), .B(new_n1077), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1060), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1039), .A2(new_n791), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(G2090), .B2(new_n1014), .ZN(new_n1084));
  NAND3_X1  g659(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1084), .B(G8), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1040), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n794), .A2(G1976), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n794), .A2(G1976), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1090), .A2(KEYINPUT120), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1093), .A2(KEYINPUT120), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(new_n1090), .C1(KEYINPUT52), .C2(new_n1091), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G305), .B(new_n786), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT49), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT121), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1009), .A2(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1095), .A2(new_n1097), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1087), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n996), .B1(new_n493), .B2(new_n972), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1020), .A2(new_n976), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n791), .A2(new_n1039), .B1(new_n1107), .B2(new_n690), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1105), .B(new_n1085), .C1(new_n1108), .C2(new_n1089), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1088), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1966), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1073), .A2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n998), .A2(new_n1003), .A3(new_n1000), .ZN(new_n1113));
  INV_X1    g688(.A(G2084), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1115), .A3(G168), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G8), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1111), .A2(new_n1073), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(G168), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT51), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1089), .B1(new_n1118), .B2(G168), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1110), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1060), .B1(new_n1080), .B2(G171), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1074), .B(new_n1076), .C1(new_n1079), .C2(new_n1078), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(G171), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1082), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1059), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G286), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1122), .B1(new_n1121), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT62), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1126), .A2(G171), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n1110), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1120), .A2(new_n1137), .A3(new_n1123), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1134), .A2(new_n1136), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1118), .A2(new_n1089), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G286), .A2(KEYINPUT63), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1109), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1088), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1104), .ZN(new_n1144));
  AOI211_X1 g719(.A(G1976), .B(G288), .C1(new_n1103), .C2(new_n1101), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G305), .A2(G1981), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1113), .A2(new_n690), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1105), .A2(new_n1085), .A3(new_n1083), .A4(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1104), .A2(new_n1140), .A3(G168), .A4(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1147), .A2(new_n1090), .B1(new_n1150), .B2(KEYINPUT63), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1139), .A2(new_n1144), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n995), .B1(new_n1129), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n986), .A2(new_n991), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT48), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n990), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n985), .A2(new_n987), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n724), .A2(G2067), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n980), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n980), .B1(new_n751), .B2(new_n981), .ZN(new_n1160));
  OR3_X1    g735(.A1(new_n980), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT46), .B1(new_n980), .B2(G1996), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1163), .B(KEYINPUT47), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1156), .A2(new_n1159), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g741(.A1(new_n960), .A2(new_n965), .ZN(new_n1168));
  NOR4_X1   g742(.A1(new_n649), .A2(G229), .A3(new_n459), .A4(G227), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n888), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1168), .A2(new_n1170), .ZN(G308));
  OAI211_X1 g745(.A(new_n888), .B(new_n1169), .C1(new_n960), .C2(new_n965), .ZN(G225));
endmodule


