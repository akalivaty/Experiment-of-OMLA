//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(G134), .B2(new_n192), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n189), .A2(KEYINPUT11), .A3(G137), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n188), .B(new_n190), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT64), .B1(new_n192), .B2(G134), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n189), .A3(G137), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n196), .A2(new_n198), .B1(G134), .B2(new_n192), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n188), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n196), .A2(new_n198), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n189), .A2(G137), .ZN(new_n204));
  OAI21_X1  g018(.A(G131), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT67), .A3(new_n195), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n208), .A2(KEYINPUT1), .A3(G146), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n212), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n215), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n217), .B1(new_n222), .B2(new_n207), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n216), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT68), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n202), .A2(new_n206), .A3(new_n221), .A4(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT2), .B(G113), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G116), .B(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(G116), .B(G119), .Z(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n227), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G143), .B(G146), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT0), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(new_n207), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT0), .B(G128), .Z(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n195), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT11), .B1(new_n189), .B2(G137), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n191), .A2(new_n192), .A3(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n188), .B1(new_n243), .B2(new_n190), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n239), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n226), .A2(new_n234), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT71), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT71), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n226), .A2(new_n245), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n248), .B(new_n250), .C1(new_n234), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT28), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT28), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n246), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(G237), .A2(G953), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G210), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n259), .B(KEYINPUT27), .Z(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n187), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT65), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n200), .B2(new_n219), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n224), .A2(new_n205), .A3(KEYINPUT65), .A4(new_n195), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n245), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n233), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n254), .B1(new_n246), .B2(new_n270), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n271), .A2(new_n255), .A3(new_n262), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n269), .A2(KEYINPUT66), .A3(new_n273), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n226), .A2(KEYINPUT30), .A3(new_n245), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n276), .A2(new_n233), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n246), .ZN(new_n280));
  AOI211_X1 g094(.A(KEYINPUT29), .B(new_n272), .C1(new_n262), .C2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(G472), .B1(new_n265), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n278), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT66), .B1(new_n269), .B2(new_n273), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n285), .A2(new_n234), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n246), .A2(new_n263), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n288), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(KEYINPUT69), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(KEYINPUT31), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n279), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n262), .B1(new_n271), .B2(new_n255), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n283), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n298), .ZN(new_n300));
  AOI211_X1 g114(.A(KEYINPUT32), .B(new_n300), .C1(new_n292), .C2(new_n296), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n282), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G104), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT3), .B1(new_n305), .B2(G107), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n307));
  INV_X1    g121(.A(G107), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(G104), .ZN(new_n309));
  INV_X1    g123(.A(G101), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(G107), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n306), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n305), .A2(G107), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n308), .A2(G104), .ZN(new_n314));
  OAI21_X1  g128(.A(G101), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n221), .A2(new_n225), .A3(KEYINPUT10), .A4(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n306), .A2(new_n309), .A3(new_n311), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT4), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G101), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n318), .A2(G101), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n312), .A2(KEYINPUT4), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n239), .B(new_n320), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n216), .A2(KEYINPUT75), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n223), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n316), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n317), .A2(new_n323), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n240), .A2(new_n244), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(G110), .B(G140), .Z(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT74), .ZN(new_n336));
  INV_X1    g150(.A(G227), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G953), .ZN(new_n338));
  XOR2_X1   g152(.A(new_n336), .B(new_n338), .Z(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n334), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n331), .A2(new_n333), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n312), .A2(new_n315), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(new_n216), .A3(new_n223), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n328), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT12), .A3(new_n333), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n212), .A2(new_n218), .A3(new_n326), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n350), .B2(new_n324), .ZN(new_n351));
  INV_X1    g165(.A(new_n346), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT76), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n328), .A2(new_n354), .A3(new_n346), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT12), .B1(new_n356), .B2(new_n333), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n349), .B1(new_n357), .B2(KEYINPUT77), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n332), .B1(new_n353), .B2(new_n355), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(KEYINPUT12), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n334), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(G469), .B(new_n344), .C1(new_n362), .C2(new_n339), .ZN(new_n363));
  NAND2_X1  g177(.A1(G469), .A2(G902), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT78), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n366));
  INV_X1    g180(.A(new_n334), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n328), .A2(new_n354), .A3(new_n346), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n354), .B1(new_n328), .B2(new_n346), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n333), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(KEYINPUT77), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n348), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT77), .B1(new_n370), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n367), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n343), .B1(new_n375), .B2(new_n340), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n366), .B(G469), .C1(new_n376), .C2(G902), .ZN(new_n377));
  INV_X1    g191(.A(G469), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n361), .A2(new_n372), .A3(new_n348), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n379), .A2(new_n341), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n339), .B1(new_n367), .B2(new_n342), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n378), .B(new_n187), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n365), .A2(new_n377), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G221), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n386), .B2(new_n187), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G113), .B(G122), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n389), .B(new_n305), .ZN(new_n390));
  INV_X1    g204(.A(G237), .ZN(new_n391));
  INV_X1    g205(.A(G953), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G214), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n208), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n258), .A2(G143), .A3(G214), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT18), .A3(G131), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G125), .B(G140), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n400), .A2(new_n210), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n210), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n401), .B2(new_n403), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n397), .B(new_n399), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n395), .ZN(new_n407));
  AOI21_X1  g221(.A(G143), .B1(new_n258), .B2(G214), .ZN(new_n408));
  OAI21_X1  g222(.A(G131), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n394), .A2(new_n188), .A3(new_n395), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(KEYINPUT83), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT82), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n409), .B2(new_n410), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n400), .A2(KEYINPUT16), .ZN(new_n416));
  INV_X1    g230(.A(G125), .ZN(new_n417));
  OR3_X1    g231(.A1(new_n417), .A2(KEYINPUT16), .A3(G140), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n210), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(G146), .A3(new_n418), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n396), .A2(KEYINPUT82), .A3(KEYINPUT17), .A4(G131), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n415), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n390), .B(new_n406), .C1(new_n413), .C2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n406), .B1(new_n413), .B2(new_n423), .ZN(new_n426));
  INV_X1    g240(.A(new_n390), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT84), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n426), .A2(new_n430), .A3(new_n427), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n425), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G475), .B1(new_n432), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n400), .A2(new_n434), .A3(KEYINPUT19), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(new_n400), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n210), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n409), .A2(new_n411), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n421), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n406), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n427), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n424), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n443), .B2(new_n445), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n433), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT8), .Z(new_n451));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n452));
  INV_X1    g266(.A(G119), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n453), .A3(G116), .ZN(new_n454));
  OAI211_X1 g268(.A(G113), .B(new_n454), .C1(new_n231), .C2(new_n452), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n230), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n345), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n316), .A2(new_n230), .A3(new_n455), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n451), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n392), .A2(G224), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n460), .A2(KEYINPUT7), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n237), .B(G125), .C1(new_n235), .C2(new_n238), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n223), .A2(new_n417), .A3(new_n216), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n462), .A2(new_n463), .A3(new_n461), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n459), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n233), .A2(new_n320), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n321), .A2(new_n322), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n458), .B(new_n450), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n458), .B1(new_n467), .B2(new_n468), .ZN(new_n471));
  INV_X1    g285(.A(new_n450), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n462), .A2(new_n463), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n460), .B(KEYINPUT79), .Z(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n478), .A3(new_n472), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G210), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n470), .A2(new_n480), .A3(new_n482), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(G234), .A2(G237), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(G952), .A3(new_n392), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(G902), .A3(G953), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT88), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT21), .B(G898), .Z(new_n491));
  OAI21_X1  g305(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G214), .B1(G237), .B2(G902), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n386), .A2(G217), .A3(new_n392), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(new_n207), .B2(G143), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n208), .A2(KEYINPUT85), .A3(G128), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n500), .A2(new_n501), .B1(new_n207), .B2(G143), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(KEYINPUT13), .A3(new_n499), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n189), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n504), .A2(KEYINPUT86), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(KEYINPUT86), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n500), .B(new_n189), .C1(G128), .C2(new_n208), .ZN(new_n507));
  XNOR2_X1  g321(.A(G116), .B(G122), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n508), .A2(G107), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(G107), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n507), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n500), .B1(G128), .B2(new_n208), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G134), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n507), .ZN(new_n515));
  INV_X1    g329(.A(G116), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n516), .A2(G122), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n308), .B1(new_n517), .B2(KEYINPUT14), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n508), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n496), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n512), .A2(new_n520), .A3(new_n496), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n187), .ZN(new_n525));
  INV_X1    g339(.A(G478), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT87), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n524), .A2(new_n187), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n449), .A2(new_n494), .A3(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n383), .A2(new_n388), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(G234), .ZN(new_n538));
  OAI21_X1  g352(.A(G217), .B1(new_n538), .B2(G902), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n453), .A2(G128), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT23), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n207), .A2(G119), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT73), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n541), .B(new_n543), .Z(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n542), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT24), .B(G110), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI22_X1  g362(.A1(new_n544), .A2(G110), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n421), .A3(new_n403), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n544), .A2(G110), .B1(new_n546), .B2(new_n548), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n420), .A2(new_n421), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT22), .B(G137), .ZN(new_n555));
  NOR3_X1   g369(.A1(new_n384), .A2(new_n538), .A3(G953), .ZN(new_n556));
  XOR2_X1   g370(.A(new_n555), .B(new_n556), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n553), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n557), .ZN(new_n561));
  AOI21_X1  g375(.A(G902), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT25), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n539), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n563), .B2(new_n562), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n559), .A2(new_n561), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n538), .B2(G217), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n282), .B(KEYINPUT72), .C1(new_n299), .C2(new_n301), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n304), .A2(new_n537), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(G101), .ZN(G3));
  AND2_X1   g387(.A1(new_n383), .A2(new_n388), .ZN(new_n574));
  INV_X1    g388(.A(G472), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n297), .B2(new_n187), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n300), .B1(new_n292), .B2(new_n296), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n576), .A2(new_n569), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n579), .B(KEYINPUT89), .Z(new_n580));
  INV_X1    g394(.A(G475), .ZN(new_n581));
  INV_X1    g395(.A(new_n431), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n430), .B1(new_n426), .B2(new_n427), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n424), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n581), .B1(new_n584), .B2(new_n187), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n446), .A2(new_n447), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n523), .ZN(new_n588));
  OAI211_X1 g402(.A(KEYINPUT91), .B(KEYINPUT33), .C1(new_n588), .C2(new_n521), .ZN(new_n589));
  OR2_X1    g403(.A1(KEYINPUT91), .A2(KEYINPUT33), .ZN(new_n590));
  NAND2_X1  g404(.A1(KEYINPUT91), .A2(KEYINPUT33), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n522), .A2(new_n523), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n526), .A2(G902), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n593), .A2(new_n594), .B1(new_n526), .B2(new_n525), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n486), .ZN(new_n597));
  INV_X1    g411(.A(new_n493), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT90), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT90), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n486), .A2(new_n600), .A3(new_n493), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n492), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n580), .A2(new_n596), .A3(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT34), .B(G104), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  AOI21_X1  g421(.A(new_n449), .B1(new_n532), .B2(new_n534), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n580), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT92), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT35), .B(G107), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  NOR2_X1   g428(.A1(new_n576), .A2(new_n577), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n383), .A2(new_n388), .A3(new_n536), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n558), .A2(KEYINPUT36), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n554), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n560), .B1(KEYINPUT36), .B2(new_n558), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n567), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(KEYINPUT93), .A3(new_n567), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n626), .A2(new_n565), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n616), .A2(new_n617), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT37), .B(G110), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  NAND2_X1  g444(.A1(new_n626), .A2(new_n565), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n383), .A2(new_n388), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n488), .B(KEYINPUT94), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n490), .B2(G900), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n608), .A2(new_n602), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n304), .A2(new_n632), .A3(new_n571), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  XNOR2_X1  g451(.A(new_n634), .B(KEYINPUT39), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n574), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT40), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n299), .A2(new_n301), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n289), .A2(new_n291), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n262), .B2(new_n252), .ZN(new_n643));
  OAI21_X1  g457(.A(G472), .B1(new_n643), .B2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n486), .B(KEYINPUT38), .Z(new_n647));
  NAND4_X1  g461(.A1(new_n627), .A2(new_n493), .A3(new_n449), .A4(new_n535), .ZN(new_n648));
  NOR4_X1   g462(.A1(new_n640), .A2(new_n646), .A3(new_n647), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n208), .ZN(G45));
  AND3_X1   g464(.A1(new_n602), .A2(new_n596), .A3(new_n634), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n304), .A2(new_n632), .A3(new_n571), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT95), .B(G146), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G48));
  AOI21_X1  g468(.A(new_n381), .B1(new_n379), .B2(new_n341), .ZN(new_n655));
  OAI21_X1  g469(.A(G469), .B1(new_n655), .B2(G902), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n382), .A2(new_n656), .A3(new_n388), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT96), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n304), .A2(new_n570), .A3(new_n659), .A4(new_n571), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n604), .A2(new_n596), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT41), .B(G113), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G15));
  AND3_X1   g478(.A1(new_n304), .A2(new_n570), .A3(new_n571), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT97), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n666), .A3(new_n610), .A4(new_n659), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT97), .B1(new_n660), .B2(new_n609), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G116), .ZN(G18));
  INV_X1    g484(.A(new_n657), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n671), .A2(new_n602), .A3(new_n631), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n449), .A2(new_n535), .ZN(new_n673));
  AND2_X1   g487(.A1(new_n673), .A2(new_n492), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n304), .A2(new_n672), .A3(new_n571), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G119), .ZN(G21));
  OAI21_X1  g490(.A(new_n535), .B1(new_n585), .B2(new_n586), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT99), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n449), .A2(KEYINPUT99), .A3(new_n535), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n492), .A2(new_n602), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n292), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n263), .B1(new_n253), .B2(new_n256), .ZN(new_n683));
  OAI21_X1  g497(.A(KEYINPUT98), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n257), .A2(new_n262), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n686), .A3(new_n292), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n684), .A2(new_n294), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n576), .B1(new_n688), .B2(new_n298), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n681), .A2(new_n689), .A3(new_n659), .A4(new_n570), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n596), .B2(new_n634), .ZN(new_n693));
  INV_X1    g507(.A(new_n634), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n587), .A2(new_n595), .A3(KEYINPUT100), .A4(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n696), .A2(new_n672), .A3(new_n689), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  XOR2_X1   g512(.A(new_n364), .B(KEYINPUT101), .Z(new_n699));
  NAND3_X1  g513(.A1(new_n382), .A2(new_n363), .A3(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n486), .A2(new_n387), .A3(new_n598), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n665), .A2(KEYINPUT102), .A3(new_n696), .A4(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n304), .A2(new_n570), .A3(new_n571), .A4(new_n702), .ZN(new_n705));
  INV_X1    g519(.A(new_n696), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n302), .A2(new_n710), .A3(new_n570), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n710), .B1(new_n302), .B2(new_n570), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n696), .A2(new_n702), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(KEYINPUT42), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  AND2_X1   g531(.A1(new_n608), .A2(new_n634), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n705), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n189), .ZN(G36));
  NOR2_X1   g535(.A1(new_n486), .A2(new_n598), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT107), .Z(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n726));
  AOI211_X1 g540(.A(new_n595), .B(new_n449), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n616), .A3(new_n631), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n724), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n729), .A2(KEYINPUT44), .A3(new_n616), .A4(new_n631), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n733), .B1(new_n732), .B2(new_n734), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n376), .B(KEYINPUT45), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n378), .ZN(new_n739));
  INV_X1    g553(.A(new_n699), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n382), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n388), .A3(new_n638), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT105), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n737), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n388), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT47), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n304), .A2(new_n571), .ZN(new_n752));
  INV_X1    g566(.A(new_n596), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n694), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n752), .A2(new_n569), .A3(new_n754), .A4(new_n722), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n755), .B(KEYINPUT109), .Z(new_n756));
  NAND2_X1  g570(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G140), .ZN(G42));
  NAND3_X1  g572(.A1(new_n570), .A2(new_n388), .A3(new_n493), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT110), .ZN(new_n760));
  INV_X1    g574(.A(new_n595), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n587), .A3(new_n761), .A4(new_n647), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n382), .A2(new_n656), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n762), .B1(KEYINPUT49), .B2(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n764), .B(new_n646), .C1(KEYINPUT49), .C2(new_n763), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n690), .B(new_n675), .C1(new_n660), .C2(new_n661), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n669), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n494), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n574), .A2(new_n578), .A3(new_n769), .A4(new_n596), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n572), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n579), .A2(new_n494), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n628), .B1(new_n774), .B2(new_n608), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n572), .A2(KEYINPUT111), .A3(new_n770), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n602), .A2(new_n679), .A3(new_n680), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n627), .A2(new_n700), .A3(new_n388), .A4(new_n634), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n645), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n636), .A2(new_n652), .A3(new_n697), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n779), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n688), .A2(new_n298), .ZN(new_n789));
  INV_X1    g603(.A(new_n576), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n627), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n714), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n673), .A2(new_n634), .A3(new_n722), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n304), .A2(new_n632), .A3(new_n571), .A4(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n793), .B(new_n795), .C1(new_n719), .C2(new_n705), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n709), .B2(new_n715), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n636), .A2(new_n697), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT112), .A3(new_n652), .A4(new_n783), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n784), .A2(new_n785), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(KEYINPUT52), .A3(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n778), .A2(new_n788), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n784), .A2(KEYINPUT52), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n800), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n805), .B1(new_n806), .B2(new_n779), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n778), .A4(new_n797), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT113), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n803), .A2(new_n809), .A3(new_n812), .A4(KEYINPUT54), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n768), .A2(KEYINPUT115), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n766), .B1(new_n667), .B2(new_n668), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n777), .A2(new_n808), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n814), .A2(new_n797), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n807), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n788), .A2(new_n801), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n773), .A2(new_n776), .A3(new_n775), .ZN(new_n824));
  INV_X1    g638(.A(new_n796), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n716), .A2(new_n824), .A3(new_n815), .A4(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n822), .B(new_n808), .C1(new_n823), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n822), .B1(new_n802), .B2(new_n808), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n821), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n811), .B(new_n813), .C1(new_n830), .C2(KEYINPUT54), .ZN(new_n831));
  INV_X1    g645(.A(new_n633), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n729), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n570), .A3(new_n689), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n671), .A2(new_n598), .A3(new_n647), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT50), .ZN(new_n837));
  INV_X1    g651(.A(new_n488), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n701), .A2(new_n382), .A3(new_n656), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n646), .A2(new_n570), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n449), .A3(new_n761), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n833), .A2(new_n839), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n842), .B2(new_n792), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT51), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n750), .B1(new_n388), .B2(new_n763), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n724), .B(new_n834), .C1(new_n846), .C2(KEYINPUT116), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(KEYINPUT116), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n834), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n846), .A2(new_n723), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT51), .B1(new_n844), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n392), .A2(G952), .ZN(new_n853));
  INV_X1    g667(.A(new_n840), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n596), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n671), .A2(new_n602), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n842), .A2(new_n713), .ZN(new_n857));
  NOR2_X1   g671(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n857), .B(new_n858), .Z(new_n859));
  AND2_X1   g673(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n860));
  OAI221_X1 g674(.A(new_n855), .B1(new_n856), .B2(new_n834), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n831), .A2(new_n849), .A3(new_n852), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(G952), .A2(G953), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n765), .B1(new_n862), .B2(new_n863), .ZN(G75));
  NOR2_X1   g678(.A1(new_n819), .A2(new_n820), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n808), .B1(new_n823), .B2(new_n826), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT114), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n867), .B2(new_n827), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n187), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(G210), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n474), .A2(new_n479), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n477), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT55), .Z(new_n874));
  AND3_X1   g688(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n874), .B1(new_n870), .B2(new_n871), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n392), .A2(G952), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G51));
  XOR2_X1   g692(.A(new_n699), .B(KEYINPUT57), .Z(new_n879));
  NOR2_X1   g693(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n868), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n655), .B(KEYINPUT118), .Z(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n869), .A2(new_n739), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n877), .B1(new_n885), .B2(new_n886), .ZN(G54));
  INV_X1    g701(.A(new_n877), .ZN(new_n888));
  AND2_X1   g702(.A1(KEYINPUT58), .A2(G475), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n869), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n443), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  AOI211_X1 g708(.A(KEYINPUT119), .B(new_n443), .C1(new_n869), .C2(new_n889), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n831), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n593), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT120), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n903), .B(new_n593), .C1(new_n831), .C2(new_n899), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n898), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n880), .B2(new_n882), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n888), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n902), .A2(new_n904), .A3(new_n907), .ZN(G63));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT121), .Z(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT60), .Z(new_n911));
  NAND2_X1  g725(.A1(new_n830), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n566), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n877), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n915));
  INV_X1    g729(.A(new_n911), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n867), .A2(new_n827), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n821), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT122), .B1(new_n918), .B2(new_n621), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  INV_X1    g734(.A(new_n621), .ZN(new_n921));
  NOR4_X1   g735(.A1(new_n868), .A2(new_n920), .A3(new_n921), .A4(new_n916), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n914), .B(new_n915), .C1(new_n919), .C2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n830), .A2(new_n621), .A3(new_n911), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n920), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n830), .A2(KEYINPUT122), .A3(new_n621), .A4(new_n911), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n915), .B1(new_n928), .B2(new_n914), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n924), .A2(new_n929), .ZN(G66));
  NAND3_X1  g744(.A1(new_n491), .A2(G224), .A3(G953), .ZN(new_n931));
  INV_X1    g745(.A(new_n778), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(G953), .ZN(new_n933));
  INV_X1    g747(.A(G898), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n872), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  AOI21_X1  g750(.A(new_n392), .B1(G227), .B2(G900), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT126), .Z(new_n938));
  NOR2_X1   g752(.A1(new_n392), .A2(G900), .ZN(new_n939));
  INV_X1    g753(.A(new_n780), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n713), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n746), .B1(new_n737), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n720), .B1(new_n751), .B2(new_n756), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n798), .A2(new_n652), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n942), .A2(new_n943), .A3(new_n716), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n939), .B1(new_n946), .B2(new_n392), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n285), .A2(new_n286), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(new_n437), .Z(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n938), .B1(new_n950), .B2(KEYINPUT125), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n952));
  OR3_X1    g766(.A1(new_n649), .A2(new_n952), .A3(new_n944), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n952), .B1(new_n649), .B2(new_n944), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n608), .A2(new_n596), .ZN(new_n956));
  OR2_X1    g770(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(KEYINPUT124), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n957), .A2(new_n722), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n959), .A2(new_n665), .A3(new_n574), .A4(new_n638), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n955), .A2(new_n747), .A3(new_n757), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n392), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n949), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(new_n947), .B2(new_n949), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n951), .B(new_n964), .ZN(G72));
  NAND2_X1  g779(.A1(G472), .A2(G902), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT63), .Z(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n961), .B2(new_n932), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n263), .A3(new_n280), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT127), .Z(new_n970));
  OAI21_X1  g784(.A(new_n967), .B1(new_n946), .B2(new_n932), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n280), .A2(new_n263), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n877), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n803), .A2(new_n809), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n280), .A2(new_n262), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n967), .B1(new_n642), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n973), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n970), .A2(new_n978), .ZN(G57));
endmodule


