//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n454), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT68), .Z(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n453), .B2(G2106), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(G101), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n467), .A2(new_n469), .A3(new_n462), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n470), .A2(G136), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n462), .A2(G112), .ZN(new_n475));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n467), .A2(new_n469), .A3(G2105), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n477), .B1(G124), .B2(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(G162));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n460), .A2(new_n483), .A3(G138), .A4(new_n462), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n470), .A2(KEYINPUT72), .A3(G138), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n467), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n482), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n487), .A2(new_n488), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n487), .A2(new_n488), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n484), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n493), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n503), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n499), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  INV_X1    g098(.A(G50), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n518), .A2(new_n520), .A3(G543), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n517), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XOR2_X1   g103(.A(new_n528), .B(KEYINPUT76), .Z(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n511), .A2(new_n513), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n521), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n531), .B(new_n532), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n521), .A2(KEYINPUT74), .A3(G543), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n525), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n540), .A2(G51), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n535), .A2(new_n541), .ZN(G168));
  AND2_X1   g117(.A1(new_n540), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n544), .A2(new_n516), .B1(new_n522), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  AND2_X1   g122(.A1(new_n540), .A2(G43), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n549), .A2(new_n516), .B1(new_n522), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT77), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT78), .Z(G188));
  NAND4_X1  g135(.A1(new_n518), .A2(new_n520), .A3(G53), .A4(G543), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n562));
  OR3_X1    g137(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT79), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n562), .B1(new_n561), .B2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n561), .A2(new_n567), .A3(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n563), .A2(new_n565), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n533), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n518), .A2(new_n520), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n533), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(G651), .A2(new_n572), .B1(new_n574), .B2(G91), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT81), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(G299));
  INV_X1    g153(.A(G171), .ZN(G301));
  INV_X1    g154(.A(G168), .ZN(G286));
  XNOR2_X1  g155(.A(G166), .B(KEYINPUT82), .ZN(G303));
  NAND2_X1  g156(.A1(new_n574), .A2(G87), .ZN(new_n582));
  INV_X1    g157(.A(new_n525), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n514), .A2(G61), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n588), .A2(new_n589), .B1(G73), .B2(G543), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n514), .A2(KEYINPUT83), .A3(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT84), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n516), .B1(new_n590), .B2(new_n591), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n574), .A2(G86), .B1(new_n583), .B2(G48), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n594), .A2(new_n597), .A3(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(new_n574), .A2(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  OAI221_X1 g177(.A(new_n600), .B1(new_n601), .B2(new_n516), .C1(new_n539), .C2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n533), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G651), .ZN(new_n608));
  INV_X1    g183(.A(G54), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n539), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g187(.A(KEYINPUT85), .B(new_n608), .C1(new_n539), .C2(new_n609), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n574), .A2(G92), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT10), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n612), .A2(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n604), .B1(G868), .B2(new_n617), .ZN(G321));
  XOR2_X1   g193(.A(G321), .B(KEYINPUT86), .Z(G284));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n576), .A2(new_n577), .ZN(new_n621));
  AOI21_X1  g196(.A(KEYINPUT81), .B1(new_n569), .B2(new_n575), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n620), .B1(G868), .B2(new_n623), .ZN(G297));
  OAI21_X1  g199(.A(new_n620), .B1(G868), .B2(new_n623), .ZN(G280));
  XNOR2_X1  g200(.A(KEYINPUT87), .B(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n617), .B1(G860), .B2(new_n626), .ZN(G148));
  INV_X1    g202(.A(new_n552), .ZN(new_n628));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n617), .A2(new_n626), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n632), .B2(new_n629), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n460), .A2(new_n464), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT12), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT13), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n479), .A2(G123), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n470), .A2(G135), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n462), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n638), .A2(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(G2427), .B(G2430), .Z(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT88), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT16), .B(G1341), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G1348), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(G14), .B1(new_n652), .B2(new_n658), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  NOR3_X1   g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(KEYINPUT17), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n664), .A2(new_n662), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n668), .B2(new_n664), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT89), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n678), .A2(new_n685), .A3(new_n681), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n684), .B(new_n686), .C1(new_n678), .C2(new_n685), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n682), .A2(new_n683), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1991), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G6), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G305), .B2(G16), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT32), .B(G1981), .Z(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(G22), .ZN(new_n703));
  MUX2_X1   g278(.A(new_n703), .B(G166), .S(G16), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(G1971), .ZN(new_n705));
  NOR2_X1   g280(.A1(G16), .A2(G23), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n586), .B2(G16), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n701), .A2(new_n702), .A3(new_n705), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT92), .Z(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n479), .A2(G119), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n470), .A2(G131), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n716), .A2(G95), .A3(G2105), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(G95), .B2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n718), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n714), .B(new_n715), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  INV_X1    g298(.A(G24), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n724), .A2(G16), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G290), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1986), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n712), .A2(new_n713), .A3(new_n723), .A4(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G19), .B(new_n628), .S(G16), .Z(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G1341), .Z(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G26), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n479), .A2(G128), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n470), .A2(G140), .ZN(new_n736));
  OR2_X1    g311(.A1(G104), .A2(G2105), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n737), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n733), .ZN(new_n741));
  MUX2_X1   g316(.A(new_n734), .B(new_n741), .S(KEYINPUT28), .Z(new_n742));
  INV_X1    g317(.A(G2067), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n617), .ZN(new_n745));
  MUX2_X1   g320(.A(G4), .B(new_n745), .S(G16), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(G1348), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(G1348), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n732), .A2(new_n744), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT94), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT26), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G105), .B2(new_n464), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n470), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n479), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G32), .B(new_n756), .S(G29), .Z(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT27), .B(G1996), .Z(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(KEYINPUT24), .A2(G34), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n733), .B1(KEYINPUT24), .B2(G34), .ZN(new_n763));
  OAI22_X1  g338(.A1(G160), .A2(new_n733), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G2084), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  NAND2_X1  g341(.A1(G171), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G5), .B2(G16), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n761), .B(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G28), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(G29), .B1(new_n770), .B2(KEYINPUT30), .ZN(new_n772));
  OR2_X1    g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  NAND2_X1  g348(.A1(KEYINPUT31), .A2(G11), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n775), .B1(new_n733), .B2(new_n643), .C1(new_n768), .C2(new_n766), .ZN(new_n776));
  INV_X1    g351(.A(G21), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G286), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n776), .B1(G1966), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n769), .B(new_n781), .C1(G1966), .C2(new_n780), .ZN(new_n782));
  NOR2_X1   g357(.A1(G29), .A2(G35), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G162), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n786), .A2(G2090), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n462), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n464), .A2(G103), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT95), .B(KEYINPUT25), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G139), .B2(new_n470), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G33), .B(new_n795), .S(G29), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT97), .B(G2072), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n764), .A2(G2084), .B1(new_n758), .B2(new_n760), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n796), .B2(new_n797), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n787), .B1(new_n802), .B2(KEYINPUT98), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(KEYINPUT98), .B2(new_n802), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n782), .B(new_n804), .C1(G2090), .C2(new_n786), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n806));
  INV_X1    g381(.A(G20), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(G16), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n806), .B(new_n808), .C1(G299), .C2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(new_n806), .B2(new_n808), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1956), .ZN(new_n811));
  NOR2_X1   g386(.A1(G27), .A2(G29), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G164), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2078), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n730), .A2(new_n750), .A3(new_n805), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  AOI22_X1  g392(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n516), .B1(new_n818), .B2(KEYINPUT100), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(KEYINPUT100), .B2(new_n818), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n536), .A2(G55), .A3(new_n538), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT101), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n574), .A2(G93), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT102), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n820), .B(KEYINPUT102), .C1(new_n824), .C2(new_n825), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n828), .A2(new_n829), .A3(new_n552), .ZN(new_n830));
  AND3_X1   g405(.A1(new_n628), .A2(new_n827), .A3(new_n826), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n617), .A2(G559), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n832), .B(new_n833), .Z(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n826), .A2(G860), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT37), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(G145));
  AOI22_X1  g416(.A1(G130), .A2(new_n479), .B1(new_n470), .B2(G142), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n844));
  INV_X1    g419(.A(G118), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n843), .A2(new_n844), .B1(new_n845), .B2(G2105), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n844), .B2(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(G162), .B(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n756), .B(new_n636), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n795), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n503), .A2(new_n506), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n739), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n720), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n472), .B(new_n643), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(G37), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n857), .B2(new_n852), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g435(.A1(new_n826), .A2(new_n629), .ZN(new_n861));
  XNOR2_X1  g436(.A(G305), .B(G288), .ZN(new_n862));
  XOR2_X1   g437(.A(G290), .B(G166), .Z(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT106), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT42), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n832), .B(new_n632), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n617), .B(new_n869), .C1(new_n621), .C2(new_n622), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(G299), .B2(new_n617), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT104), .B1(new_n623), .B2(new_n745), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(KEYINPUT105), .A3(new_n870), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n623), .A2(new_n745), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n867), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT41), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n874), .A2(new_n870), .B1(new_n623), .B2(new_n745), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n878), .B1(new_n883), .B2(new_n867), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n866), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n861), .B1(new_n885), .B2(new_n629), .ZN(G295));
  OAI21_X1  g461(.A(new_n861), .B1(new_n885), .B2(new_n629), .ZN(G331));
  INV_X1    g462(.A(new_n864), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n828), .A2(new_n829), .A3(new_n552), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n628), .A2(new_n827), .A3(new_n826), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(G301), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G301), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(new_n893), .A3(G286), .ZN(new_n894));
  OAI21_X1  g469(.A(G171), .B1(new_n830), .B2(new_n831), .ZN(new_n895));
  AOI21_X1  g470(.A(G168), .B1(new_n895), .B2(new_n891), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n877), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT107), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(G168), .A3(new_n891), .ZN(new_n899));
  OAI21_X1  g474(.A(G286), .B1(new_n892), .B2(new_n893), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n879), .A2(new_n882), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n902), .B(new_n877), .C1(new_n894), .C2(new_n896), .ZN(new_n903));
  AND4_X1   g478(.A1(new_n888), .A2(new_n898), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G37), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n899), .A3(KEYINPUT41), .ZN(new_n906));
  INV_X1    g481(.A(new_n877), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n864), .B1(new_n906), .B2(new_n880), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT109), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n898), .A2(new_n901), .A3(new_n888), .A4(new_n903), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n908), .B(new_n864), .C1(new_n880), .C2(new_n906), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n905), .A4(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(KEYINPUT43), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n898), .A2(new_n901), .A3(new_n903), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n864), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n905), .A4(new_n913), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n925), .B1(new_n923), .B2(KEYINPUT108), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n912), .A2(KEYINPUT110), .A3(KEYINPUT43), .A4(new_n916), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n919), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n913), .A2(new_n905), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n922), .B1(new_n929), .B2(new_n921), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n904), .A2(new_n911), .A3(KEYINPUT43), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(new_n925), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n933), .ZN(G397));
  XNOR2_X1  g509(.A(KEYINPUT111), .B(G1384), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n503), .B2(new_n506), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(KEYINPUT45), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n461), .A2(new_n462), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n464), .A2(G101), .ZN(new_n939));
  AND4_X1   g514(.A1(G40), .A2(new_n938), .A3(new_n471), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n941), .A2(new_n942), .A3(G1996), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n941), .B2(G1996), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n739), .B(new_n743), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n756), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n943), .B(new_n944), .C1(new_n941), .C2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n756), .B(G1996), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n720), .A2(new_n722), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n740), .A2(new_n743), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n941), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT126), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n720), .A2(new_n722), .ZN(new_n957));
  NOR4_X1   g532(.A1(new_n946), .A2(new_n950), .A3(new_n957), .A4(new_n952), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(new_n941), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n960));
  OR3_X1    g535(.A1(new_n941), .A2(G1986), .A3(G290), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n960), .B2(new_n961), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n949), .A2(new_n956), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n593), .A2(KEYINPUT84), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n598), .B1(new_n595), .B2(new_n596), .ZN(new_n966));
  OAI21_X1  g541(.A(G1981), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1981), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n594), .A2(new_n968), .A3(new_n597), .A4(new_n598), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT49), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(G1384), .B1(new_n503), .B2(new_n506), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n940), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G8), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n967), .A2(KEYINPUT49), .A3(new_n969), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n586), .A2(G1976), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(G8), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n586), .A2(G1976), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n981), .A2(KEYINPUT52), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(KEYINPUT52), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n979), .A2(KEYINPUT114), .A3(new_n983), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g563(.A1(G303), .A2(G8), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT55), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n499), .A2(new_n507), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n490), .B2(new_n498), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n940), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(G2090), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n465), .A2(G40), .A3(new_n471), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(KEYINPUT45), .B2(new_n936), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT112), .B(G1971), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n976), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n987), .A2(new_n988), .B1(new_n991), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n499), .A2(new_n507), .A3(new_n1009), .A4(new_n992), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT113), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n940), .B1(new_n973), .B2(new_n1009), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1010), .A2(KEYINPUT113), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(G2090), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n990), .B1(new_n1017), .B2(new_n976), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1008), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1004), .ZN(new_n1020));
  INV_X1    g595(.A(G2078), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT53), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n766), .B2(new_n998), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n940), .A2(KEYINPUT45), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n974), .A2(KEYINPUT115), .A3(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n499), .A2(new_n507), .A3(KEYINPUT45), .A4(new_n992), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n940), .C1(new_n973), .C2(KEYINPUT45), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1026), .A2(new_n1021), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT124), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1024), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1023), .A2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1019), .A2(G301), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1036));
  INV_X1    g611(.A(G1966), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n996), .B1(KEYINPUT50), .B2(new_n993), .ZN(new_n1039));
  INV_X1    g614(.A(G2084), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n976), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G286), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(G168), .A3(new_n1041), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G8), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n1047), .B2(new_n1045), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1043), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT62), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(new_n1043), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1035), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1007), .A2(new_n991), .ZN(new_n1056));
  INV_X1    g631(.A(new_n969), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G288), .A2(G1976), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n979), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n977), .ZN(new_n1060));
  OAI22_X1  g635(.A1(new_n1056), .A2(new_n985), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1042), .A2(G168), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1019), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n990), .A2(KEYINPUT116), .ZN(new_n1065));
  OR2_X1    g640(.A1(new_n1007), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1063), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n985), .A2(new_n1062), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1007), .A2(new_n1065), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1061), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1055), .A2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(G171), .B(KEYINPUT54), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n936), .A2(KEYINPUT45), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(KEYINPUT53), .A3(new_n1021), .A4(new_n940), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1076), .A2(new_n937), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(KEYINPUT125), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1023), .B(new_n1078), .C1(KEYINPUT125), .C2(new_n1077), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1008), .A2(new_n1018), .A3(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1080), .B(new_n1051), .C1(new_n1073), .C2(new_n1034), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n1082));
  INV_X1    g657(.A(G1956), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1001), .A2(new_n1003), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n576), .B(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1082), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1012), .B1(KEYINPUT113), .B2(new_n1010), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n508), .A2(new_n1094), .A3(new_n1009), .A4(new_n992), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1956), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1096), .A2(new_n1091), .A3(new_n1086), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT119), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1084), .A2(new_n1087), .A3(new_n1090), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1092), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1090), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1082), .B1(new_n1103), .B2(new_n1097), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT58), .B(G1341), .Z(new_n1105));
  NAND2_X1  g680(.A1(new_n974), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1004), .B2(G1996), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n552), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1107), .A2(new_n1110), .A3(new_n552), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1104), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT120), .B1(new_n1102), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1348), .B1(new_n994), .B2(new_n997), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n974), .A2(G2067), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1117), .ZN(new_n1119));
  OAI211_X1 g694(.A(KEYINPUT118), .B(new_n1119), .C1(new_n1039), .C2(G1348), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT60), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n617), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT121), .B1(new_n1126), .B2(new_n745), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n745), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1118), .A2(new_n1125), .A3(new_n1120), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1092), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(new_n1104), .A4(new_n1112), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1114), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1121), .A2(new_n745), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1099), .B1(new_n1136), .B2(new_n1103), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1081), .B1(new_n1138), .B2(KEYINPUT122), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1135), .A2(new_n1140), .A3(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1072), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(G290), .B(G1986), .Z(new_n1143));
  AOI21_X1  g718(.A(new_n941), .B1(new_n958), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n964), .B1(new_n1142), .B2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n930), .A2(new_n931), .ZN(new_n1148));
  OAI21_X1  g722(.A(G319), .B1(new_n659), .B2(new_n660), .ZN(new_n1149));
  NOR2_X1   g723(.A1(G227), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g724(.A1(new_n695), .A2(new_n859), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g725(.A(new_n1147), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1153));
  OAI211_X1 g727(.A(new_n1153), .B(KEYINPUT127), .C1(new_n930), .C2(new_n931), .ZN(new_n1154));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1154), .ZN(G308));
  NAND2_X1  g729(.A1(new_n932), .A2(new_n1153), .ZN(G225));
endmodule


