//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996, new_n997;
  XNOR2_X1  g000(.A(KEYINPUT11), .B(G169gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(G113gat), .B(G141gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT84), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT12), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n205), .A2(KEYINPUT84), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(KEYINPUT84), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT12), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT86), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NOR3_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G43gat), .B(G50gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT15), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT14), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n217), .A3(new_n218), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n223), .A2(new_n214), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n220), .A2(KEYINPUT15), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226));
  INV_X1    g025(.A(G43gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(G50gat), .ZN(new_n228));
  INV_X1    g027(.A(G50gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n229), .A2(G43gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n224), .A2(new_n225), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n213), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n221), .A2(new_n232), .A3(KEYINPUT86), .A4(KEYINPUT17), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G15gat), .B(G22gat), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT16), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G8gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n241), .B(new_n242), .C1(G1gat), .C2(new_n238), .ZN(new_n243));
  INV_X1    g042(.A(G15gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G22gat), .ZN(new_n245));
  INV_X1    g044(.A(G22gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G15gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n240), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(G1gat), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(G8gat), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n221), .A2(new_n232), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT85), .B1(new_n252), .B2(KEYINPUT17), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT85), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n233), .A2(new_n254), .A3(new_n234), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n237), .A2(new_n251), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n243), .A2(new_n250), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(new_n233), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n256), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT90), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n260), .A2(KEYINPUT90), .A3(new_n261), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n212), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n256), .A2(KEYINPUT18), .A3(new_n257), .A4(new_n259), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT87), .B1(new_n258), .B2(new_n233), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n259), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n257), .B(KEYINPUT13), .Z(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT88), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT88), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n271), .A2(new_n275), .A3(new_n272), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n266), .A2(new_n267), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n267), .A2(new_n274), .A3(new_n276), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT89), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT89), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n267), .A2(new_n274), .A3(new_n281), .A4(new_n276), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n282), .A3(new_n262), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n212), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G230gat), .A2(G233gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT97), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G57gat), .B(G64gat), .Z(new_n289));
  OR2_X1    g088(.A1(G71gat), .A2(G78gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G71gat), .A2(G78gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT9), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n289), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G57gat), .B(G64gat), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n291), .B(new_n290), .C1(new_n296), .C2(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G99gat), .A2(G106gat), .ZN(new_n299));
  INV_X1    g098(.A(G85gat), .ZN(new_n300));
  INV_X1    g099(.A(G92gat), .ZN(new_n301));
  AOI22_X1  g100(.A1(KEYINPUT8), .A2(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G85gat), .A2(G92gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT95), .ZN(new_n308));
  XOR2_X1   g107(.A(G99gat), .B(G106gat), .Z(new_n309));
  AND2_X1   g108(.A1(new_n305), .A2(new_n306), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT95), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(new_n302), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n309), .B1(new_n308), .B2(new_n312), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n298), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n309), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n307), .A2(KEYINPUT95), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n311), .B1(new_n310), .B2(new_n302), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n295), .A2(new_n297), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT10), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n321), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(KEYINPUT10), .A3(new_n320), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n288), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G120gat), .B(G148gat), .ZN(new_n328));
  INV_X1    g127(.A(G176gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G204gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n322), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n327), .B(new_n333), .C1(new_n334), .C2(new_n288), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT10), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n313), .A2(new_n314), .A3(new_n298), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n287), .B1(new_n339), .B2(new_n325), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n334), .A2(new_n288), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n332), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n335), .A2(new_n342), .A3(KEYINPUT98), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT98), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n344), .B(new_n332), .C1(new_n340), .C2(new_n341), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n285), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  OR2_X1    g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(KEYINPUT2), .ZN(new_n351));
  XNOR2_X1  g150(.A(G141gat), .B(G148gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(KEYINPUT76), .ZN(new_n353));
  INV_X1    g152(.A(G148gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G141gat), .ZN(new_n355));
  INV_X1    g154(.A(G141gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G148gat), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT76), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n351), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n349), .B(new_n350), .C1(new_n352), .C2(KEYINPUT2), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(G197gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n331), .ZN(new_n364));
  NAND2_X1  g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365));
  OR2_X1    g164(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(G218gat), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT22), .ZN(new_n369));
  AOI221_X4 g168(.A(G211gat), .B1(new_n364), .B2(new_n365), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G211gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n369), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n364), .A2(new_n365), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n362), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  AND2_X1   g174(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT22), .B1(new_n378), .B2(G218gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n373), .ZN(new_n380));
  OAI21_X1  g179(.A(G211gat), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n372), .A2(new_n371), .A3(new_n373), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(G218gat), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n375), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n361), .B1(new_n384), .B2(KEYINPUT3), .ZN(new_n385));
  INV_X1    g184(.A(G228gat), .ZN(new_n386));
  INV_X1    g185(.A(G233gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(new_n383), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n359), .A2(new_n391), .A3(new_n360), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n385), .A2(new_n388), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n361), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n393), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n402));
  OAI22_X1  g201(.A1(new_n401), .A2(new_n402), .B1(new_n386), .B2(new_n387), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n385), .A2(new_n395), .A3(KEYINPUT80), .A4(new_n388), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n406), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n398), .A2(new_n403), .A3(new_n408), .A4(new_n404), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT31), .B(G50gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT79), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G22gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n407), .A2(new_n413), .A3(new_n409), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT0), .B(G57gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G85gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(G134gat), .ZN(new_n424));
  INV_X1    g223(.A(G120gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(G113gat), .ZN(new_n426));
  INV_X1    g225(.A(G113gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G120gat), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT1), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G127gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT1), .B(G127gat), .C1(new_n426), .C2(new_n428), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n424), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n430), .ZN(new_n434));
  XNOR2_X1  g233(.A(G113gat), .B(G120gat), .ZN(new_n435));
  OAI21_X1  g234(.A(G127gat), .B1(new_n435), .B2(KEYINPUT1), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n436), .A3(G134gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n361), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n433), .A2(new_n437), .A3(new_n359), .A4(new_n360), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n423), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT5), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT78), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n423), .ZN(new_n444));
  INV_X1    g243(.A(new_n440), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n433), .A2(new_n437), .B1(new_n359), .B2(new_n360), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(KEYINPUT4), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n361), .A2(KEYINPUT3), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(new_n438), .A3(new_n392), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n444), .B1(new_n440), .B2(new_n455), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n443), .A2(new_n449), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n452), .B(new_n459), .C1(new_n440), .C2(new_n455), .ZN(new_n460));
  NOR3_X1   g259(.A1(new_n460), .A2(KEYINPUT5), .A3(new_n444), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n422), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n444), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n439), .A2(new_n440), .A3(new_n423), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT39), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(KEYINPUT81), .A3(KEYINPUT39), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n460), .A2(new_n470), .A3(new_n444), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(KEYINPUT40), .A3(new_n421), .A4(new_n471), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n462), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G183gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT69), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(G183gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT27), .ZN(new_n478));
  NOR2_X1   g277(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n482));
  INV_X1    g281(.A(G190gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n474), .A2(new_n483), .ZN(new_n485));
  AND2_X1   g284(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n483), .B1(new_n486), .B2(new_n479), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n485), .B1(new_n487), .B2(KEYINPUT28), .ZN(new_n488));
  INV_X1    g287(.A(G169gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n329), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n490), .A2(KEYINPUT26), .ZN(new_n491));
  NAND2_X1  g290(.A1(G169gat), .A2(G176gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT67), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(G169gat), .A3(G176gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n490), .A2(KEYINPUT26), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n484), .A2(new_n488), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT23), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n490), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT65), .B(G176gat), .Z(new_n503));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT23), .A4(new_n489), .ZN(new_n505));
  AND3_X1   g304(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n474), .A2(new_n483), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT25), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(KEYINPUT65), .B(G176gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n489), .A2(KEYINPUT23), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT66), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n502), .A2(new_n505), .A3(new_n510), .A4(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n496), .B(new_n501), .C1(G176gat), .C2(new_n512), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n516));
  AOI21_X1  g315(.A(G190gat), .B1(new_n475), .B2(new_n477), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n506), .ZN(new_n518));
  INV_X1    g317(.A(new_n507), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n506), .B2(new_n516), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n515), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT25), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n499), .B(new_n514), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n525), .B1(new_n524), .B2(new_n393), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(new_n390), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n525), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n389), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G8gat), .B(G36gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(G64gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(new_n301), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(KEYINPUT30), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n536), .B(KEYINPUT75), .Z(new_n540));
  OAI211_X1 g339(.A(new_n538), .B(KEYINPUT30), .C1(new_n533), .C2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n469), .A2(new_n421), .A3(new_n471), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT40), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n473), .A2(new_n539), .A3(new_n541), .A4(new_n544), .ZN(new_n545));
  OR3_X1    g344(.A1(new_n526), .A2(new_n531), .A3(new_n389), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n546), .B(KEYINPUT37), .C1(new_n390), .C2(new_n528), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT82), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT37), .B1(new_n529), .B2(new_n532), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n551), .A2(KEYINPUT38), .A3(new_n540), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n529), .A2(KEYINPUT37), .A3(new_n532), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n536), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT38), .B1(new_n555), .B2(new_n551), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n450), .A2(new_n452), .A3(new_n456), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n448), .B1(new_n447), .B2(KEYINPUT5), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n441), .A2(KEYINPUT78), .A3(new_n442), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n461), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n421), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n462), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(KEYINPUT6), .B(new_n422), .C1(new_n457), .C2(new_n461), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n556), .A2(new_n564), .A3(new_n565), .A4(new_n538), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n417), .B(new_n545), .C1(new_n553), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n539), .A2(new_n541), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n570), .A2(new_n416), .A3(new_n415), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT70), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n524), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n506), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT69), .B(G183gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(G190gat), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n520), .B1(new_n576), .B2(new_n516), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT25), .B1(new_n577), .B2(new_n515), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n578), .A2(KEYINPUT70), .A3(new_n499), .A4(new_n514), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n438), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G227gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT64), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n524), .A2(new_n572), .A3(new_n437), .A4(new_n433), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT32), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G15gat), .B(G43gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(G71gat), .B(G99gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n585), .B(KEYINPUT32), .C1(new_n587), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n580), .A2(new_n584), .B1(G227gat), .B2(G233gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT71), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT34), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n584), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n582), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n600), .B(new_n601), .C1(KEYINPUT71), .C2(new_n596), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n601), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT71), .B1(new_n599), .B2(new_n581), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n598), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n594), .A3(new_n592), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT36), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT72), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n595), .A2(KEYINPUT72), .A3(new_n598), .A4(new_n602), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(KEYINPUT36), .A3(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n567), .A2(new_n571), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n611), .A2(new_n612), .B1(new_n416), .B2(new_n415), .ZN(new_n616));
  INV_X1    g415(.A(new_n570), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n608), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n417), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n568), .A2(new_n569), .A3(new_n615), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n614), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT83), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n614), .B(KEYINPUT83), .C1(new_n618), .C2(new_n622), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n348), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n298), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G183gat), .B(G211gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT94), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n632), .B(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT19), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n320), .A2(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n251), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT93), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT92), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT93), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n639), .B(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT92), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n637), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G231gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n387), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(KEYINPUT92), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n640), .A2(new_n641), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT19), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n646), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n649), .B1(new_n646), .B2(new_n652), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n636), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n652), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT19), .B1(new_n650), .B2(new_n651), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n646), .A2(new_n649), .A3(new_n652), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n659), .A3(new_n635), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT96), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n313), .A2(new_n314), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n237), .A2(new_n664), .A3(new_n253), .A4(new_n255), .ZN(new_n665));
  AND3_X1   g464(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n324), .B2(new_n233), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n483), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n483), .A3(new_n667), .ZN(new_n670));
  AOI21_X1  g469(.A(G218gat), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n672), .A2(new_n362), .A3(new_n668), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n663), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n362), .B1(new_n672), .B2(new_n668), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n669), .A2(G218gat), .A3(new_n670), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT96), .ZN(new_n677));
  XNOR2_X1  g476(.A(G134gat), .B(G162gat), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n674), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n677), .A2(new_n681), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n662), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n627), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n569), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g488(.A1(new_n539), .A2(new_n541), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n627), .A2(new_n685), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G8gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT99), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT16), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n242), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n242), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n686), .A2(new_n690), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(KEYINPUT42), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n693), .B1(new_n699), .B2(new_n700), .ZN(G1325gat));
  AOI21_X1  g500(.A(G15gat), .B1(new_n686), .B2(new_n619), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n609), .A2(new_n613), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n686), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(G15gat), .B2(new_n704), .ZN(G1326gat));
  INV_X1    g504(.A(new_n417), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n686), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT43), .B(G22gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  AND3_X1   g508(.A1(new_n627), .A2(new_n662), .A3(new_n684), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n217), .A3(new_n687), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(KEYINPUT45), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT44), .B1(new_n623), .B2(new_n684), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n625), .A2(new_n626), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n661), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n655), .A2(KEYINPUT100), .A3(new_n660), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(new_n348), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n717), .A2(new_n687), .A3(new_n722), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n712), .A2(new_n713), .B1(new_n217), .B2(new_n723), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n710), .A2(new_n218), .A3(new_n690), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT101), .B(KEYINPUT46), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n717), .A2(new_n690), .A3(new_n722), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G36gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(G1329gat));
  NAND3_X1  g530(.A1(new_n710), .A2(new_n227), .A3(new_n619), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n716), .ZN(new_n733));
  INV_X1    g532(.A(new_n714), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n733), .A2(new_n703), .A3(new_n734), .A4(new_n722), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(G43gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n732), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n732), .B2(new_n736), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(G1330gat));
  INV_X1    g539(.A(KEYINPUT102), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n627), .A2(new_n662), .A3(new_n684), .A4(new_n706), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n229), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n717), .A2(G50gat), .A3(new_n706), .A4(new_n722), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n741), .B(KEYINPUT48), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(KEYINPUT48), .ZN(new_n747));
  AND4_X1   g546(.A1(new_n746), .A2(new_n743), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n745), .A2(new_n748), .ZN(G1331gat));
  NOR4_X1   g548(.A1(new_n662), .A2(new_n684), .A3(new_n285), .A4(new_n347), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n623), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n569), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(G57gat), .Z(G1332gat));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n751), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n690), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  OAI21_X1  g557(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(G1333gat));
  NOR3_X1   g558(.A1(new_n751), .A2(G71gat), .A3(new_n608), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n703), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(G71gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n755), .A2(new_n706), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT104), .B(G78gat), .Z(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n661), .A2(new_n285), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n769), .A2(KEYINPUT106), .A3(new_n346), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT106), .B1(new_n769), .B2(new_n346), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n717), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n569), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n623), .A2(new_n684), .A3(new_n769), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n775), .A2(KEYINPUT108), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n623), .A2(KEYINPUT51), .A3(new_n684), .A4(new_n769), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n300), .A3(new_n687), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n774), .B1(new_n788), .B2(new_n347), .ZN(G1336gat));
  NAND4_X1  g588(.A1(new_n733), .A2(new_n690), .A3(new_n734), .A4(new_n772), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G92gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT111), .B1(new_n775), .B2(new_n776), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n775), .A2(KEYINPUT111), .A3(new_n776), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n783), .A2(KEYINPUT107), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n783), .A2(KEYINPUT107), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n568), .A2(new_n347), .A3(G92gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT110), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n791), .A2(new_n792), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n790), .A2(KEYINPUT109), .A3(G92gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n781), .B2(new_n785), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n791), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n800), .A2(new_n801), .B1(new_n803), .B2(new_n804), .ZN(G1337gat));
  NOR3_X1   g604(.A1(new_n608), .A2(G99gat), .A3(new_n347), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT112), .Z(new_n807));
  NAND2_X1  g606(.A1(new_n787), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n703), .ZN(new_n809));
  OAI21_X1  g608(.A(G99gat), .B1(new_n773), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1338gat));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n417), .A2(G106gat), .A3(new_n347), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT113), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n717), .A2(new_n706), .A3(new_n772), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n797), .A2(new_n815), .B1(new_n816), .B2(G106gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(G106gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n812), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n814), .B1(new_n782), .B2(new_n786), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n812), .A2(new_n817), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  AOI21_X1  g620(.A(new_n257), .B1(new_n256), .B2(new_n259), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n271), .A2(new_n272), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n205), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n824), .B(KEYINPUT115), .Z(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n278), .A3(new_n346), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n333), .B1(new_n340), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n339), .A2(new_n325), .A3(new_n287), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n327), .A2(new_n829), .A3(KEYINPUT54), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n212), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n279), .A2(KEYINPUT89), .B1(new_n261), .B2(new_n260), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n834), .B1(new_n835), .B2(new_n282), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n212), .B(new_n279), .C1(new_n264), .C2(new_n265), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n830), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n839), .A2(new_n840), .A3(new_n335), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n839), .B2(new_n335), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n826), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n682), .A2(new_n683), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n825), .A2(new_n278), .A3(new_n833), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n839), .A2(new_n335), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n839), .A2(new_n840), .A3(new_n335), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n684), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n721), .B1(new_n846), .B2(new_n853), .ZN(new_n854));
  NOR4_X1   g653(.A1(new_n662), .A2(new_n684), .A3(new_n285), .A4(new_n346), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n616), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n690), .A2(new_n569), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n427), .A3(new_n285), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n719), .A2(new_n720), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n852), .A2(new_n285), .A3(new_n833), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n684), .B1(new_n863), .B2(new_n826), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n845), .A2(new_n847), .A3(new_n843), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n285), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n685), .A2(new_n867), .A3(new_n347), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n620), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n858), .ZN(new_n870));
  OAI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n861), .A2(new_n871), .ZN(G1340gat));
  NAND3_X1  g671(.A1(new_n860), .A2(new_n425), .A3(new_n346), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n869), .A2(new_n346), .A3(new_n858), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT116), .B1(new_n874), .B2(G120gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT117), .Z(G1341gat));
  AOI21_X1  g677(.A(G127gat), .B1(new_n860), .B2(new_n661), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n870), .A2(new_n430), .A3(new_n862), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(G1342gat));
  NAND3_X1  g680(.A1(new_n860), .A2(new_n424), .A3(new_n684), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n885));
  OAI21_X1  g684(.A(G134gat), .B1(new_n870), .B2(new_n845), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(KEYINPUT118), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(G1343gat));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n868), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n706), .A3(new_n809), .ZN(new_n890));
  NOR4_X1   g689(.A1(new_n890), .A2(G141gat), .A3(new_n867), .A4(new_n859), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(KEYINPUT58), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n703), .A2(new_n859), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n285), .A2(new_n335), .A3(new_n833), .A4(new_n839), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n684), .B1(new_n894), .B2(new_n826), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n662), .B1(new_n895), .B2(new_n865), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n417), .B1(new_n896), .B2(new_n868), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n856), .A2(KEYINPUT57), .A3(new_n417), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n899), .A2(new_n900), .A3(new_n867), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n892), .B1(new_n356), .B2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT119), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  INV_X1    g703(.A(new_n893), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n826), .B1(new_n838), .B2(new_n849), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n845), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n661), .B1(new_n907), .B2(new_n853), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n706), .B1(new_n908), .B2(new_n855), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n905), .B1(new_n909), .B2(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n889), .A2(new_n898), .A3(new_n706), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n285), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n891), .B1(new_n913), .B2(G141gat), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n902), .B1(new_n914), .B2(new_n915), .ZN(G1344gat));
  OAI21_X1  g715(.A(KEYINPUT119), .B1(new_n899), .B2(new_n900), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n910), .A2(new_n904), .A3(new_n911), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n347), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT120), .B1(new_n897), .B2(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT120), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n909), .A2(new_n921), .A3(new_n898), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n889), .A2(KEYINPUT57), .A3(new_n706), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(new_n346), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n893), .A2(KEYINPUT59), .ZN(new_n926));
  OAI22_X1  g725(.A1(new_n919), .A2(KEYINPUT59), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n890), .A2(new_n859), .ZN(new_n928));
  AOI21_X1  g727(.A(G148gat), .B1(new_n928), .B2(new_n346), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n927), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n929), .ZN(G1345gat));
  AOI21_X1  g729(.A(G155gat), .B1(new_n928), .B2(new_n661), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n862), .B1(new_n917), .B2(new_n918), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g732(.A(G162gat), .B1(new_n928), .B2(new_n684), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n845), .B1(new_n917), .B2(new_n918), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n935), .B2(G162gat), .ZN(G1347gat));
  INV_X1    g735(.A(new_n620), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n690), .A2(new_n569), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT121), .Z(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n939), .C1(new_n854), .C2(new_n855), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n867), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n856), .A2(new_n857), .ZN(new_n942));
  INV_X1    g741(.A(new_n938), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n489), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n941), .B1(new_n944), .B2(new_n867), .ZN(G1348gat));
  NOR3_X1   g744(.A1(new_n940), .A2(new_n503), .A3(new_n347), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n946), .A2(KEYINPUT122), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n946), .A2(KEYINPUT122), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n346), .A3(new_n943), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n947), .B(new_n948), .C1(new_n329), .C2(new_n949), .ZN(G1349gat));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT123), .B1(new_n940), .B2(new_n862), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n869), .A2(new_n953), .A3(new_n721), .A4(new_n939), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n954), .A3(new_n575), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n486), .A2(new_n479), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n661), .A3(new_n957), .A4(new_n943), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n955), .B2(new_n958), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n955), .A2(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(KEYINPUT60), .A3(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n961), .A2(new_n965), .ZN(G1350gat));
  OAI21_X1  g765(.A(G190gat), .B1(new_n940), .B2(new_n845), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n942), .A2(new_n483), .A3(new_n684), .A4(new_n943), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n968), .B2(new_n969), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n939), .A2(new_n809), .ZN(new_n975));
  XOR2_X1   g774(.A(new_n975), .B(KEYINPUT127), .Z(new_n976));
  NAND2_X1  g775(.A1(new_n924), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n867), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n890), .A2(new_n687), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n690), .ZN(new_n981));
  NOR4_X1   g780(.A1(new_n890), .A2(KEYINPUT126), .A3(new_n687), .A4(new_n568), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n363), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n978), .B1(new_n983), .B2(new_n867), .ZN(G1352gat));
  NOR2_X1   g783(.A1(new_n347), .A2(G204gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n980), .A2(new_n690), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT62), .Z(new_n987));
  AND3_X1   g786(.A1(new_n924), .A2(new_n346), .A3(new_n976), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n987), .B1(new_n331), .B2(new_n988), .ZN(G1353gat));
  OAI221_X1 g788(.A(new_n661), .B1(new_n377), .B2(new_n376), .C1(new_n981), .C2(new_n982), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n924), .A2(new_n661), .A3(new_n976), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n991), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT63), .B1(new_n991), .B2(G211gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  OAI21_X1  g793(.A(G218gat), .B1(new_n977), .B2(new_n845), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n981), .A2(new_n982), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n684), .A2(new_n362), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(G1355gat));
endmodule


