//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(KEYINPUT66), .B1(G567), .B2(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XOR2_X1   g035(.A(KEYINPUT67), .B(G2105), .Z(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n462), .A2(G137), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT67), .B(G2105), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OR3_X1    g048(.A1(new_n467), .A2(KEYINPUT69), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT69), .B1(new_n467), .B2(new_n473), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(G160));
  OAI221_X1 g051(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n461), .C2(G112), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n462), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT70), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n462), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n477), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n462), .A2(new_n472), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT71), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n462), .A2(new_n472), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n486), .B1(G124), .B2(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .ZN(new_n496));
  INV_X1    g071(.A(G126), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(new_n478), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n498), .B2(new_n462), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n462), .B(KEYINPUT68), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n461), .A2(G138), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n506), .A2(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n518), .A2(new_n521), .ZN(G166));
  XOR2_X1   g097(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n507), .A2(new_n508), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n512), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n526), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n525), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n535), .B1(new_n529), .B2(new_n530), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n513), .A2(KEYINPUT72), .A3(new_n514), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n538), .A2(G63), .A3(G651), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n534), .A2(new_n539), .ZN(G168));
  NAND2_X1  g115(.A1(new_n538), .A2(G64), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n520), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n544), .A2(new_n510), .B1(new_n516), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n548), .A2(new_n510), .B1(new_n516), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n536), .A2(new_n537), .A3(G56), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n520), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n552), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI211_X1 g139(.A(KEYINPUT75), .B(new_n563), .C1(new_n510), .C2(new_n564), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n515), .A2(G65), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  XOR2_X1   g142(.A(new_n567), .B(KEYINPUT76), .Z(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n532), .A2(G91), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n565), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT75), .B1(new_n510), .B2(new_n564), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n527), .A2(new_n573), .A3(G53), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G168), .ZN(G286));
  INV_X1    g153(.A(G166), .ZN(G303));
  AOI22_X1  g154(.A1(G87), .A2(new_n532), .B1(new_n527), .B2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n581), .A2(KEYINPUT77), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n581), .A2(KEYINPUT77), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n515), .A2(G61), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(KEYINPUT78), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n585), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n520), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  INV_X1    g164(.A(G86), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n589), .A2(new_n510), .B1(new_n516), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n520), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n532), .A2(G85), .ZN(new_n596));
  XOR2_X1   g171(.A(KEYINPUT79), .B(G47), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n527), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT80), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n598), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n595), .B1(new_n599), .B2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n532), .A2(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G79), .ZN(new_n608));
  OR3_X1    g183(.A1(new_n608), .A2(new_n512), .A3(KEYINPUT81), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT81), .B1(new_n608), .B2(new_n512), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n531), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n604), .B1(G868), .B2(new_n615), .ZN(G284));
  OAI21_X1  g191(.A(new_n604), .B1(G868), .B2(new_n615), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n622), .B2(G860), .ZN(G148));
  NOR2_X1   g198(.A1(new_n557), .A2(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n615), .A2(new_n622), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n464), .A2(new_n469), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n491), .A2(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n461), .C2(G111), .ZN(new_n636));
  INV_X1    g211(.A(G135), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n484), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND3_X1  g214(.A1(new_n633), .A2(new_n634), .A3(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n643), .A2(new_n646), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n641), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n655), .ZN(new_n657));
  INV_X1    g232(.A(new_n641), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(new_n653), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n662), .B1(new_n656), .B2(new_n659), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n667));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n672), .B1(new_n670), .B2(new_n668), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(new_n669), .B2(new_n670), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(new_n670), .A3(new_n668), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  NOR3_X1   g252(.A1(new_n673), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  OR3_X1    g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n682), .A2(new_n685), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n682), .A2(new_n686), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n687), .A2(new_n690), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT88), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n694), .B(new_n696), .ZN(new_n706));
  INV_X1    g281(.A(new_n699), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n703), .B1(new_n700), .B2(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(G229));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G27), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(G164), .B2(new_n712), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2078), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NOR2_X1   g291(.A1(G168), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n716), .B2(G21), .ZN(new_n718));
  INV_X1    g293(.A(G1966), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT31), .B(G11), .ZN(new_n722));
  INV_X1    g297(.A(G28), .ZN(new_n723));
  AOI21_X1  g298(.A(G29), .B1(new_n723), .B2(KEYINPUT30), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT100), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT99), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n727), .A2(new_n723), .A3(KEYINPUT30), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n723), .B2(KEYINPUT30), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(new_n725), .C2(KEYINPUT100), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n722), .B1(new_n726), .B2(new_n730), .C1(new_n638), .C2(new_n712), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n720), .A2(new_n721), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT93), .B(G2067), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n712), .A2(G26), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT28), .Z(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n736));
  INV_X1    g311(.A(G116), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n472), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n483), .B2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n491), .A2(G128), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(G29), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n715), .B(new_n732), .C1(new_n733), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n712), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n712), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT29), .Z(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(KEYINPUT101), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(KEYINPUT101), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n716), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n619), .B2(new_n716), .ZN(new_n753));
  INV_X1    g328(.A(G1956), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n743), .A2(new_n749), .A3(new_n750), .A4(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n469), .A2(KEYINPUT96), .A3(G105), .ZN(new_n760));
  AOI21_X1  g335(.A(KEYINPUT96), .B1(new_n469), .B2(G105), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n491), .B2(G129), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n483), .A2(G141), .ZN(new_n765));
  AND3_X1   g340(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n769), .B(KEYINPUT98), .C1(G29), .C2(G32), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT98), .B2(new_n769), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT27), .B(G1996), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n746), .A2(new_n747), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n775), .B2(KEYINPUT24), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT95), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n775), .A2(KEYINPUT24), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n776), .B2(KEYINPUT95), .ZN(new_n779));
  AOI22_X1  g354(.A1(G160), .A2(G29), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n774), .B1(G2084), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n712), .A2(G33), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT25), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n483), .A2(G139), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n464), .A2(G127), .ZN(new_n786));
  NAND2_X1  g361(.A1(G115), .A2(G2104), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n461), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n784), .B(new_n785), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n782), .B1(new_n792), .B2(new_n712), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n716), .A2(G19), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n557), .B2(new_n716), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n793), .A2(G2072), .B1(G1341), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n780), .A2(G2084), .ZN(new_n797));
  NOR2_X1   g372(.A1(G4), .A2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT92), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n614), .B2(new_n716), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n733), .B2(new_n742), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n793), .A2(G2072), .B1(G1341), .B2(new_n795), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n716), .A2(G5), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G171), .B2(new_n716), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1961), .ZN(new_n806));
  NOR4_X1   g381(.A1(new_n797), .A2(new_n802), .A3(new_n803), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n781), .A2(new_n796), .A3(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n756), .A2(new_n773), .A3(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G23), .B(G288), .S(G16), .Z(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT33), .B(G1976), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n592), .A2(G16), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G6), .B2(G16), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT32), .B(G1981), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n815), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n716), .A2(G22), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n716), .ZN(new_n821));
  INV_X1    g396(.A(G1971), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n813), .A2(new_n818), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT91), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT34), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(G290), .A2(G16), .ZN(new_n828));
  INV_X1    g403(.A(G24), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n829), .A2(KEYINPUT90), .A3(G16), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT90), .B1(new_n829), .B2(G16), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(G1986), .Z(new_n833));
  OR2_X1    g408(.A1(G25), .A2(G29), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(G107), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n835), .B1(new_n472), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n491), .B2(G119), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n483), .A2(KEYINPUT89), .A3(G131), .ZN(new_n839));
  AOI21_X1  g414(.A(KEYINPUT89), .B1(new_n483), .B2(G131), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n834), .B1(new_n841), .B2(new_n712), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n833), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(new_n825), .B2(new_n826), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n827), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT36), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT36), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n827), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n810), .B1(new_n849), .B2(new_n851), .ZN(G311));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n809), .ZN(G150));
  NAND3_X1  g429(.A1(new_n536), .A2(new_n537), .A3(G67), .ZN(new_n855));
  INV_X1    g430(.A(G80), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(new_n512), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G651), .ZN(new_n858));
  AOI22_X1  g433(.A1(G93), .A2(new_n532), .B1(new_n527), .B2(G55), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n553), .A2(new_n554), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(G651), .A3(new_n556), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  INV_X1    g440(.A(new_n550), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n864), .A2(new_n866), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(KEYINPUT102), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n557), .A2(new_n865), .A3(KEYINPUT103), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT103), .B1(new_n557), .B2(new_n865), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n860), .B1(new_n557), .B2(new_n865), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n552), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT74), .B1(new_n551), .B2(new_n552), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n877), .A2(new_n878), .A3(new_n520), .ZN(new_n879));
  OAI211_X1 g454(.A(KEYINPUT102), .B(new_n870), .C1(new_n879), .C2(new_n550), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n614), .A2(new_n622), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  XNOR2_X1  g460(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(G860), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n862), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n895), .B(KEYINPUT105), .Z(G145));
  INV_X1    g471(.A(new_n792), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n504), .B1(new_n766), .B2(new_n767), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n763), .A2(new_n765), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT97), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(G164), .A3(new_n901), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n898), .A2(new_n902), .A3(new_n741), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n741), .B1(new_n898), .B2(new_n902), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n897), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n741), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n766), .A2(new_n767), .A3(new_n504), .ZN(new_n907));
  AOI21_X1  g482(.A(G164), .B1(new_n900), .B2(new_n901), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n898), .A2(new_n902), .A3(new_n741), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n792), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n841), .B(new_n630), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n483), .A2(G142), .ZN(new_n914));
  OAI21_X1  g489(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n915));
  INV_X1    g490(.A(G118), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n472), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G130), .ZN(new_n919));
  INV_X1    g494(.A(new_n491), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n913), .B(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G162), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n474), .A2(new_n475), .ZN(new_n925));
  INV_X1    g500(.A(new_n638), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n925), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n927), .A3(G162), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n921), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n913), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n913), .A2(new_n934), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n911), .A3(new_n905), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n923), .A2(new_n933), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT106), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n912), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n922), .A2(new_n905), .A3(KEYINPUT106), .A4(new_n911), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n930), .A2(new_n932), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G37), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n939), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n948));
  NAND2_X1  g523(.A1(G299), .A2(new_n614), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n571), .A2(new_n607), .A3(new_n575), .A4(new_n613), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n948), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n949), .A2(new_n953), .A3(new_n950), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n949), .B2(new_n950), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n954), .B1(new_n957), .B2(new_n948), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n882), .B(new_n625), .ZN(new_n959));
  MUX2_X1   g534(.A(new_n958), .B(new_n952), .S(new_n959), .Z(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n602), .A2(new_n599), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n581), .B(KEYINPUT77), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n962), .A2(new_n963), .A3(new_n580), .A4(new_n595), .ZN(new_n964));
  NAND2_X1  g539(.A1(G290), .A2(G288), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n592), .B(G166), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n965), .A3(new_n961), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n967), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n971), .B2(new_n966), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n960), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n960), .A2(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(G868), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G868), .B2(new_n868), .ZN(G295));
  OAI21_X1  g552(.A(new_n976), .B1(G868), .B2(new_n868), .ZN(G331));
  NAND2_X1  g553(.A1(new_n972), .A2(KEYINPUT112), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n969), .B(new_n980), .C1(new_n971), .C2(new_n966), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(G171), .B(G168), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n875), .A2(new_n876), .A3(new_n880), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n875), .A2(new_n880), .B1(new_n868), .B2(new_n867), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(G171), .B(G168), .Z(new_n987));
  NAND3_X1  g562(.A1(new_n874), .A2(new_n881), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(KEYINPUT110), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n874), .A2(new_n987), .A3(new_n990), .A4(new_n881), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n989), .A2(new_n958), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n986), .A2(KEYINPUT111), .A3(new_n988), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n882), .A2(new_n994), .A3(new_n983), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n951), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n982), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n995), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n952), .ZN(new_n999));
  INV_X1    g574(.A(new_n972), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n989), .A2(new_n958), .A3(new_n991), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(new_n1002), .A3(new_n945), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n998), .A2(new_n957), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n951), .B1(new_n989), .B2(new_n991), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n982), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n945), .A4(new_n1002), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1002), .A2(new_n945), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(new_n1007), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT44), .B1(new_n1014), .B2(new_n1008), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(G397));
  INV_X1    g592(.A(G40), .ZN(new_n1018));
  OR3_X1    g593(.A1(new_n467), .A2(new_n1018), .A3(new_n473), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT113), .B(G1384), .ZN(new_n1020));
  AND2_X1   g595(.A1(new_n504), .A2(new_n1020), .ZN(new_n1021));
  OR3_X1    g596(.A1(new_n1019), .A2(new_n1021), .A3(KEYINPUT45), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT114), .ZN(new_n1023));
  INV_X1    g598(.A(G2067), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n741), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1996), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(new_n768), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1022), .A2(G1996), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1023), .A2(new_n1027), .B1(new_n768), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1023), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n841), .B(new_n843), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1022), .ZN(new_n1033));
  XNOR2_X1  g608(.A(G290), .B(G1986), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n504), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n467), .A2(new_n1018), .A3(new_n473), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n499), .B2(new_n503), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1961), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1021), .A2(KEYINPUT45), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G2078), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n504), .A2(KEYINPUT45), .A3(new_n1020), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1047), .A2(new_n1040), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1038), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G2078), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1040), .A4(new_n1050), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n1048), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1055), .B2(new_n1048), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1046), .B(new_n1051), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1036), .B1(new_n1060), .B2(G171), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(new_n1048), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT122), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1064), .A2(new_n1057), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1041), .A2(KEYINPUT45), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(new_n1019), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1067), .B(new_n1049), .C1(new_n1052), .C2(new_n1038), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(G301), .A3(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1061), .A2(new_n1062), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1062), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT56), .B(G2072), .Z(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1067), .A2(new_n1073), .A3(new_n1050), .A4(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1050), .B(new_n1040), .C1(KEYINPUT45), .C2(new_n1041), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n1077), .B2(new_n1074), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1044), .A2(new_n754), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1081), .A2(KEYINPUT57), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(KEYINPUT57), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n619), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(G299), .A2(new_n1081), .A3(KEYINPUT57), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1044), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1040), .A2(new_n1024), .A3(new_n1041), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n614), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1086), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1076), .A2(new_n1078), .A3(new_n1092), .A4(new_n1079), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1087), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1089), .A2(new_n1090), .A3(new_n614), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT60), .B1(new_n1095), .B2(new_n1091), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT58), .B(G1341), .Z(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1019), .B2(new_n1038), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT120), .B(G1996), .Z(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1077), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n557), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1103), .A3(new_n557), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n614), .A2(KEYINPUT60), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1089), .A2(new_n1090), .A3(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1096), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1093), .B(KEYINPUT61), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1094), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(G301), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1060), .A2(G171), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1036), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1040), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1038), .A2(new_n1052), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n719), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G2084), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1039), .A2(new_n1118), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G8), .ZN(new_n1121));
  NOR2_X1   g696(.A1(G168), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT121), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1114), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1121), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n1125), .A2(KEYINPUT51), .A3(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G303), .A2(G8), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT55), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1044), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT115), .B(G2090), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1131), .A2(new_n1132), .B1(new_n1077), .B2(new_n822), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1130), .B1(new_n1133), .B2(new_n1121), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1121), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n1136), .B2(G288), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT52), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT49), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT116), .B(G1981), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n588), .A2(new_n591), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(G1981), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n592), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1139), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1141), .B(KEYINPUT49), .C1(new_n1143), .C2(new_n592), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1145), .A2(new_n1135), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1135), .B(new_n1148), .C1(new_n1136), .C2(G288), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1138), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1130), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1077), .A2(new_n822), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1132), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1044), .A2(new_n1154), .ZN(new_n1155));
  OAI211_X1 g730(.A(G8), .B(new_n1152), .C1(new_n1153), .C2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1134), .A2(new_n1151), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1128), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1110), .A2(new_n1113), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1072), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT124), .B1(new_n1128), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1157), .B1(new_n1128), .B2(new_n1161), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1126), .A2(new_n1127), .A3(new_n1164), .A4(KEYINPUT62), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1162), .A2(new_n1163), .A3(new_n1111), .A4(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n963), .A2(new_n1136), .A3(new_n580), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1142), .B1(new_n1147), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1135), .ZN(new_n1170));
  OAI22_X1  g745(.A1(new_n1156), .A2(new_n1150), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT63), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT117), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1125), .A2(new_n1173), .A3(G168), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1173), .B1(new_n1125), .B2(G168), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1172), .B1(new_n1177), .B2(new_n1157), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1134), .A2(new_n1151), .A3(new_n1156), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1176), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1174), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1179), .A2(KEYINPUT63), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1171), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1166), .A2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1035), .B1(new_n1160), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1028), .A2(KEYINPUT46), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT125), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1025), .A2(new_n768), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1023), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1028), .A2(KEYINPUT46), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(KEYINPUT126), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1186), .B(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1194), .A2(new_n1195), .A3(new_n1190), .A4(new_n1189), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1192), .A2(new_n1196), .A3(KEYINPUT47), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT47), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n838), .B(new_n843), .C1(new_n839), .C2(new_n840), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  AOI22_X1  g775(.A1(new_n1029), .A2(new_n1200), .B1(new_n1024), .B2(new_n906), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1022), .A2(G1986), .A3(G290), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT48), .ZN(new_n1203));
  OAI22_X1  g778(.A1(new_n1201), .A2(new_n1030), .B1(new_n1032), .B2(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1197), .A2(new_n1198), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1185), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1208));
  NOR2_X1   g782(.A1(new_n459), .A2(G227), .ZN(new_n1209));
  OAI21_X1  g783(.A(new_n1209), .B1(new_n705), .B2(new_n709), .ZN(new_n1210));
  NOR2_X1   g784(.A1(G401), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n946), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g786(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g787(.A(new_n1208), .B1(new_n1010), .B2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g788(.A(KEYINPUT127), .B(new_n1212), .C1(new_n1004), .C2(new_n1009), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n1214), .A2(new_n1215), .ZN(G308));
  NAND2_X1  g790(.A1(new_n1010), .A2(new_n1213), .ZN(G225));
endmodule


