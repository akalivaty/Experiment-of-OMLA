

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598;

  XNOR2_X1 U327 ( .A(G211GAT), .B(KEYINPUT85), .ZN(n348) );
  XNOR2_X1 U328 ( .A(n428), .B(n427), .ZN(n430) );
  XNOR2_X1 U329 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U330 ( .A(KEYINPUT94), .B(KEYINPUT26), .ZN(n295) );
  XOR2_X1 U331 ( .A(n349), .B(G204GAT), .Z(n296) );
  XNOR2_X1 U332 ( .A(n437), .B(n436), .ZN(n465) );
  INV_X1 U333 ( .A(KEYINPUT95), .ZN(n379) );
  XNOR2_X1 U334 ( .A(n335), .B(KEYINPUT24), .ZN(n336) );
  XNOR2_X1 U335 ( .A(n337), .B(n336), .ZN(n340) );
  XNOR2_X1 U336 ( .A(n469), .B(KEYINPUT47), .ZN(n470) );
  XNOR2_X1 U337 ( .A(n471), .B(n470), .ZN(n476) );
  XNOR2_X1 U338 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U339 ( .A(n419), .B(n369), .ZN(n370) );
  XNOR2_X1 U340 ( .A(n371), .B(n370), .ZN(n375) );
  XNOR2_X1 U341 ( .A(n383), .B(n295), .ZN(n581) );
  XNOR2_X1 U342 ( .A(n418), .B(KEYINPUT37), .ZN(n530) );
  XNOR2_X1 U343 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U344 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U345 ( .A(n496), .B(n495), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT101), .B(KEYINPUT38), .Z(n457) );
  XOR2_X1 U348 ( .A(G85GAT), .B(G92GAT), .Z(n420) );
  XOR2_X1 U349 ( .A(G162GAT), .B(G50GAT), .Z(n334) );
  XOR2_X1 U350 ( .A(G134GAT), .B(G43GAT), .Z(n364) );
  XNOR2_X1 U351 ( .A(n334), .B(n364), .ZN(n299) );
  XOR2_X1 U352 ( .A(G36GAT), .B(KEYINPUT7), .Z(n298) );
  XNOR2_X1 U353 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n297) );
  XNOR2_X1 U354 ( .A(n298), .B(n297), .ZN(n444) );
  XNOR2_X1 U355 ( .A(n299), .B(n444), .ZN(n303) );
  XOR2_X1 U356 ( .A(G190GAT), .B(G106GAT), .Z(n301) );
  NAND2_X1 U357 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U359 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U360 ( .A(G99GAT), .B(KEYINPUT65), .Z(n305) );
  XNOR2_X1 U361 ( .A(KEYINPUT9), .B(KEYINPUT64), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n306), .B(KEYINPUT10), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U365 ( .A(n420), .B(n309), .Z(n311) );
  XNOR2_X1 U366 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n310) );
  XOR2_X1 U367 ( .A(n311), .B(n310), .Z(n570) );
  XNOR2_X1 U368 ( .A(KEYINPUT36), .B(n570), .ZN(n593) );
  XOR2_X1 U369 ( .A(KEYINPUT78), .B(G22GAT), .Z(n313) );
  XNOR2_X1 U370 ( .A(G64GAT), .B(G15GAT), .ZN(n312) );
  XNOR2_X1 U371 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U372 ( .A(KEYINPUT76), .B(KEYINPUT79), .Z(n315) );
  XNOR2_X1 U373 ( .A(G155GAT), .B(KEYINPUT14), .ZN(n314) );
  XNOR2_X1 U374 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U375 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U376 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n319) );
  NAND2_X1 U377 ( .A1(G231GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U378 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U379 ( .A(KEYINPUT15), .B(n320), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n331) );
  XOR2_X1 U381 ( .A(KEYINPUT77), .B(G183GAT), .Z(n324) );
  XNOR2_X1 U382 ( .A(G127GAT), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U383 ( .A(n324), .B(n323), .ZN(n329) );
  XOR2_X1 U384 ( .A(G1GAT), .B(G8GAT), .Z(n451) );
  XOR2_X1 U385 ( .A(n451), .B(G78GAT), .Z(n327) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n325) );
  XNOR2_X1 U387 ( .A(n325), .B(KEYINPUT70), .ZN(n431) );
  XNOR2_X1 U388 ( .A(n431), .B(G71GAT), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U390 ( .A(n329), .B(n328), .Z(n330) );
  XOR2_X1 U391 ( .A(n331), .B(n330), .Z(n489) );
  INV_X1 U392 ( .A(n489), .ZN(n591) );
  XOR2_X1 U393 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n333) );
  XNOR2_X1 U394 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n332) );
  XNOR2_X1 U395 ( .A(n333), .B(n332), .ZN(n394) );
  XNOR2_X1 U396 ( .A(n334), .B(n394), .ZN(n337) );
  AND2_X1 U397 ( .A1(G228GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U398 ( .A(G148GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n338), .B(G78GAT), .ZN(n432) );
  XOR2_X1 U400 ( .A(n432), .B(KEYINPUT22), .Z(n339) );
  XNOR2_X1 U401 ( .A(n340), .B(n339), .ZN(n343) );
  INV_X1 U402 ( .A(n343), .ZN(n341) );
  NAND2_X1 U403 ( .A1(n341), .A2(KEYINPUT87), .ZN(n345) );
  INV_X1 U404 ( .A(KEYINPUT87), .ZN(n342) );
  NAND2_X1 U405 ( .A1(n343), .A2(n342), .ZN(n344) );
  NAND2_X1 U406 ( .A1(n345), .A2(n344), .ZN(n347) );
  XOR2_X1 U407 ( .A(G141GAT), .B(G22GAT), .Z(n441) );
  XNOR2_X1 U408 ( .A(n441), .B(KEYINPUT23), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n348), .B(G197GAT), .ZN(n349) );
  XNOR2_X1 U411 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n350) );
  XOR2_X1 U412 ( .A(n296), .B(n350), .Z(n371) );
  INV_X1 U413 ( .A(n371), .ZN(n351) );
  XOR2_X1 U414 ( .A(n352), .B(n351), .Z(n480) );
  XOR2_X1 U415 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n354) );
  NAND2_X1 U416 ( .A1(G227GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U418 ( .A(KEYINPUT82), .B(n355), .ZN(n368) );
  XOR2_X1 U419 ( .A(G113GAT), .B(G15GAT), .Z(n440) );
  XOR2_X1 U420 ( .A(G127GAT), .B(KEYINPUT0), .Z(n390) );
  XNOR2_X1 U421 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n356), .B(KEYINPUT18), .ZN(n357) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(n357), .ZN(n359) );
  XOR2_X1 U424 ( .A(G190GAT), .B(KEYINPUT19), .Z(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n376) );
  XNOR2_X1 U426 ( .A(n390), .B(n376), .ZN(n361) );
  XOR2_X1 U427 ( .A(KEYINPUT83), .B(G176GAT), .Z(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U429 ( .A(n440), .B(n362), .Z(n366) );
  XNOR2_X1 U430 ( .A(G120GAT), .B(G99GAT), .ZN(n363) );
  XNOR2_X1 U431 ( .A(n363), .B(G71GAT), .ZN(n433) );
  XNOR2_X1 U432 ( .A(n364), .B(n433), .ZN(n365) );
  XNOR2_X1 U433 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U434 ( .A(n368), .B(n367), .ZN(n487) );
  INV_X1 U435 ( .A(n487), .ZN(n410) );
  XOR2_X1 U436 ( .A(G64GAT), .B(G176GAT), .Z(n419) );
  XNOR2_X1 U437 ( .A(G92GAT), .B(G36GAT), .ZN(n369) );
  XOR2_X1 U438 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n373) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n378) );
  XNOR2_X1 U442 ( .A(G8GAT), .B(n376), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n533) );
  NOR2_X1 U444 ( .A1(n410), .A2(n533), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n381) );
  NOR2_X1 U446 ( .A1(n480), .A2(n381), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n382), .B(KEYINPUT25), .ZN(n385) );
  NAND2_X1 U448 ( .A1(n480), .A2(n410), .ZN(n383) );
  XNOR2_X1 U449 ( .A(n533), .B(KEYINPUT27), .ZN(n412) );
  OR2_X1 U450 ( .A1(n581), .A2(n412), .ZN(n384) );
  NAND2_X1 U451 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n386), .B(KEYINPUT96), .ZN(n409) );
  XOR2_X1 U453 ( .A(G85GAT), .B(G134GAT), .Z(n388) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(G162GAT), .ZN(n387) );
  XNOR2_X1 U455 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U456 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U459 ( .A(n393), .B(KEYINPUT89), .Z(n396) );
  XNOR2_X1 U460 ( .A(n394), .B(KEYINPUT90), .ZN(n395) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U462 ( .A(G1GAT), .B(G148GAT), .Z(n398) );
  XNOR2_X1 U463 ( .A(G57GAT), .B(G120GAT), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U465 ( .A(n400), .B(n399), .Z(n408) );
  XOR2_X1 U466 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n402) );
  XNOR2_X1 U467 ( .A(KEYINPUT4), .B(KEYINPUT88), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U469 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n404) );
  XNOR2_X1 U470 ( .A(G113GAT), .B(G141GAT), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U472 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n531) );
  NAND2_X1 U474 ( .A1(n409), .A2(n531), .ZN(n415) );
  XOR2_X1 U475 ( .A(n480), .B(KEYINPUT28), .Z(n538) );
  INV_X1 U476 ( .A(n538), .ZN(n548) );
  INV_X1 U477 ( .A(n487), .ZN(n545) );
  XOR2_X1 U478 ( .A(KEYINPUT84), .B(n545), .Z(n411) );
  NOR2_X1 U479 ( .A1(n548), .A2(n411), .ZN(n413) );
  NOR2_X1 U480 ( .A1(n531), .A2(n412), .ZN(n544) );
  NAND2_X1 U481 ( .A1(n413), .A2(n544), .ZN(n414) );
  NAND2_X1 U482 ( .A1(n415), .A2(n414), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n416), .B(KEYINPUT97), .ZN(n501) );
  NOR2_X1 U484 ( .A1(n591), .A2(n501), .ZN(n417) );
  NAND2_X1 U485 ( .A1(n593), .A2(n417), .ZN(n418) );
  XOR2_X1 U486 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n422) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U488 ( .A(n422), .B(n421), .ZN(n428) );
  XOR2_X1 U489 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n424) );
  XNOR2_X1 U490 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n423) );
  XOR2_X1 U491 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U492 ( .A1(G230GAT), .A2(G233GAT), .ZN(n425) );
  INV_X1 U493 ( .A(KEYINPUT72), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n431), .B(KEYINPUT74), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U497 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n439) );
  XNOR2_X1 U498 ( .A(G50GAT), .B(G43GAT), .ZN(n438) );
  XNOR2_X1 U499 ( .A(n439), .B(n438), .ZN(n455) );
  XOR2_X1 U500 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U501 ( .A1(G229GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U502 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n444), .B(KEYINPUT66), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n445), .B(KEYINPUT67), .ZN(n446) );
  XOR2_X1 U505 ( .A(n447), .B(n446), .Z(n453) );
  XOR2_X1 U506 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n449) );
  XNOR2_X1 U507 ( .A(G169GAT), .B(G197GAT), .ZN(n448) );
  XNOR2_X1 U508 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U511 ( .A(n455), .B(n454), .Z(n582) );
  INV_X1 U512 ( .A(n582), .ZN(n573) );
  NOR2_X1 U513 ( .A1(n465), .A2(n573), .ZN(n502) );
  NAND2_X1 U514 ( .A1(n530), .A2(n502), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U516 ( .A(KEYINPUT100), .B(n458), .ZN(n513) );
  NOR2_X1 U517 ( .A1(n513), .A2(n545), .ZN(n462) );
  XNOR2_X1 U518 ( .A(KEYINPUT40), .B(KEYINPUT102), .ZN(n460) );
  INV_X1 U519 ( .A(G43GAT), .ZN(n459) );
  NOR2_X1 U520 ( .A1(n531), .A2(n513), .ZN(n464) );
  XNOR2_X1 U521 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n464), .B(n463), .ZN(G1328GAT) );
  INV_X1 U523 ( .A(n570), .ZN(n497) );
  XOR2_X1 U524 ( .A(n465), .B(KEYINPUT41), .Z(n562) );
  AND2_X1 U525 ( .A1(n582), .A2(n562), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n466), .B(KEYINPUT46), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n467), .A2(n591), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n497), .A2(n468), .ZN(n471) );
  INV_X1 U529 ( .A(KEYINPUT111), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n593), .A2(n591), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT45), .B(n472), .Z(n473) );
  NAND2_X1 U532 ( .A1(n473), .A2(n573), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n474), .A2(n465), .ZN(n475) );
  NOR2_X1 U534 ( .A1(n476), .A2(n475), .ZN(n542) );
  XNOR2_X1 U535 ( .A(n542), .B(KEYINPUT48), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n477), .A2(n533), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(KEYINPUT54), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n479), .A2(n531), .ZN(n580) );
  NOR2_X1 U539 ( .A1(n480), .A2(n580), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT55), .B(n481), .ZN(n483) );
  INV_X1 U541 ( .A(KEYINPUT118), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n483), .A2(n482), .ZN(n486) );
  INV_X1 U543 ( .A(n483), .ZN(n484) );
  NAND2_X1 U544 ( .A1(KEYINPUT118), .A2(n484), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n488) );
  NAND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n572) );
  NOR2_X1 U547 ( .A1(n572), .A2(n489), .ZN(n492) );
  XNOR2_X1 U548 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(G183GAT), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(G1350GAT) );
  NOR2_X1 U551 ( .A1(n572), .A2(n497), .ZN(n496) );
  XNOR2_X1 U552 ( .A(KEYINPUT122), .B(KEYINPUT58), .ZN(n494) );
  INV_X1 U553 ( .A(G190GAT), .ZN(n493) );
  NAND2_X1 U554 ( .A1(n591), .A2(n497), .ZN(n498) );
  XNOR2_X1 U555 ( .A(n498), .B(KEYINPUT80), .ZN(n499) );
  XNOR2_X1 U556 ( .A(n499), .B(KEYINPUT16), .ZN(n500) );
  NOR2_X1 U557 ( .A1(n501), .A2(n500), .ZN(n519) );
  NAND2_X1 U558 ( .A1(n502), .A2(n519), .ZN(n510) );
  NOR2_X1 U559 ( .A1(n531), .A2(n510), .ZN(n504) );
  XNOR2_X1 U560 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U562 ( .A(G1GAT), .B(n505), .Z(G1324GAT) );
  NOR2_X1 U563 ( .A1(n533), .A2(n510), .ZN(n507) );
  XNOR2_X1 U564 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n507), .B(n506), .ZN(G1325GAT) );
  NOR2_X1 U566 ( .A1(n545), .A2(n510), .ZN(n509) );
  XNOR2_X1 U567 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(G1326GAT) );
  NOR2_X1 U569 ( .A1(n538), .A2(n510), .ZN(n511) );
  XOR2_X1 U570 ( .A(G22GAT), .B(n511), .Z(G1327GAT) );
  NOR2_X1 U571 ( .A1(n533), .A2(n513), .ZN(n512) );
  XOR2_X1 U572 ( .A(G36GAT), .B(n512), .Z(G1329GAT) );
  NOR2_X1 U573 ( .A1(n538), .A2(n513), .ZN(n515) );
  XNOR2_X1 U574 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(G1331GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n517) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(n521) );
  INV_X1 U579 ( .A(n562), .ZN(n575) );
  NOR2_X1 U580 ( .A1(n575), .A2(n582), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(KEYINPUT104), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n519), .A2(n529), .ZN(n525) );
  NOR2_X1 U583 ( .A1(n531), .A2(n525), .ZN(n520) );
  XOR2_X1 U584 ( .A(n521), .B(n520), .Z(G1332GAT) );
  NOR2_X1 U585 ( .A1(n533), .A2(n525), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n523), .B(n522), .ZN(G1333GAT) );
  NOR2_X1 U588 ( .A1(n545), .A2(n525), .ZN(n524) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n524), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n538), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G78GAT), .B(n528), .ZN(G1335GAT) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n537) );
  NOR2_X1 U595 ( .A1(n531), .A2(n537), .ZN(n532) );
  XOR2_X1 U596 ( .A(G85GAT), .B(n532), .Z(G1336GAT) );
  NOR2_X1 U597 ( .A1(n533), .A2(n537), .ZN(n535) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U600 ( .A1(n545), .A2(n537), .ZN(n536) );
  XOR2_X1 U601 ( .A(G99GAT), .B(n536), .Z(G1338GAT) );
  NOR2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U603 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U605 ( .A(G106GAT), .B(n541), .Z(G1339GAT) );
  XOR2_X1 U606 ( .A(n542), .B(KEYINPUT48), .Z(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n560) );
  NOR2_X1 U608 ( .A1(n545), .A2(n560), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT112), .B(n546), .Z(n547) );
  NOR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n556), .A2(n582), .ZN(n549) );
  XNOR2_X1 U612 ( .A(n549), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U614 ( .A1(n556), .A2(n562), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(G120GAT), .B(n552), .Z(G1341GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n554) );
  NAND2_X1 U618 ( .A1(n556), .A2(n591), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U620 ( .A(G127GAT), .B(n555), .Z(G1342GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U622 ( .A1(n556), .A2(n570), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U624 ( .A(G134GAT), .B(n559), .Z(G1343GAT) );
  NOR2_X1 U625 ( .A1(n581), .A2(n560), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n582), .A2(n569), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n561), .ZN(G1344GAT) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n564) );
  NAND2_X1 U630 ( .A1(n569), .A2(n562), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  XOR2_X1 U633 ( .A(G155GAT), .B(KEYINPUT117), .Z(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n591), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(G169GAT), .B(n574), .Z(G1348GAT) );
  NOR2_X1 U640 ( .A1(n572), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n577) );
  XNOR2_X1 U642 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1349GAT) );
  XOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .Z(n584) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n594) );
  NAND2_X1 U647 ( .A1(n594), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n586) );
  XOR2_X1 U649 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n588) );
  NAND2_X1 U652 ( .A1(n594), .A2(n465), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n590) );
  XOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT124), .Z(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  NAND2_X1 U656 ( .A1(n591), .A2(n594), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n592), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n598) );
  XOR2_X1 U659 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n596) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U661 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n598), .B(n597), .ZN(G1355GAT) );
endmodule

