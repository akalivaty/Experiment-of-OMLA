//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n555, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT65), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n462));
  OAI211_X1 g037(.A(new_n462), .B(G125), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G137), .A3(new_n467), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n458), .A2(new_n459), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n467), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n467), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n476), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT66), .ZN(G162));
  NAND3_X1  g059(.A1(new_n470), .A2(G126), .A3(G2105), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT67), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n467), .A2(G114), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n491), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n485), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n467), .A3(G138), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n474), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n496), .A2(new_n467), .A3(G138), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT68), .B1(new_n470), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n467), .C1(new_n458), .C2(new_n459), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n494), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .A3(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(G50), .A3(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n511), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n520), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(new_n521), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n506), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n515), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT7), .Z(new_n530));
  AND3_X1   g105(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n531));
  AOI211_X1 g106(.A(new_n530), .B(new_n531), .C1(new_n523), .C2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n512), .A2(KEYINPUT72), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n516), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n533), .A2(G51), .A3(G543), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND3_X1  g113(.A1(new_n533), .A2(G543), .A3(new_n535), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT73), .B(G52), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n523), .A2(G90), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n506), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(new_n523), .A2(G81), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n522), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n539), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(G43), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  AND2_X1   g134(.A1(G53), .A2(G543), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n533), .A2(new_n535), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(KEYINPUT75), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n522), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(G91), .A2(new_n523), .B1(new_n566), .B2(G651), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n533), .A2(new_n570), .A3(new_n535), .A4(new_n560), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  OR2_X1    g149(.A1(new_n515), .A2(new_n527), .ZN(G303));
  NAND4_X1  g150(.A1(new_n533), .A2(G49), .A3(G543), .A4(new_n535), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n525), .A2(G74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n523), .A2(G87), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n522), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(G48), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n522), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(new_n512), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n506), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n523), .A2(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n539), .ZN(G290));
  NAND4_X1  g171(.A1(new_n510), .A2(new_n525), .A3(G92), .A4(new_n511), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n533), .A2(G54), .A3(G543), .A4(new_n535), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n525), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n506), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G284));
  OAI21_X1  g181(.A(new_n605), .B1(G171), .B2(new_n604), .ZN(G321));
  NOR2_X1   g182(.A1(G286), .A2(new_n604), .ZN(new_n608));
  XOR2_X1   g183(.A(G299), .B(KEYINPUT76), .Z(new_n609));
  AOI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n604), .ZN(G297));
  AOI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n604), .ZN(G280));
  INV_X1    g186(.A(G860), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n603), .B1(G559), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT77), .ZN(G148));
  AND2_X1   g189(.A1(new_n546), .A2(new_n550), .ZN(new_n615));
  INV_X1    g190(.A(G43), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n539), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(new_n604), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n603), .A2(G559), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n618), .B1(new_n620), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n475), .A2(G135), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT79), .Z(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(G123), .B2(new_n479), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n470), .A2(new_n468), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT12), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2100), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(G2096), .ZN(new_n639));
  NAND4_X1  g214(.A1(new_n632), .A2(new_n637), .A3(new_n638), .A4(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n646), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT81), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n650), .A2(new_n654), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n662), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n662), .A2(KEYINPUT83), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(KEYINPUT83), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n661), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n662), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(new_n631), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT85), .B(G2100), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT20), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n680), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n680), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G229));
  INV_X1    g270(.A(G29), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G25), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n479), .A2(G119), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT86), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n475), .A2(G131), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n467), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n700), .B(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT87), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n698), .B1(new_n705), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n706), .B(new_n708), .Z(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G24), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n593), .B1(new_n552), .B2(G47), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1986), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G1971), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n710), .A2(G22), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G303), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n716), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OR2_X1    g298(.A1(G16), .A2(G23), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n576), .A2(new_n578), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(G288), .A2(KEYINPUT90), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n724), .B1(new_n729), .B2(new_n710), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT33), .B(G1976), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n718), .A2(new_n719), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n733), .A2(G1971), .A3(new_n720), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n588), .A2(G16), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G6), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT32), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1981), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n736), .A2(KEYINPUT32), .ZN(new_n739));
  INV_X1    g314(.A(G1981), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n736), .A2(KEYINPUT32), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n723), .A2(new_n732), .A3(new_n734), .A4(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n715), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(KEYINPUT93), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT92), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n744), .B2(new_n746), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n744), .A2(new_n751), .A3(new_n746), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n748), .B(new_n750), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G35), .ZN(new_n756));
  OR3_X1    g331(.A1(new_n756), .A2(KEYINPUT103), .A3(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT103), .B1(new_n756), .B2(G29), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n757), .B(new_n758), .C1(G162), .C2(new_n696), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT29), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(G2090), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT104), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n553), .B2(G16), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT94), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(G1341), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G1341), .B2(new_n766), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n630), .A2(G29), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT101), .ZN(new_n770));
  NOR2_X1   g345(.A1(G27), .A2(G29), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G164), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n696), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n475), .A2(G140), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n479), .A2(G128), .ZN(new_n778));
  OR2_X1    g353(.A1(G104), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(new_n696), .ZN(new_n783));
  INV_X1    g358(.A(G2067), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n770), .A2(new_n774), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(G28), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n696), .B1(new_n787), .B2(G28), .ZN(new_n789));
  AND2_X1   g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NOR2_X1   g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  OAI22_X1  g366(.A1(new_n788), .A2(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT25), .ZN(new_n793));
  NAND2_X1  g368(.A1(G103), .A2(G2104), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(G2105), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n475), .A2(G139), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n467), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n696), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n696), .B2(G33), .ZN(new_n802));
  INV_X1    g377(.A(G2072), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n792), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G2084), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n696), .B1(KEYINPUT24), .B2(G34), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(KEYINPUT24), .B2(G34), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n472), .B2(G29), .ZN(new_n808));
  OAI221_X1 g383(.A(new_n804), .B1(new_n803), .B2(new_n802), .C1(new_n805), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G5), .A2(G16), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G171), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1961), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n786), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT27), .B(G1996), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n475), .A2(G141), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT95), .ZN(new_n818));
  NAND3_X1  g393(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT96), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT26), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n479), .A2(G129), .B1(G105), .B2(new_n468), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n818), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n696), .ZN(new_n824));
  NOR2_X1   g399(.A1(G29), .A2(G32), .ZN(new_n825));
  OR3_X1    g400(.A1(new_n824), .A2(KEYINPUT97), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(KEYINPUT97), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n816), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n710), .A2(G21), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(G168), .B2(new_n710), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT100), .B(G1966), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n832), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n828), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n826), .A2(new_n816), .A3(new_n827), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n761), .A2(new_n762), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n813), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G4), .A2(G16), .ZN(new_n840));
  INV_X1    g415(.A(new_n603), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(G16), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n760), .A2(G2090), .B1(G1348), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n808), .A2(new_n805), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT102), .Z(new_n845));
  INV_X1    g420(.A(G1348), .ZN(new_n846));
  INV_X1    g421(.A(new_n842), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n710), .A2(G20), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT23), .Z(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G299), .B2(G16), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G1956), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n843), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n768), .A2(new_n839), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n754), .A2(new_n752), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n855), .A2(new_n747), .ZN(new_n856));
  XOR2_X1   g431(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n857));
  OAI211_X1 g432(.A(new_n755), .B(new_n854), .C1(new_n856), .C2(new_n857), .ZN(G150));
  INV_X1    g433(.A(G150), .ZN(G311));
  NAND2_X1  g434(.A1(G80), .A2(G543), .ZN(new_n860));
  INV_X1    g435(.A(G67), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n522), .B2(new_n861), .ZN(new_n862));
  AOI22_X1  g437(.A1(G93), .A2(new_n523), .B1(new_n862), .B2(G651), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n533), .A2(G55), .A3(G543), .A4(new_n535), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n841), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n617), .A2(new_n865), .ZN(new_n870));
  INV_X1    g445(.A(new_n865), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n553), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n869), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT105), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n612), .B1(new_n875), .B2(KEYINPUT39), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n867), .B1(new_n877), .B2(new_n878), .ZN(G145));
  XNOR2_X1  g454(.A(new_n629), .B(KEYINPUT106), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G160), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n823), .B(new_n800), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n475), .A2(G142), .B1(G130), .B2(new_n479), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n467), .A2(KEYINPUT107), .A3(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT107), .B1(new_n467), .B2(G118), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n884), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n634), .Z(new_n889));
  XNOR2_X1  g464(.A(new_n883), .B(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n495), .B1(new_n474), .B2(new_n497), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n470), .A2(new_n499), .A3(KEYINPUT68), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n503), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n487), .A2(KEYINPUT67), .A3(new_n489), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n492), .B1(new_n491), .B2(new_n486), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n894), .A2(new_n895), .B1(new_n479), .B2(G126), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n782), .B(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n705), .B(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n890), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n890), .A2(new_n899), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n882), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n882), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(G37), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n907));
  NOR2_X1   g482(.A1(G290), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n909));
  OAI21_X1  g484(.A(G166), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(G290), .A2(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(G303), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n729), .A2(new_n588), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n727), .A2(G305), .A3(new_n728), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n910), .A2(new_n915), .A3(new_n913), .A4(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n568), .A2(new_n572), .A3(new_n841), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n841), .B1(new_n568), .B2(new_n572), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT41), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(G299), .A2(new_n603), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n568), .A2(new_n572), .A3(new_n841), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(new_n929), .A3(KEYINPUT108), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n923), .A2(new_n924), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n927), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n873), .A2(new_n620), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n619), .A2(new_n870), .A3(new_n872), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT110), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(KEYINPUT110), .A3(new_n938), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n922), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n920), .B(KEYINPUT42), .ZN(new_n943));
  INV_X1    g518(.A(new_n941), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(G868), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT111), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n871), .A2(G868), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n943), .B1(new_n944), .B2(new_n939), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n922), .A2(new_n941), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n604), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT111), .B1(new_n953), .B2(new_n948), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(G295));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n949), .ZN(G331));
  NOR2_X1   g531(.A1(new_n617), .A2(new_n865), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n552), .A2(G43), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n958), .A2(new_n615), .B1(new_n864), .B2(new_n863), .ZN(new_n959));
  OAI21_X1  g534(.A(G168), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n870), .A2(new_n872), .A3(G286), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(G171), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n961), .ZN(new_n963));
  AOI21_X1  g538(.A(G286), .B1(new_n870), .B2(new_n872), .ZN(new_n964));
  OAI21_X1  g539(.A(G301), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n930), .A2(new_n933), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n960), .A2(G171), .A3(new_n961), .ZN(new_n967));
  AOI21_X1  g542(.A(G171), .B1(new_n960), .B2(new_n961), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n931), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n920), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n904), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n925), .A2(new_n929), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n962), .A3(new_n965), .ZN(new_n973));
  AOI211_X1 g548(.A(KEYINPUT112), .B(new_n920), .C1(new_n973), .C2(new_n969), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n969), .ZN(new_n976));
  INV_X1    g551(.A(new_n920), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT43), .ZN(new_n979));
  NOR4_X1   g554(.A1(new_n971), .A2(new_n974), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n971), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n966), .A2(new_n969), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n977), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT43), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT44), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n986));
  NOR4_X1   g561(.A1(new_n971), .A2(new_n974), .A3(new_n978), .A4(KEYINPUT43), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n979), .B1(new_n981), .B2(new_n983), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n989), .ZN(G397));
  AOI21_X1  g565(.A(G1384), .B1(new_n893), .B2(new_n896), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(KEYINPUT113), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n991), .B2(KEYINPUT113), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n471), .A2(G40), .A3(new_n469), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n465), .B2(G2105), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n705), .B(new_n708), .Z(new_n1000));
  XNOR2_X1  g575(.A(new_n823), .B(G1996), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n781), .B(new_n784), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1000), .A2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(G290), .A2(G1986), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G290), .A2(G1986), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n999), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT123), .B1(G286), .B2(G8), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT123), .ZN(new_n1011));
  INV_X1    g586(.A(G8), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1011), .B(new_n1012), .C1(new_n532), .C2(new_n536), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n993), .A2(G1384), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n997), .B1(G164), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n831), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n897), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(new_n996), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n466), .A2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n893), .B2(new_n896), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1027), .A3(new_n805), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1012), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT124), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1014), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g606(.A(KEYINPUT124), .B(new_n1012), .C1(new_n1019), .C2(new_n1028), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT125), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT125), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1035), .B(KEYINPUT51), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1014), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1037), .A2(KEYINPUT51), .A3(new_n1029), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1014), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT126), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1038), .B1(new_n1033), .B2(KEYINPUT125), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1041), .B1(new_n1046), .B2(new_n1036), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT62), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(G2090), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1022), .A2(new_n1027), .A3(KEYINPUT115), .A4(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT114), .B(G1971), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1052), .A2(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1012), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT116), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G166), .A2(new_n1012), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1060), .A2(new_n1063), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1069), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1051), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1056), .A2(new_n1057), .B1(new_n1072), .B2(new_n1053), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1012), .B2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n727), .A2(G1976), .A3(new_n728), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n991), .A2(new_n997), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n1012), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT52), .ZN(new_n1080));
  INV_X1    g655(.A(G1976), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT52), .B1(G288), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT118), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1078), .A3(new_n1075), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G305), .A2(G1981), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n588), .A2(new_n740), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(KEYINPUT49), .A3(new_n1088), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1078), .A3(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1080), .A2(new_n1086), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT53), .B1(new_n1055), .B2(new_n773), .ZN(new_n1095));
  INV_X1    g670(.A(G1961), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1096), .B2(new_n1051), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1055), .A2(KEYINPUT53), .A3(new_n773), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1070), .A2(new_n1074), .A3(new_n1094), .A4(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1044), .A2(new_n1049), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1029), .A2(G168), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1070), .A2(new_n1074), .A3(new_n1094), .A4(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT63), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1071), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1103), .A2(KEYINPUT63), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(new_n1070), .A3(new_n1094), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1107), .A2(new_n1071), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1093), .A2(new_n1081), .A3(new_n725), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1088), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1112), .A2(new_n1094), .B1(new_n1078), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  INV_X1    g691(.A(G1956), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1055), .A2(new_n1116), .B1(new_n1051), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(KEYINPUT120), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n567), .A2(KEYINPUT119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(KEYINPUT57), .ZN(new_n1121));
  NAND2_X1  g696(.A1(G299), .A2(new_n1121), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n568), .B(new_n572), .C1(KEYINPUT57), .C2(new_n1120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1118), .A2(KEYINPUT120), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1124), .A2(new_n1118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1051), .A2(new_n846), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1077), .A2(new_n784), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n603), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1125), .A2(new_n1126), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n1124), .B2(new_n1118), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1127), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1124), .A2(new_n1118), .A3(new_n1132), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1128), .A2(new_n603), .A3(new_n1129), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1130), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n603), .A2(KEYINPUT60), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1128), .A2(new_n1129), .A3(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(KEYINPUT58), .B(G1341), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1076), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1076), .A2(KEYINPUT122), .A3(new_n1141), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT121), .B(G1996), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1144), .B(new_n1145), .C1(new_n1056), .C2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1147), .A2(new_n1148), .A3(new_n553), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1147), .B2(new_n553), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1138), .B(new_n1140), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1131), .B1(new_n1136), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1070), .A2(new_n1074), .A3(new_n1094), .ZN(new_n1153));
  XOR2_X1   g728(.A(G171), .B(KEYINPUT54), .Z(new_n1154));
  INV_X1    g729(.A(new_n995), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1017), .A2(new_n1156), .A3(G2078), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1154), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1158), .A2(new_n1097), .B1(new_n1159), .B2(new_n1154), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1152), .A2(new_n1153), .A3(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1111), .B(new_n1115), .C1(new_n1161), .C2(new_n1047), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1009), .B1(new_n1102), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n705), .A2(new_n708), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1004), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n782), .A2(new_n784), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n998), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1006), .A2(new_n998), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1005), .A2(new_n999), .B1(KEYINPUT48), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1168), .A2(KEYINPUT48), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n998), .A2(G1996), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT46), .Z(new_n1173));
  OAI21_X1  g748(.A(new_n999), .B1(new_n823), .B2(new_n1003), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AND2_X1   g750(.A1(new_n1175), .A2(KEYINPUT47), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(KEYINPUT47), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT127), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1163), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g755(.A(G319), .B1(new_n656), .B2(new_n657), .ZN(new_n1182));
  NOR3_X1   g756(.A1(G229), .A2(G227), .A3(new_n1182), .ZN(new_n1183));
  OAI211_X1 g757(.A(new_n905), .B(new_n1183), .C1(new_n987), .C2(new_n988), .ZN(G225));
  INV_X1    g758(.A(G225), .ZN(G308));
endmodule


