//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n588, new_n589,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  AND2_X1   g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(new_n462));
  OAI21_X1  g037(.A(G2105), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(new_n459), .B(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n472), .ZN(new_n477));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI22_X1  g055(.A1(new_n477), .A2(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n476), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n476), .B2(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n481), .B1(new_n486), .B2(G124), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT71), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NOR2_X1   g064(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT73), .A2(KEYINPUT4), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n491), .A2(G138), .A3(new_n472), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n469), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n490), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n459), .A2(new_n494), .A3(new_n491), .A4(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n472), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n459), .B2(new_n504), .ZN(new_n505));
  AND4_X1   g080(.A1(new_n503), .A2(new_n466), .A3(new_n468), .A4(new_n504), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT74), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n466), .A2(new_n468), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n466), .A2(new_n468), .A3(new_n504), .A4(new_n503), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n496), .A2(new_n466), .A3(new_n468), .A4(new_n491), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n500), .B1(new_n513), .B2(new_n490), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n512), .A2(new_n514), .A3(new_n515), .A4(new_n497), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n508), .A2(new_n516), .ZN(G164));
  INV_X1    g092(.A(KEYINPUT75), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT75), .A3(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n520), .A2(new_n522), .B1(KEYINPUT6), .B2(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT76), .A2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G50), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n529), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n525), .A2(new_n527), .ZN(new_n535));
  INV_X1    g110(.A(G62), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n533), .A2(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  NAND3_X1  g116(.A1(new_n528), .A2(G63), .A3(G651), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT77), .Z(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT78), .B(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n544), .B(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n523), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n546), .B1(G51), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n523), .A2(new_n528), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G89), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n543), .A2(new_n548), .A3(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  NAND2_X1  g127(.A1(new_n549), .A2(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n547), .A2(G52), .ZN(new_n554));
  NAND2_X1  g129(.A1(G77), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G64), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n535), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n553), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G171));
  AOI22_X1  g135(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n519), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n549), .A2(G81), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n547), .A2(G43), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  AND3_X1   g142(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G36), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(G188));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n547), .A2(new_n573), .A3(G53), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT79), .B1(new_n531), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(KEYINPUT9), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n535), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n549), .A2(G91), .B1(new_n581), .B2(G651), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT9), .ZN(new_n583));
  OAI211_X1 g158(.A(KEYINPUT79), .B(new_n583), .C1(new_n531), .C2(new_n575), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n559), .B(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G301));
  NAND2_X1  g165(.A1(new_n547), .A2(G49), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n549), .A2(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(G288));
  AOI22_X1  g169(.A1(G86), .A2(new_n549), .B1(new_n547), .B2(G48), .ZN(new_n595));
  NAND2_X1  g170(.A1(G73), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G61), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n535), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n599), .A2(KEYINPUT81), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n599), .A2(KEYINPUT81), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n549), .A2(G85), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT82), .B(G47), .Z(new_n605));
  OAI221_X1 g180(.A(new_n603), .B1(new_n519), .B2(new_n604), .C1(new_n531), .C2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT84), .B(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n535), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n519), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(new_n609), .ZN(new_n612));
  AND3_X1   g187(.A1(new_n523), .A2(G92), .A3(new_n528), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n614));
  AOI22_X1  g189(.A1(new_n613), .A2(new_n614), .B1(new_n547), .B2(G54), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n589), .B2(new_n618), .ZN(G284));
  OAI21_X1  g195(.A(new_n619), .B1(new_n589), .B2(new_n618), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n586), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G868), .B2(new_n586), .ZN(G280));
  INV_X1    g199(.A(new_n617), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT86), .B(G559), .Z(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(G860), .B2(new_n626), .ZN(G148));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n486), .A2(G123), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n476), .A2(G135), .A3(new_n472), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT87), .Z(new_n634));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n635), .A2(new_n472), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n472), .B2(G111), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G2104), .A3(new_n638), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n632), .B(new_n634), .C1(new_n636), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n465), .A2(G2105), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n459), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(new_n646), .ZN(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2438), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(KEYINPUT14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT89), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2084), .B(G2090), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT90), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(KEYINPUT17), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n673));
  AOI211_X1 g248(.A(new_n668), .B(new_n672), .C1(new_n671), .C2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n670), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  OAI221_X1 g265(.A(new_n687), .B1(new_n685), .B2(new_n683), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n690), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT91), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n700), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(G1971), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(G1971), .ZN(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT32), .B(G1981), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(new_n705), .B2(new_n706), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G23), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT92), .Z(new_n710));
  INV_X1    g285(.A(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g286(.A1(G288), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n592), .A2(new_n591), .A3(KEYINPUT93), .A4(new_n593), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n710), .B1(new_n714), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n708), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT34), .Z(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  INV_X1    g296(.A(G131), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n472), .A2(G107), .ZN(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n724));
  OAI22_X1  g299(.A1(new_n477), .A2(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n486), .B2(G119), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(new_n720), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT35), .B(G1991), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G24), .B(G290), .S(G16), .Z(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G1986), .Z(new_n732));
  NAND3_X1  g307(.A1(new_n719), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT36), .ZN(new_n734));
  NOR2_X1   g309(.A1(G29), .A2(G35), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G162), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT29), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G2090), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT31), .B(G11), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT98), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n741), .A2(G28), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n720), .B1(new_n741), .B2(G28), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT24), .ZN(new_n744));
  INV_X1    g319(.A(G34), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n744), .B2(new_n745), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n720), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n740), .B1(new_n742), .B2(new_n743), .C1(new_n748), .C2(G2084), .ZN(new_n749));
  NAND2_X1  g324(.A1(G168), .A2(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G16), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n749), .B(new_n754), .C1(G2084), .C2(new_n748), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n700), .A2(G19), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n566), .B2(new_n700), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n755), .B1(new_n720), .B2(new_n640), .C1(G1341), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G27), .A2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G164), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n625), .A2(new_n700), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G4), .B2(new_n700), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n761), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n767), .A2(G2072), .B1(G29), .B2(G33), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n642), .A2(G103), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  INV_X1    g346(.A(G139), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n770), .B1(new_n472), .B2(new_n771), .C1(new_n477), .C2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT96), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n768), .B1(new_n775), .B2(G29), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(KEYINPUT97), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G29), .A2(G32), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT26), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n783), .A2(new_n784), .B1(G105), .B2(new_n642), .ZN(new_n785));
  INV_X1    g360(.A(G141), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n477), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n486), .B2(G129), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n780), .B1(new_n788), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT27), .B(G1996), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n776), .A2(new_n767), .A3(G2072), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n779), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n751), .A2(new_n752), .B1(new_n757), .B2(G1341), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n758), .A2(new_n766), .A3(new_n793), .A4(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(G128), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n485), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G140), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n472), .A2(G116), .ZN(new_n804));
  OAI21_X1  g379(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n805));
  OAI22_X1  g380(.A1(new_n477), .A2(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G29), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n720), .A2(G26), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT95), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G2067), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT23), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n700), .A2(G20), .ZN(new_n818));
  AOI211_X1 g393(.A(new_n817), .B(new_n818), .C1(G299), .C2(G16), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT99), .B(G1956), .Z(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n816), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n734), .A2(new_n738), .A3(new_n800), .A4(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NAND2_X1  g402(.A1(new_n549), .A2(G93), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n547), .A2(G55), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n828), .B(new_n829), .C1(new_n519), .C2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n566), .B1(KEYINPUT100), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(KEYINPUT100), .B2(new_n831), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n565), .A2(new_n831), .A3(KEYINPUT100), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n625), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n831), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(new_n640), .B(new_n474), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n808), .A2(new_n788), .ZN(new_n848));
  INV_X1    g423(.A(new_n788), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(new_n807), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n512), .A2(new_n514), .A3(new_n497), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n848), .B2(new_n850), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n775), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n855), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n857), .A2(new_n853), .A3(new_n773), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n726), .B(new_n644), .ZN(new_n859));
  OR2_X1    g434(.A1(G106), .A2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n861));
  INV_X1    g436(.A(G142), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n477), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n486), .A2(G130), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n859), .B(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n856), .A2(new_n858), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n868), .B1(new_n856), .B2(new_n858), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n488), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n874), .A2(new_n870), .A3(G162), .A4(new_n869), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n847), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n875), .A3(new_n847), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g456(.A1(new_n831), .A2(new_n618), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n835), .B(new_n628), .Z(new_n884));
  XNOR2_X1  g459(.A(new_n586), .B(new_n617), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT104), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n885), .B(KEYINPUT41), .Z(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n883), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n883), .B2(new_n887), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n714), .B(G303), .ZN(new_n892));
  XOR2_X1   g467(.A(G305), .B(G290), .Z(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT42), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n891), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n882), .B1(new_n896), .B2(new_n618), .ZN(G295));
  OAI21_X1  g472(.A(new_n882), .B1(new_n896), .B2(new_n618), .ZN(G331));
  MUX2_X1   g473(.A(new_n589), .B(new_n559), .S(G286), .Z(new_n899));
  OR2_X1    g474(.A1(new_n835), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n835), .A2(new_n899), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n885), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT106), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n900), .A2(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n888), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n903), .A3(new_n888), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n894), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n878), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n894), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n906), .B(KEYINPUT107), .C1(new_n886), .C2(new_n905), .ZN(new_n913));
  INV_X1    g488(.A(new_n894), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n905), .A2(KEYINPUT107), .A3(new_n886), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n878), .A4(new_n909), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n878), .A3(new_n909), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n910), .A2(new_n911), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n924), .B(KEYINPUT44), .C1(new_n925), .C2(KEYINPUT43), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n923), .A2(KEYINPUT108), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n921), .B1(new_n926), .B2(new_n927), .ZN(G397));
  AND3_X1   g503(.A1(new_n493), .A2(new_n497), .A3(new_n501), .ZN(new_n929));
  AOI21_X1  g504(.A(G1384), .B1(new_n929), .B2(new_n512), .ZN(new_n930));
  XOR2_X1   g505(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n463), .A2(new_n473), .A3(G40), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n807), .B(G2067), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n788), .B(G1996), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n726), .B(new_n729), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g515(.A1(G290), .A2(G1986), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT110), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(G1986), .B2(G290), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(G1986), .A3(G290), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n935), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n934), .B1(new_n930), .B2(KEYINPUT45), .ZN(new_n949));
  INV_X1    g524(.A(G2078), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n508), .A2(new_n952), .A3(new_n516), .ZN(new_n953));
  INV_X1    g528(.A(new_n931), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT53), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n952), .B1(new_n502), .B2(new_n507), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n463), .A2(new_n473), .A3(G40), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(KEYINPUT114), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT114), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT45), .B1(new_n851), .B2(new_n952), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n934), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n508), .A2(new_n952), .A3(new_n516), .A4(new_n931), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n962), .A2(new_n965), .A3(new_n950), .A4(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n957), .B1(new_n967), .B2(KEYINPUT121), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT114), .B1(new_n960), .B2(new_n961), .ZN(new_n969));
  INV_X1    g544(.A(new_n966), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT121), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n950), .A4(new_n962), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n934), .B1(new_n930), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(G1961), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT122), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n974), .A2(KEYINPUT122), .A3(new_n980), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n956), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT123), .B1(new_n985), .B2(G301), .ZN(new_n986));
  INV_X1    g561(.A(new_n956), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT122), .B1(new_n974), .B2(new_n980), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n982), .B(new_n979), .C1(new_n968), .C2(new_n973), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT123), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n589), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n951), .A2(KEYINPUT53), .A3(new_n933), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n987), .A2(new_n980), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n994), .A2(new_n589), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n986), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n961), .A2(new_n930), .A3(new_n815), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT117), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n975), .A2(new_n978), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n764), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n934), .B1(new_n958), .B2(new_n976), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(new_n953), .B2(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(G1956), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n578), .B2(new_n585), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n577), .A2(KEYINPUT57), .A3(new_n584), .A4(new_n582), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT56), .B(G2072), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n955), .A2(new_n949), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1008), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1004), .A2(new_n1015), .A3(new_n625), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1008), .A2(new_n1014), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1012), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT60), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n625), .B1(new_n1004), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1001), .A2(new_n1003), .A3(KEYINPUT60), .A4(new_n617), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1022), .A2(new_n1023), .B1(new_n1021), .B2(new_n1004), .ZN(new_n1024));
  INV_X1    g599(.A(G1996), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n955), .A2(new_n1025), .A3(new_n949), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n955), .A2(KEYINPUT118), .A3(new_n949), .A4(new_n1025), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n961), .A2(new_n930), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT58), .B(G1341), .Z(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n566), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(KEYINPUT59), .A3(new_n566), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1008), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1012), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1019), .A2(KEYINPUT61), .A3(new_n1015), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1036), .A2(new_n1037), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1024), .B1(new_n1043), .B2(KEYINPUT119), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1045), .A2(new_n1046), .A3(new_n1037), .A4(new_n1036), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1020), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n994), .B2(G171), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n990), .B2(new_n589), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n712), .B2(new_n713), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1030), .A2(G8), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1057), .B(KEYINPUT55), .Z(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT111), .B(G1971), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n955), .B2(new_n949), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1002), .A2(G2090), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1058), .B(G8), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n595), .A2(new_n599), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G1981), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(G305), .B2(G1981), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT49), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1054), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1052), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1067), .A2(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1006), .A2(G2090), .ZN(new_n1072));
  OAI21_X1  g647(.A(G8), .B1(new_n1072), .B2(new_n1060), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1057), .B(KEYINPUT55), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1056), .A2(new_n1062), .A3(new_n1071), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1002), .B2(G2084), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n965), .A2(new_n966), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n964), .A2(new_n963), .A3(new_n934), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n752), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G2084), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n975), .A2(KEYINPUT115), .A3(new_n978), .A4(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1077), .B(G8), .C1(new_n1085), .C2(G286), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G168), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1085), .B2(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT51), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1076), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1051), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1048), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n999), .A2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g671(.A(G1976), .B(G288), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1097));
  NOR2_X1   g672(.A1(G305), .A2(G1981), .ZN(new_n1098));
  OAI211_X1 g673(.A(G8), .B(new_n1030), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1056), .A2(new_n1071), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1062), .B2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1102));
  NAND3_X1  g677(.A1(new_n1085), .A2(G8), .A3(G168), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(new_n1076), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1056), .A2(new_n1062), .A3(new_n1071), .ZN(new_n1105));
  OAI21_X1  g680(.A(G8), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1074), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT63), .ZN(new_n1108));
  OR3_X1    g683(.A1(new_n1105), .A2(new_n1103), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1101), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1096), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n986), .A2(new_n992), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1077), .B(new_n1088), .C1(new_n1085), .C2(G8), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT62), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1092), .A2(new_n1117), .A3(new_n1089), .A4(new_n1086), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1076), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1112), .A2(new_n1113), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1113), .B1(new_n1112), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n948), .B1(new_n1111), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n935), .A2(new_n1025), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT46), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n936), .A2(new_n788), .ZN(new_n1127));
  INV_X1    g702(.A(new_n935), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT47), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n941), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT48), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n726), .A2(new_n729), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n938), .A2(new_n1133), .B1(G2067), .B2(new_n808), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n940), .A2(new_n1132), .B1(new_n1134), .B2(new_n935), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT125), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1124), .A2(KEYINPUT126), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1110), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1141), .B1(new_n999), .B2(new_n1095), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n990), .A2(new_n991), .A3(new_n589), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n991), .B1(new_n990), .B2(new_n589), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT124), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1112), .A2(new_n1120), .A3(new_n1113), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n947), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1140), .B1(new_n1150), .B2(new_n1137), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1139), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g727(.A(G319), .ZN(new_n1154));
  NOR4_X1   g728(.A1(G229), .A2(new_n1154), .A3(G401), .A4(G227), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n879), .A2(new_n878), .ZN(new_n1156));
  OAI211_X1 g730(.A(new_n919), .B(new_n1155), .C1(new_n1156), .C2(new_n876), .ZN(G225));
  NAND2_X1  g731(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1158));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n1159));
  NAND4_X1  g733(.A1(new_n880), .A2(new_n1159), .A3(new_n919), .A4(new_n1155), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1160), .ZN(G308));
endmodule


