//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n589, new_n592, new_n594, new_n595, new_n596, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT69), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n466), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n469), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n469), .B2(new_n473), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n472), .B1(new_n479), .B2(G2105), .ZN(G160));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n464), .A2(new_n467), .A3(new_n469), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n470), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(G136), .B2(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(new_n468), .A2(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n489), .B1(new_n475), .B2(new_n476), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n464), .A2(new_n467), .A3(G126), .A4(new_n469), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n464), .A2(new_n467), .A3(new_n469), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G102), .A2(G2104), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n468), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n492), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n507), .B2(KEYINPUT70), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(G88), .A2(new_n515), .B1(new_n517), .B2(G50), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n512), .A2(new_n518), .ZN(G166));
  XOR2_X1   g094(.A(KEYINPUT71), .B(G89), .Z(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n514), .A2(new_n520), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n522), .A2(new_n526), .ZN(G168));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n504), .A2(new_n505), .ZN(new_n530));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n534), .B1(new_n533), .B2(new_n532), .ZN(new_n535));
  AOI22_X1  g110(.A1(G90), .A2(new_n515), .B1(new_n517), .B2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(G81), .A2(new_n515), .B1(new_n517), .B2(G43), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n544));
  XOR2_X1   g119(.A(new_n544), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  NAND2_X1  g123(.A1(new_n517), .A2(G53), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT9), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n515), .A2(G91), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n550), .B(new_n551), .C1(new_n528), .C2(new_n552), .ZN(G299));
  INV_X1    g128(.A(G168), .ZN(G286));
  INV_X1    g129(.A(G166), .ZN(G303));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n515), .A2(new_n556), .A3(G87), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n556), .B1(new_n515), .B2(G87), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n506), .A2(G74), .ZN(new_n560));
  AOI22_X1  g135(.A1(G651), .A2(new_n560), .B1(new_n517), .B2(G49), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(G288));
  NAND2_X1  g137(.A1(new_n506), .A2(G61), .ZN(new_n563));
  NAND2_X1  g138(.A1(G73), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n528), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n506), .A2(new_n513), .A3(G86), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G305));
  AOI22_X1  g145(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n528), .ZN(new_n572));
  INV_X1    g147(.A(G85), .ZN(new_n573));
  INV_X1    g148(.A(G47), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n514), .A2(new_n573), .B1(new_n516), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G290));
  INV_X1    g152(.A(G868), .ZN(new_n578));
  NOR2_X1   g153(.A1(G301), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n517), .A2(G54), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT10), .B1(new_n515), .B2(G92), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n580), .B1(new_n528), .B2(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT76), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n579), .B1(new_n586), .B2(new_n578), .ZN(G284));
  AOI21_X1  g162(.A(new_n579), .B1(new_n586), .B2(new_n578), .ZN(G321));
  NAND2_X1  g163(.A1(G299), .A2(new_n578), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(new_n578), .B2(G168), .ZN(G297));
  OAI21_X1  g165(.A(new_n589), .B1(new_n578), .B2(G168), .ZN(G280));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n586), .B1(new_n592), .B2(G860), .ZN(G148));
  OAI21_X1  g168(.A(KEYINPUT77), .B1(new_n542), .B2(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n586), .A2(new_n592), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G868), .ZN(new_n596));
  MUX2_X1   g171(.A(KEYINPUT77), .B(new_n594), .S(new_n596), .Z(G323));
  XNOR2_X1  g172(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g173(.A(G123), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n468), .A2(G111), .ZN(new_n600));
  OAI21_X1  g175(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n601));
  OAI22_X1  g176(.A1(new_n484), .A2(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(G135), .B2(new_n487), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT81), .Z(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(G2096), .Z(new_n605));
  NOR2_X1   g180(.A1(new_n466), .A2(G2104), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT68), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n469), .A2(new_n473), .A3(new_n474), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n462), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(KEYINPUT80), .B(G2100), .Z(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n613), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n605), .A2(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT83), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2427), .B(G2430), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n623), .A2(KEYINPUT14), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(G1341), .B(G1348), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n625), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G14), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n629), .A2(new_n632), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(G401));
  XNOR2_X1  g211(.A(G2072), .B(G2078), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(KEYINPUT17), .Z(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2084), .B(G2090), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT84), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n637), .A2(new_n639), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n641), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT85), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n639), .A3(new_n637), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  NAND3_X1  g223(.A1(new_n638), .A2(new_n643), .A3(new_n640), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT86), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1971), .B(G1976), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT19), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1956), .B(G2474), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n655), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  MUX2_X1   g245(.A(G23), .B(G288), .S(G16), .Z(new_n671));
  XOR2_X1   g246(.A(KEYINPUT33), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT91), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G22), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G166), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(G1971), .Z(new_n678));
  NOR2_X1   g253(.A1(G6), .A2(G16), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n569), .B2(G16), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT32), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n674), .A2(new_n678), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  OAI21_X1  g262(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n688));
  INV_X1    g263(.A(G107), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(G2105), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  INV_X1    g266(.A(G119), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n484), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT88), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n487), .A2(G131), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G25), .B(new_n698), .S(G29), .Z(new_n699));
  XOR2_X1   g274(.A(KEYINPUT35), .B(G1991), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT89), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n699), .A2(new_n701), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n675), .A2(G24), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n576), .B2(new_n675), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1986), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g282(.A1(new_n686), .A2(new_n687), .A3(new_n702), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT36), .Z(new_n709));
  NAND2_X1  g284(.A1(G168), .A2(G16), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n710), .B(new_n711), .C1(G16), .C2(G21), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(new_n710), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(G1966), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT97), .Z(new_n715));
  XOR2_X1   g290(.A(KEYINPUT31), .B(G11), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT96), .B(G28), .Z(new_n717));
  OR2_X1    g292(.A1(new_n717), .A2(KEYINPUT30), .ZN(new_n718));
  AOI21_X1  g293(.A(G29), .B1(new_n717), .B2(KEYINPUT30), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n604), .A2(new_n722), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n721), .B(new_n723), .C1(new_n713), .C2(G1966), .ZN(new_n724));
  INV_X1    g299(.A(G1961), .ZN(new_n725));
  NOR2_X1   g300(.A1(G171), .A2(new_n675), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G5), .B2(new_n675), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n715), .B(new_n724), .C1(new_n725), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n722), .A2(G32), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT26), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n733), .A2(new_n734), .B1(G105), .B2(new_n462), .ZN(new_n735));
  INV_X1    g310(.A(G129), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n484), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G141), .B2(new_n487), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n730), .B1(new_n738), .B2(new_n722), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT27), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1996), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n675), .A2(G19), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT92), .Z(new_n743));
  INV_X1    g318(.A(new_n542), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G16), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(G1341), .Z(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  NAND2_X1  g322(.A1(G164), .A2(G29), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G27), .B2(G29), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n722), .A2(G35), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT99), .Z(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G162), .B2(new_n722), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT29), .B(G2090), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n675), .A2(G4), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n586), .B2(new_n675), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G1348), .ZN(new_n758));
  AND4_X1   g333(.A1(new_n741), .A2(new_n750), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n675), .A2(G20), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT23), .Z(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT100), .B(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G160), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT24), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n766), .A2(G34), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n722), .B1(new_n766), .B2(G34), .ZN(new_n768));
  OAI22_X1  g343(.A1(new_n765), .A2(new_n722), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2084), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n727), .A2(new_n725), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n764), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n757), .A2(G1348), .B1(new_n747), .B2(new_n749), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT94), .B(KEYINPUT25), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G139), .B2(new_n487), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n610), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n468), .B2(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G33), .B(new_n781), .S(G29), .Z(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G2072), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n722), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  OR2_X1    g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n788));
  INV_X1    g363(.A(G128), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n484), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G140), .B2(new_n487), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n786), .B1(new_n791), .B2(new_n722), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT93), .B(G2067), .Z(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n783), .A2(new_n784), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n774), .A2(new_n775), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n729), .A2(new_n759), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n709), .A2(new_n798), .ZN(G311));
  INV_X1    g374(.A(G311), .ZN(G150));
  AOI22_X1  g375(.A1(G93), .A2(new_n515), .B1(new_n517), .B2(G55), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n528), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n541), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n744), .B2(new_n803), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n585), .A2(new_n592), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n809));
  AOI21_X1  g384(.A(G860), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n803), .A2(G860), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT37), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(G145));
  XNOR2_X1  g389(.A(new_n698), .B(new_n613), .ZN(new_n815));
  INV_X1    g390(.A(G142), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n470), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT102), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n820));
  INV_X1    g395(.A(G118), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(new_n484), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G130), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n815), .B(new_n825), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n791), .B(new_n502), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n781), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n738), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n826), .A2(KEYINPUT103), .A3(new_n829), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n832), .B(new_n833), .C1(new_n826), .C2(new_n829), .ZN(new_n834));
  XOR2_X1   g409(.A(G160), .B(KEYINPUT101), .Z(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G162), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n604), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n829), .ZN(new_n840));
  INV_X1    g415(.A(new_n826), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n842), .B2(new_n830), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n839), .A2(KEYINPUT40), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT40), .B1(new_n839), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(G395));
  XOR2_X1   g421(.A(new_n595), .B(KEYINPUT104), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n805), .ZN(new_n848));
  XOR2_X1   g423(.A(G299), .B(new_n584), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT105), .B(KEYINPUT41), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(KEYINPUT41), .B2(new_n850), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n847), .A2(new_n805), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n847), .A2(new_n805), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n850), .ZN(new_n859));
  XNOR2_X1  g434(.A(G288), .B(G290), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(G166), .B(new_n569), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n864), .A2(new_n863), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT42), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n856), .A2(new_n859), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n868), .B1(new_n856), .B2(new_n859), .ZN(new_n870));
  OAI21_X1  g445(.A(G868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n803), .A2(new_n578), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(G295));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n872), .ZN(G331));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n875));
  AOI21_X1  g450(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n876));
  NOR2_X1   g451(.A1(G301), .A2(KEYINPUT107), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n805), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n805), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n849), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n854), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n867), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n882), .B2(new_n884), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n875), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n849), .A2(new_n852), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(KEYINPUT41), .B2(new_n849), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n883), .A2(new_n850), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n867), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n895), .A2(KEYINPUT43), .A3(new_n887), .A4(new_n886), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT44), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n888), .B2(new_n889), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n895), .A2(new_n875), .A3(new_n887), .A4(new_n886), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n898), .A2(new_n903), .ZN(G397));
  INV_X1    g479(.A(G8), .ZN(new_n905));
  NOR2_X1   g480(.A1(G166), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT108), .B1(G160), .B2(G40), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n468), .B1(new_n477), .B2(new_n478), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  INV_X1    g485(.A(G40), .ZN(new_n911));
  NOR4_X1   g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n472), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(G1384), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT45), .B1(new_n502), .B2(new_n914), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n913), .A2(KEYINPUT109), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n919));
  INV_X1    g494(.A(new_n472), .ZN(new_n920));
  INV_X1    g495(.A(new_n478), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n610), .B2(G125), .ZN(new_n922));
  OAI211_X1 g497(.A(G40), .B(new_n920), .C1(new_n922), .C2(new_n468), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n910), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n479), .A2(G2105), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(KEYINPUT108), .A3(G40), .A4(new_n920), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n926), .A3(new_n915), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n919), .B1(new_n927), .B2(new_n916), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT110), .B(G1971), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n918), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n918), .A2(new_n928), .A3(KEYINPUT111), .A4(new_n929), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT50), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n502), .B2(new_n914), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n908), .A2(new_n935), .A3(new_n912), .ZN(new_n936));
  INV_X1    g511(.A(G2090), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n502), .A2(new_n914), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n502), .A2(KEYINPUT112), .A3(new_n914), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n934), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(new_n937), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(G8), .B(new_n907), .C1(new_n932), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n924), .A2(new_n926), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n938), .A2(KEYINPUT50), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n502), .A2(KEYINPUT112), .A3(new_n914), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT112), .B1(new_n502), .B2(new_n914), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT50), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n937), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n930), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G8), .ZN(new_n954));
  INV_X1    g529(.A(new_n907), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n940), .A2(new_n924), .A3(new_n926), .A4(new_n941), .ZN(new_n957));
  INV_X1    g532(.A(G1976), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT52), .B1(G288), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n559), .A2(G1976), .A3(new_n561), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n957), .A2(new_n959), .A3(G8), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n569), .A2(new_n682), .ZN(new_n962));
  OAI21_X1  g537(.A(G1981), .B1(new_n565), .B2(new_n568), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n962), .B(new_n963), .C1(KEYINPUT114), .C2(KEYINPUT49), .ZN(new_n964));
  NAND2_X1  g539(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(KEYINPUT114), .A3(KEYINPUT49), .A4(new_n962), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n957), .A2(G8), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n957), .A2(G8), .A3(new_n960), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n970), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT113), .B1(new_n970), .B2(KEYINPUT52), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n945), .A2(new_n956), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT124), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n949), .A2(new_n950), .A3(KEYINPUT50), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n938), .A2(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n924), .A3(new_n926), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n977), .A2(new_n979), .A3(G2084), .ZN(new_n980));
  INV_X1    g555(.A(new_n927), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n949), .B2(new_n950), .ZN(new_n983));
  AOI21_X1  g558(.A(G1966), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(G8), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(G286), .A2(G8), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n986), .B(KEYINPUT120), .Z(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(KEYINPUT51), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n989));
  INV_X1    g564(.A(G1966), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT45), .B1(new_n940), .B2(new_n941), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n927), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n936), .A2(new_n770), .A3(new_n942), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n905), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n987), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT62), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n980), .B2(new_n984), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n988), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n747), .A2(KEYINPUT53), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n991), .A2(new_n927), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT121), .B(G1961), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n936), .B2(new_n942), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT122), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n981), .A2(new_n983), .A3(KEYINPUT53), .A4(new_n747), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT122), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n977), .A2(new_n979), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1005), .B(new_n1006), .C1(new_n1007), .C2(new_n1002), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n918), .A2(new_n928), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(G2078), .ZN(new_n1012));
  AOI21_X1  g587(.A(G301), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n975), .A2(new_n976), .A3(new_n999), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n907), .B1(new_n953), .B2(G8), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n973), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n999), .A2(new_n1016), .A3(new_n945), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT124), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n996), .A2(new_n998), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n988), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT62), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1014), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1023));
  XNOR2_X1  g598(.A(G299), .B(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1956), .B1(new_n948), .B2(new_n951), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n927), .A2(new_n916), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1024), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT116), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1024), .B(new_n1031), .C1(new_n1025), .C2(new_n1028), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n936), .A2(new_n942), .ZN(new_n1033));
  INV_X1    g608(.A(G1348), .ZN(new_n1034));
  INV_X1    g609(.A(new_n957), .ZN(new_n1035));
  INV_X1    g610(.A(G2067), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1033), .A2(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1030), .B(new_n1032), .C1(new_n585), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n948), .A2(new_n951), .ZN(new_n1039));
  INV_X1    g614(.A(G1956), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  XOR2_X1   g616(.A(G299), .B(new_n1023), .Z(new_n1042));
  INV_X1    g617(.A(new_n1028), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1037), .A2(KEYINPUT60), .A3(new_n586), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n1007), .A2(G1348), .B1(G2067), .B2(new_n957), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n585), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1030), .A2(KEYINPUT61), .A3(new_n1032), .A4(new_n1044), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT58), .B(G1341), .Z(new_n1055));
  AND2_X1   g630(.A1(new_n957), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT117), .B(G1996), .Z(new_n1057));
  NOR3_X1   g632(.A1(new_n927), .A2(new_n916), .A3(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n542), .B(new_n1054), .C1(new_n1056), .C2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT59), .B1(new_n1062), .B2(new_n744), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n957), .A2(new_n1055), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(KEYINPUT119), .A3(new_n542), .A4(new_n1054), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1061), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1044), .A2(new_n1029), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1045), .B1(new_n1053), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1000), .B1(new_n923), .B2(KEYINPUT123), .ZN(new_n1076));
  AND4_X1   g651(.A1(new_n915), .A2(new_n1075), .A3(new_n917), .A4(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1003), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1012), .A2(G301), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1074), .B1(new_n1080), .B2(new_n1013), .ZN(new_n1081));
  AOI21_X1  g656(.A(G2078), .B1(new_n918), .B2(new_n928), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1078), .B1(new_n1082), .B2(KEYINPUT53), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1074), .B1(new_n1083), .B2(G171), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1009), .A2(G301), .A3(new_n1012), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1019), .A2(new_n988), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1073), .A2(new_n975), .A3(new_n1081), .A4(new_n1086), .ZN(new_n1087));
  AND4_X1   g662(.A1(new_n958), .A2(new_n968), .A3(new_n559), .A4(new_n561), .ZN(new_n1088));
  INV_X1    g663(.A(new_n962), .ZN(new_n1089));
  OAI211_X1 g664(.A(G8), .B(new_n957), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n945), .B2(new_n973), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n945), .A2(new_n974), .A3(new_n956), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n994), .A2(G168), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n932), .B2(new_n944), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n955), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n973), .A2(new_n1094), .A3(new_n1092), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(new_n945), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1091), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1022), .A2(new_n1087), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n946), .A2(new_n917), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n698), .A2(new_n701), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n791), .B(G2067), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n738), .B(G1996), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n698), .A2(new_n701), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  XOR2_X1   g683(.A(new_n576), .B(G1986), .Z(new_n1109));
  OAI21_X1  g684(.A(new_n1102), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1101), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1105), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1104), .B1(new_n1112), .B2(new_n1102), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1036), .B2(new_n791), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1114), .A2(KEYINPUT125), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(KEYINPUT125), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1102), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1102), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT46), .ZN(new_n1122));
  OR3_X1    g697(.A1(new_n1121), .A2(new_n1122), .A3(G1996), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1105), .A2(new_n738), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1102), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1122), .B1(new_n1121), .B2(G1996), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT47), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1121), .A2(G1986), .A3(G290), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT48), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n1108), .A2(new_n1102), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT127), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(KEYINPUT127), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1128), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1119), .A2(new_n1120), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1111), .A2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g712(.A1(new_n839), .A2(new_n843), .ZN(new_n1139));
  OAI21_X1  g713(.A(G319), .B1(new_n634), .B2(new_n635), .ZN(new_n1140));
  NOR3_X1   g714(.A1(G229), .A2(G227), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g715(.A1(new_n1139), .A2(new_n901), .A3(new_n1141), .ZN(G225));
  INV_X1    g716(.A(G225), .ZN(G308));
endmodule


