//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G104), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n190), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n191), .B1(new_n196), .B2(KEYINPUT77), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n192), .A2(G104), .ZN(new_n199));
  AOI21_X1  g013(.A(G107), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n189), .B1(new_n197), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT76), .B(G104), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT3), .B1(new_n204), .B2(G107), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n194), .A2(KEYINPUT3), .A3(G107), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n204), .B2(G107), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(new_n189), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT78), .B1(new_n203), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT67), .B1(new_n211), .B2(G116), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  INV_X1    g027(.A(G116), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n214), .A2(G119), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G113), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n220), .B2(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT2), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT68), .B1(new_n219), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n217), .B1(new_n212), .B2(new_n215), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n231), .A3(new_n227), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n221), .A2(new_n223), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n200), .A2(new_n201), .B1(G104), .B2(new_n190), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n196), .A2(KEYINPUT77), .ZN(new_n235));
  OAI21_X1  g049(.A(G101), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(new_n208), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n210), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n198), .A2(new_n199), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(new_n241), .B2(new_n190), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n198), .A2(new_n199), .A3(G107), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n190), .A3(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(G101), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(new_n208), .A3(KEYINPUT4), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n219), .A2(new_n228), .ZN(new_n248));
  AND4_X1   g062(.A1(new_n231), .A2(new_n216), .A3(new_n218), .A4(new_n227), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n231), .B1(new_n230), .B2(new_n227), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n189), .B1(new_n205), .B2(new_n207), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n247), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT82), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n247), .A2(new_n251), .A3(new_n254), .A4(KEYINPUT82), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n239), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G110), .B(G122), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n239), .A2(new_n257), .A3(new_n260), .A4(new_n258), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(KEYINPUT6), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n259), .A2(new_n265), .A3(new_n261), .ZN(new_n266));
  OR2_X1    g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  INV_X1    g082(.A(G146), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(G143), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G146), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n267), .B(new_n268), .C1(new_n270), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n271), .B2(G146), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n269), .A2(KEYINPUT65), .A3(G143), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(G146), .ZN(new_n277));
  INV_X1    g091(.A(new_n268), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G125), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT1), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n275), .A2(new_n276), .A3(new_n284), .A4(new_n277), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(KEYINPUT66), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G128), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n269), .A2(G143), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n286), .A2(new_n288), .B1(new_n289), .B2(KEYINPUT1), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n270), .A2(new_n272), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n285), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G125), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n282), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G224), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n294), .B(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n264), .A2(new_n266), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT84), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n264), .A2(new_n300), .A3(new_n266), .A4(new_n297), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G902), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT87), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n223), .A2(new_n305), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n223), .A2(new_n305), .B1(new_n230), .B2(KEYINPUT5), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n306), .A2(new_n307), .B1(new_n229), .B2(new_n232), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n210), .A2(new_n238), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n221), .A2(new_n223), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n249), .B2(new_n250), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n236), .A2(new_n208), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n260), .B(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n304), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  AOI211_X1 g132(.A(KEYINPUT87), .B(new_n316), .C1(new_n309), .C2(new_n313), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT7), .ZN(new_n321));
  INV_X1    g135(.A(new_n296), .ZN(new_n322));
  OAI22_X1  g136(.A1(new_n282), .A2(new_n293), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT88), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT7), .B1(new_n296), .B2(KEYINPUT89), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(KEYINPUT89), .B2(new_n296), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n281), .B(new_n326), .C1(G125), .C2(new_n292), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT90), .ZN(new_n328));
  OR2_X1    g142(.A1(new_n323), .A2(KEYINPUT88), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n263), .A2(new_n324), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n303), .B1(new_n320), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n302), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(G210), .B1(G237), .B2(G902), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n302), .A2(new_n332), .A3(new_n334), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n188), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT66), .B(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G119), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n211), .A2(G128), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT71), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT24), .B(G110), .Z(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT72), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT72), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n343), .A2(new_n349), .A3(new_n345), .A4(new_n346), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT16), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT16), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G125), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n269), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(G125), .ZN(new_n359));
  INV_X1    g173(.A(G125), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(G146), .B(new_n356), .C1(new_n362), .C2(new_n354), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT23), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n365), .B1(new_n211), .B2(G128), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n341), .B(new_n366), .C1(new_n340), .C2(new_n365), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G110), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n351), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n363), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n353), .A2(KEYINPUT73), .A3(G146), .A4(new_n356), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n352), .A2(new_n269), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n367), .A2(G110), .ZN(new_n377));
  INV_X1    g191(.A(new_n346), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n340), .A2(new_n344), .A3(new_n341), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n344), .B1(new_n340), .B2(new_n341), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n376), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT22), .B(G137), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n295), .A2(G221), .A3(G234), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n384), .B(new_n385), .Z(new_n386));
  NAND3_X1  g200(.A1(new_n371), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n369), .B1(new_n348), .B2(new_n350), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n382), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT74), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT25), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n391), .A2(new_n392), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n395), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n387), .A2(new_n390), .A3(new_n397), .A4(new_n393), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(G234), .B2(new_n303), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n387), .A2(new_n390), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n400), .A2(G902), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(G472), .A2(G902), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n273), .A2(new_n279), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT11), .ZN(new_n409));
  INV_X1    g223(.A(G134), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(G137), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(G137), .ZN(new_n412));
  INV_X1    g226(.A(G137), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT11), .A3(G134), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G131), .ZN(new_n416));
  INV_X1    g230(.A(G131), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n411), .A2(new_n414), .A3(new_n417), .A4(new_n412), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n408), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n413), .A2(G134), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n410), .A2(G137), .ZN(new_n422));
  OAI21_X1  g236(.A(G131), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n292), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT64), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT30), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n429));
  AOI211_X1 g243(.A(KEYINPUT64), .B(new_n429), .C1(new_n420), .C2(new_n425), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n251), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT69), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n426), .A2(new_n432), .A3(new_n251), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n419), .A2(new_n408), .B1(new_n424), .B2(new_n292), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n229), .A2(new_n232), .B1(new_n219), .B2(new_n228), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT69), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(G237), .A2(G953), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G210), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(KEYINPUT27), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G101), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n431), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT31), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT31), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n431), .A2(new_n437), .A3(new_n445), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n426), .A2(new_n251), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT28), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT70), .B1(new_n434), .B2(new_n435), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n432), .B1(new_n426), .B2(new_n251), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT69), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT70), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n426), .A2(new_n453), .A3(new_n251), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n450), .A2(new_n451), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n449), .B1(new_n455), .B2(KEYINPUT28), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(new_n442), .ZN(new_n457));
  OAI211_X1 g271(.A(KEYINPUT32), .B(new_n407), .C1(new_n447), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n426), .A2(new_n251), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n449), .B1(new_n460), .B2(KEYINPUT28), .ZN(new_n461));
  INV_X1    g275(.A(new_n442), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n462), .B(new_n449), .C1(new_n455), .C2(KEYINPUT28), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n429), .B1(new_n434), .B2(KEYINPUT64), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n280), .B1(new_n418), .B2(new_n416), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n418), .A2(new_n423), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n289), .A2(KEYINPUT1), .ZN(new_n470));
  OAI22_X1  g284(.A1(new_n470), .A2(new_n339), .B1(new_n270), .B2(new_n272), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n471), .B2(new_n285), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n427), .B(KEYINPUT30), .C1(new_n468), .C2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n435), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n451), .A2(new_n452), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n462), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n465), .B1(new_n466), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G472), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n458), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n444), .B(new_n446), .C1(new_n442), .C2(new_n456), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT32), .B1(new_n481), .B2(new_n407), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n406), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G110), .B(G140), .ZN(new_n485));
  INV_X1    g299(.A(G227), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G953), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n485), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n275), .A2(new_n277), .A3(new_n276), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n489), .B1(new_n470), .B2(new_n283), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n285), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n236), .A2(new_n208), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT10), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n280), .B1(new_n252), .B2(new_n253), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n247), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n471), .B2(new_n285), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n210), .A2(new_n238), .A3(new_n496), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n419), .B(KEYINPUT79), .Z(new_n498));
  AND3_X1   g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n419), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n500), .B1(new_n495), .B2(new_n497), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n488), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT81), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n505));
  INV_X1    g319(.A(new_n488), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n292), .B1(new_n210), .B2(new_n238), .ZN(new_n508));
  INV_X1    g322(.A(new_n492), .ZN(new_n509));
  OAI211_X1 g323(.A(KEYINPUT80), .B(new_n419), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT12), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n500), .A2(KEYINPUT12), .ZN(new_n512));
  OAI211_X1 g326(.A(KEYINPUT80), .B(new_n512), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n507), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(KEYINPUT81), .B(new_n488), .C1(new_n499), .C2(new_n501), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n504), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G469), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n303), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n511), .A2(new_n505), .A3(new_n513), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n488), .B(KEYINPUT75), .Z(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR3_X1    g335(.A1(new_n499), .A2(new_n501), .A3(new_n488), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(G469), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(G469), .A2(G902), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G221), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT9), .B(G234), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n526), .B1(new_n528), .B2(new_n303), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n295), .A2(G952), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(G234), .B2(G237), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n303), .B(new_n295), .C1(G234), .C2(G237), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT21), .B(G898), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n283), .A2(G143), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n339), .B2(G143), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n410), .ZN(new_n540));
  OR2_X1    g354(.A1(KEYINPUT93), .A2(G122), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT93), .A2(G122), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n214), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n214), .A2(G122), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n190), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n547));
  OR3_X1    g361(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT14), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(KEYINPUT14), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n545), .B2(KEYINPUT14), .ZN(new_n550));
  AND4_X1   g364(.A1(new_n544), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n540), .B(new_n546), .C1(new_n190), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n545), .ZN(new_n553));
  OAI21_X1  g367(.A(G107), .B1(new_n543), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n546), .A2(new_n554), .B1(new_n410), .B2(new_n539), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n339), .A2(G143), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n538), .A2(KEYINPUT13), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n538), .A2(KEYINPUT13), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n559), .A2(KEYINPUT94), .A3(G134), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT94), .B1(new_n559), .B2(G134), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n555), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n527), .A2(new_n399), .A3(G953), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n552), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n552), .B2(new_n562), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n303), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G478), .ZN(new_n567));
  NOR2_X1   g381(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT96), .A2(KEYINPUT15), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n303), .B(new_n573), .C1(new_n564), .C2(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n438), .A2(G143), .A3(G214), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(G143), .B1(new_n438), .B2(G214), .ZN(new_n578));
  OAI21_X1  g392(.A(G131), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n438), .A2(G214), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n271), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n417), .A3(new_n576), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(KEYINPUT17), .B(G131), .C1(new_n577), .C2(new_n578), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(new_n358), .A3(new_n363), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n352), .A2(new_n269), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(KEYINPUT91), .B2(new_n375), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n362), .A2(KEYINPUT91), .A3(G146), .ZN(new_n589));
  AND4_X1   g403(.A1(KEYINPUT18), .A2(new_n581), .A3(G131), .A4(new_n576), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n581), .A2(new_n576), .B1(KEYINPUT18), .B2(G131), .ZN(new_n591));
  OAI22_X1  g405(.A1(new_n588), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G113), .B(G122), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(new_n194), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n586), .B2(new_n592), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n303), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(G475), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT20), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n579), .A2(new_n582), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n352), .A2(KEYINPUT19), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n352), .A2(KEYINPUT19), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n269), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n601), .A2(new_n604), .A3(new_n373), .A4(new_n374), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n592), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n594), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n595), .ZN(new_n609));
  NOR2_X1   g423(.A1(G475), .A2(G902), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n600), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n610), .ZN(new_n612));
  AOI211_X1 g426(.A(KEYINPUT20), .B(new_n612), .C1(new_n608), .C2(new_n595), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n599), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT92), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT92), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n616), .B(new_n599), .C1(new_n611), .C2(new_n613), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n537), .B(new_n575), .C1(new_n615), .C2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n338), .A2(new_n484), .A3(new_n532), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT97), .B(G101), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G3));
  INV_X1    g435(.A(G472), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n481), .B2(new_n303), .ZN(new_n623));
  INV_X1    g437(.A(new_n407), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n474), .A2(new_n475), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n445), .B1(new_n625), .B2(new_n442), .ZN(new_n626));
  INV_X1    g440(.A(new_n446), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n457), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n406), .ZN(new_n632));
  OAI21_X1  g446(.A(KEYINPUT98), .B1(new_n531), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n303), .B1(new_n447), .B2(new_n457), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G472), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n481), .A2(new_n407), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n405), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n638), .A2(new_n525), .A3(new_n639), .A4(new_n530), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n537), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT33), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT99), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n643), .A2(KEYINPUT99), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n644), .B(new_n645), .C1(new_n564), .C2(new_n565), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n552), .A2(new_n562), .ZN(new_n647));
  INV_X1    g461(.A(new_n563), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n552), .A2(new_n562), .A3(new_n563), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n649), .A2(KEYINPUT99), .A3(new_n643), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n567), .A2(G902), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n566), .A2(new_n567), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n615), .A2(new_n617), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n338), .A2(new_n642), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n641), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT34), .B(G104), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  AOI21_X1  g477(.A(new_n334), .B1(new_n302), .B2(new_n332), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n335), .B(new_n331), .C1(new_n299), .C2(new_n301), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n187), .B(new_n642), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n575), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n614), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n667), .A2(new_n633), .A3(new_n640), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT35), .B(G107), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  OAI21_X1  g486(.A(KEYINPUT100), .B1(new_n389), .B2(new_n382), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n389), .A2(KEYINPUT100), .A3(new_n382), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n388), .A2(KEYINPUT36), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n675), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n676), .B1(new_n679), .B2(new_n673), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n403), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n401), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n637), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n338), .A2(new_n532), .A3(new_n618), .A4(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT37), .B(G110), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G12));
  OAI21_X1  g502(.A(new_n187), .B1(new_n664), .B2(new_n665), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(new_n531), .ZN(new_n690));
  INV_X1    g504(.A(new_n534), .ZN(new_n691));
  INV_X1    g505(.A(new_n535), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n691), .B1(new_n692), .B2(G900), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT101), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n668), .A2(new_n614), .A3(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n695), .B(new_n683), .C1(new_n480), .C2(new_n482), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  NAND2_X1  g513(.A1(new_n336), .A2(new_n337), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n700), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n694), .B(KEYINPUT39), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n532), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT40), .ZN(new_n706));
  INV_X1    g520(.A(new_n625), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n442), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n460), .A2(new_n442), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n709), .A2(G902), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n622), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n482), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n458), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n658), .A2(new_n668), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NOR4_X1   g530(.A1(new_n714), .A2(new_n716), .A3(new_n188), .A4(new_n683), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT40), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n532), .A2(new_n718), .A3(new_n704), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n703), .A2(new_n706), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  INV_X1    g535(.A(new_n694), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n615), .A2(new_n656), .A3(new_n617), .A4(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n723), .B(new_n683), .C1(new_n480), .C2(new_n482), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n690), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  NAND2_X1  g541(.A1(new_n516), .A2(new_n303), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n530), .A3(new_n518), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n730), .A2(new_n483), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT103), .B1(new_n660), .B2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n667), .A2(new_n734), .A3(new_n659), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NAND3_X1  g552(.A1(new_n667), .A2(new_n669), .A3(new_n731), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G116), .ZN(G18));
  INV_X1    g554(.A(new_n730), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n618), .B(new_n683), .C1(new_n480), .C2(new_n482), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n338), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G119), .ZN(G21));
  AND4_X1   g559(.A1(new_n530), .A2(new_n729), .A3(new_n518), .A4(new_n642), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n405), .A2(KEYINPUT107), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n401), .A2(new_n404), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n474), .A2(new_n475), .A3(new_n462), .ZN(new_n751));
  OAI22_X1  g565(.A1(new_n751), .A2(new_n445), .B1(new_n461), .B2(new_n442), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n627), .B1(new_n752), .B2(KEYINPUT104), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n460), .A2(KEYINPUT28), .ZN(new_n754));
  INV_X1    g568(.A(new_n449), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n756), .A2(new_n462), .B1(new_n443), .B2(KEYINPUT31), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI211_X1 g573(.A(KEYINPUT105), .B(new_n624), .C1(new_n753), .C2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n635), .A2(KEYINPUT106), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n623), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n446), .B1(new_n757), .B2(new_n758), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n752), .A2(KEYINPUT104), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n407), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n762), .A2(new_n764), .B1(new_n767), .B2(KEYINPUT105), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n746), .A2(new_n750), .A3(new_n761), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n700), .A2(new_n187), .A3(new_n715), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(G122), .Z(G24));
  AOI211_X1 g586(.A(KEYINPUT106), .B(new_n622), .C1(new_n481), .C2(new_n303), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n763), .B1(new_n634), .B2(G472), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n624), .B1(new_n753), .B2(new_n759), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT105), .ZN(new_n776));
  OAI22_X1  g590(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n723), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n684), .A4(new_n760), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n689), .A2(new_n730), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G125), .ZN(G27));
  INV_X1    g596(.A(KEYINPUT108), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n525), .B2(new_n530), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n664), .A2(new_n665), .A3(new_n188), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n525), .A2(new_n783), .A3(new_n530), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n785), .A2(new_n786), .A3(new_n484), .A4(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n778), .A2(KEYINPUT42), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n336), .A2(new_n187), .A3(new_n337), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n525), .A2(new_n783), .A3(new_n530), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n784), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n458), .B(new_n479), .C1(new_n482), .C2(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n630), .A2(KEYINPUT109), .A3(KEYINPUT32), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n750), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT110), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n799), .B(new_n750), .C1(new_n795), .C2(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n793), .A2(new_n801), .A3(new_n723), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n790), .B1(new_n802), .B2(KEYINPUT42), .ZN(new_n803));
  XOR2_X1   g617(.A(KEYINPUT111), .B(G131), .Z(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G33));
  INV_X1    g619(.A(new_n695), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n788), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n410), .ZN(G36));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n521), .A2(new_n522), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(G469), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n810), .A2(new_n811), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n814), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n517), .B1(new_n810), .B2(new_n811), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT46), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n820), .B1(G469), .B2(G902), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(KEYINPUT113), .A3(new_n518), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n819), .A2(new_n524), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n820), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n524), .A2(KEYINPUT46), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n827), .B1(new_n815), .B2(new_n818), .ZN(new_n828));
  INV_X1    g642(.A(new_n518), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n704), .A2(new_n530), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n658), .A2(new_n656), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(KEYINPUT43), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT114), .B(KEYINPUT43), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n658), .B2(new_n656), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n631), .B2(new_n684), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n637), .A2(KEYINPUT115), .A3(new_n683), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n786), .B1(new_n845), .B2(KEYINPUT44), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(KEYINPUT44), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT116), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT116), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n845), .A2(new_n850), .A3(KEYINPUT44), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n834), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G137), .ZN(G39));
  NAND2_X1  g668(.A1(new_n831), .A2(new_n530), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT47), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT47), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n831), .A2(new_n857), .A3(new_n530), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n458), .A2(new_n479), .ZN(new_n859));
  INV_X1    g673(.A(new_n482), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n791), .A2(new_n861), .A3(new_n406), .A4(new_n778), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(G140), .ZN(G42));
  NOR2_X1   g678(.A1(new_n841), .A2(new_n691), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n791), .A2(new_n730), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n801), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT48), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n777), .A2(new_n760), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n865), .A2(new_n750), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n533), .B1(new_n870), .B2(new_n780), .ZN(new_n871));
  INV_X1    g685(.A(new_n659), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n866), .A2(new_n406), .A3(new_n534), .A4(new_n714), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n868), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n700), .B(new_n701), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n730), .A2(new_n187), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n870), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT50), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n777), .A2(new_n684), .A3(new_n760), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n866), .A2(new_n879), .A3(new_n865), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT118), .Z(new_n881));
  AOI211_X1 g695(.A(new_n656), .B(new_n873), .C1(new_n615), .C2(new_n617), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n729), .A2(new_n518), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n884), .A2(new_n530), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n856), .B2(new_n858), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n870), .A2(new_n786), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n874), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n889), .B2(new_n888), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n716), .A2(new_n683), .A3(new_n694), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n338), .A2(new_n532), .A3(new_n713), .A4(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n338), .B(new_n532), .C1(new_n725), .C2(new_n697), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n781), .A2(KEYINPUT52), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n781), .A2(new_n894), .A3(new_n893), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT52), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n896), .A3(new_n899), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n658), .A2(new_n656), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n668), .B2(new_n658), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n667), .A2(new_n633), .A3(new_n640), .A4(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n906), .A2(new_n686), .A3(new_n739), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n744), .B1(new_n769), .B2(new_n770), .ZN(new_n908));
  INV_X1    g722(.A(new_n619), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n910), .A3(new_n736), .ZN(new_n911));
  INV_X1    g725(.A(new_n800), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT109), .B1(new_n630), .B2(KEYINPUT32), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n482), .A2(new_n794), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n859), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n799), .B1(new_n915), .B2(new_n750), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n723), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT42), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n788), .A2(new_n789), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n793), .A2(new_n484), .A3(new_n695), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n575), .A2(new_n614), .A3(new_n694), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n683), .B(new_n922), .C1(new_n480), .C2(new_n482), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n791), .A2(new_n531), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n793), .B2(new_n779), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n911), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n903), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n906), .A2(new_n686), .A3(new_n739), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n619), .B(new_n744), .C1(new_n770), .C2(new_n769), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n879), .A2(new_n723), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n531), .A2(new_n923), .ZN(new_n933));
  OAI22_X1  g747(.A1(new_n932), .A2(new_n918), .B1(new_n791), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n934), .A2(new_n807), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n931), .A2(new_n803), .A3(new_n935), .A4(new_n736), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n900), .A2(new_n895), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT53), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT54), .B1(new_n928), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n903), .A2(new_n927), .A3(KEYINPUT53), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n938), .B1(new_n936), .B2(new_n937), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(KEYINPUT54), .B2(new_n943), .ZN(new_n944));
  OAI22_X1  g758(.A1(new_n891), .A2(new_n944), .B1(G952), .B2(G953), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n835), .A2(new_n188), .A3(new_n529), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n714), .A2(new_n750), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(KEYINPUT49), .B2(new_n884), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n875), .C1(KEYINPUT49), .C2(new_n884), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n945), .A2(new_n949), .ZN(G75));
  AOI21_X1  g764(.A(new_n303), .B1(new_n941), .B2(new_n942), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(G210), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT56), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n264), .A2(new_n266), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n297), .ZN(new_n956));
  XOR2_X1   g770(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT120), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n956), .B(new_n958), .Z(new_n959));
  NAND2_X1  g773(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n295), .A2(G952), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n954), .A2(new_n959), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(G51));
  INV_X1    g779(.A(KEYINPUT54), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n943), .B(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n524), .B(KEYINPUT57), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n516), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n951), .A2(new_n815), .A3(new_n818), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n961), .B1(new_n969), .B2(new_n970), .ZN(G54));
  AND2_X1   g785(.A1(KEYINPUT58), .A2(G475), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n951), .A2(new_n609), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n609), .B1(new_n951), .B2(new_n972), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n974), .A3(new_n961), .ZN(G60));
  XNOR2_X1  g789(.A(new_n652), .B(KEYINPUT121), .ZN(new_n976));
  NAND2_X1  g790(.A1(G478), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT59), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n962), .B1(new_n967), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n976), .B1(new_n944), .B2(new_n978), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(G63));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT60), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n943), .A2(new_n681), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT61), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n985), .B1(new_n941), .B2(new_n942), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n962), .B1(new_n989), .B2(new_n402), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n983), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT61), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n989), .B2(new_n681), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n943), .A2(new_n986), .ZN(new_n994));
  INV_X1    g808(.A(new_n402), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n993), .A2(new_n996), .A3(KEYINPUT123), .A4(new_n962), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n991), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT122), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n987), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n989), .A2(KEYINPUT122), .A3(new_n681), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1000), .A2(new_n996), .A3(new_n962), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n992), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n998), .A2(new_n1003), .ZN(G66));
  INV_X1    g818(.A(G224), .ZN(new_n1005));
  OAI21_X1  g819(.A(G953), .B1(new_n536), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n911), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1006), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n955), .B1(G898), .B2(new_n295), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(G69));
  INV_X1    g824(.A(KEYINPUT124), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n921), .A2(new_n781), .A3(new_n894), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n770), .B1(new_n800), .B2(new_n798), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n846), .B1(KEYINPUT116), .B2(new_n848), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1013), .B1(new_n1014), .B2(new_n851), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n831), .A2(new_n833), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n803), .B(new_n1012), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  AND3_X1   g831(.A1(new_n831), .A2(new_n857), .A3(new_n530), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n857), .B1(new_n831), .B2(new_n530), .ZN(new_n1019));
  INV_X1    g833(.A(new_n862), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1011), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n834), .B1(new_n852), .B2(new_n1013), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1012), .A2(new_n803), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n863), .A2(new_n1023), .A3(new_n1024), .A4(KEYINPUT124), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1022), .A2(new_n295), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n428), .A2(new_n430), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n602), .A2(new_n603), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1027), .B(new_n1028), .Z(new_n1029));
  AOI21_X1  g843(.A(new_n1029), .B1(G900), .B2(G953), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n720), .A2(new_n781), .A3(new_n894), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT62), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n720), .A2(KEYINPUT62), .A3(new_n781), .A4(new_n894), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n484), .A2(new_n905), .ZN(new_n1037));
  NOR3_X1   g851(.A1(new_n705), .A2(new_n1037), .A3(new_n791), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1038), .B1(new_n834), .B2(new_n852), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n863), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1029), .B1(new_n1040), .B2(G953), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1031), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(G900), .ZN(new_n1043));
  OAI21_X1  g857(.A(G953), .B1(new_n486), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT125), .Z(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1031), .A2(new_n1041), .A3(new_n1045), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1047), .A2(new_n1048), .ZN(G72));
  NAND4_X1  g863(.A1(new_n863), .A2(new_n1039), .A3(new_n1036), .A4(new_n1007), .ZN(new_n1050));
  NAND2_X1  g864(.A1(G472), .A2(G902), .ZN(new_n1051));
  XOR2_X1   g865(.A(new_n1051), .B(KEYINPUT63), .Z(new_n1052));
  NAND2_X1  g866(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g867(.A(new_n708), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n707), .A2(new_n442), .ZN(new_n1056));
  INV_X1    g870(.A(new_n1056), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n1057), .A2(new_n708), .A3(new_n1052), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1058), .B1(new_n928), .B2(new_n939), .ZN(new_n1059));
  AND3_X1   g873(.A1(new_n1055), .A2(new_n962), .A3(new_n1059), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n1022), .A2(new_n1007), .A3(new_n1025), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n1061), .A2(new_n1052), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1062), .A2(new_n1056), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n1060), .A2(new_n1063), .A3(KEYINPUT126), .ZN(new_n1064));
  INV_X1    g878(.A(KEYINPUT126), .ZN(new_n1065));
  NAND3_X1  g879(.A1(new_n1055), .A2(new_n962), .A3(new_n1059), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1057), .B1(new_n1061), .B2(new_n1052), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1064), .A2(new_n1068), .ZN(G57));
endmodule


