//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n212), .B(new_n218), .C1(G116), .C2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(new_n205), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n202), .A2(G50), .ZN(new_n232));
  OAI22_X1  g0032(.A1(new_n227), .A2(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n209), .B(new_n233), .C1(new_n227), .C2(new_n228), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT76), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT14), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G41), .B2(G45), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n256), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n216), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT68), .B(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n264), .A2(new_n215), .B1(new_n236), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n262), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n263), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n258), .B1(new_n211), .B2(new_n261), .C1(new_n271), .C2(new_n260), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n273));
  XOR2_X1   g0073(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n254), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n272), .B(new_n273), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n277), .B(G169), .C1(new_n252), .C2(new_n253), .ZN(new_n278));
  INV_X1    g0078(.A(G179), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n272), .A2(KEYINPUT13), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n280), .B1(new_n273), .B2(new_n272), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n276), .B(new_n278), .C1(new_n279), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n229), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n262), .A2(G20), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT70), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G77), .B1(G20), .B2(new_n210), .ZN(new_n288));
  INV_X1    g0088(.A(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n262), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n285), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT11), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n255), .A2(new_n210), .A3(G13), .A4(G20), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(KEYINPUT11), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n255), .A2(G20), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n285), .A2(G68), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n294), .A2(new_n296), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT77), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n282), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n274), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G190), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n281), .A2(new_n305), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n304), .A2(new_n306), .A3(new_n300), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g0109(.A(KEYINPUT8), .B(G58), .Z(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT69), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n287), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n291), .A2(G150), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n289), .B1(new_n201), .B2(new_n214), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n255), .A2(G13), .A3(G20), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n316), .A2(new_n284), .B1(new_n214), .B2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n284), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n320), .A2(KEYINPUT72), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(KEYINPUT72), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(new_n298), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(new_n214), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G223), .ZN(new_n328));
  INV_X1    g0128(.A(G222), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n270), .B1(new_n328), .B2(new_n265), .C1(new_n264), .C2(new_n329), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(new_n259), .C1(G77), .C2(new_n270), .ZN(new_n331));
  INV_X1    g0131(.A(new_n261), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G226), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n258), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G190), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n319), .A2(KEYINPUT9), .A3(new_n324), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n334), .A2(G200), .B1(new_n338), .B2(KEYINPUT10), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n327), .A2(new_n336), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n338), .A2(KEYINPUT10), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(new_n337), .A2(new_n339), .ZN(new_n343));
  INV_X1    g0143(.A(new_n341), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(new_n336), .A4(new_n327), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n334), .A2(new_n275), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n335), .A2(new_n279), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n325), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n270), .B1(new_n211), .B2(new_n265), .C1(new_n264), .C2(new_n236), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n259), .C1(G107), .C2(new_n270), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n332), .A2(G244), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n258), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT73), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT73), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n350), .A2(new_n354), .A3(new_n258), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G190), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(G200), .A3(new_n355), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT15), .B(G87), .Z(new_n359));
  AOI22_X1  g0159(.A1(new_n310), .A2(new_n291), .B1(new_n359), .B2(new_n286), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n289), .B2(new_n220), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n284), .B1(new_n220), .B2(new_n318), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n285), .A2(G77), .A3(new_n298), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n357), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n342), .A2(new_n345), .A3(new_n348), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G58), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n210), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n201), .ZN(new_n370));
  INV_X1    g0170(.A(G159), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(new_n290), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n267), .A2(KEYINPUT78), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT78), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n375), .A3(G33), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(new_n289), .A3(new_n268), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n210), .B1(new_n377), .B2(KEYINPUT7), .ZN(new_n378));
  NOR2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT7), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n289), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n372), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n285), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n374), .A2(KEYINPUT3), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n267), .A2(KEYINPUT78), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n262), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n389), .A2(KEYINPUT7), .A3(new_n289), .A4(new_n269), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n382), .B1(new_n270), .B2(G20), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n210), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n386), .B1(new_n392), .B2(new_n372), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n311), .A2(new_n318), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n323), .A2(new_n311), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n385), .A2(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n332), .A2(G232), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n264), .A2(new_n328), .B1(new_n215), .B2(new_n265), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n376), .A2(new_n268), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n398), .A2(new_n399), .B1(G33), .B2(G87), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n397), .B(new_n258), .C1(new_n400), .C2(new_n260), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n401), .A2(new_n305), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(G200), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n396), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n396), .A2(KEYINPUT17), .A3(new_n402), .A4(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n385), .A2(new_n393), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n395), .A2(new_n394), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n401), .A2(new_n279), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n401), .A2(G169), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT18), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT18), .B1(new_n410), .B2(new_n413), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n406), .B(new_n407), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n353), .A2(new_n275), .A3(new_n355), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n364), .ZN(new_n419));
  AOI21_X1  g0219(.A(G179), .B1(new_n353), .B2(new_n355), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NOR4_X1   g0221(.A1(new_n309), .A2(new_n367), .A3(new_n417), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT80), .ZN(new_n423));
  INV_X1    g0223(.A(G41), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT5), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT5), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(KEYINPUT80), .B2(G41), .ZN(new_n427));
  INV_X1    g0227(.A(G45), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(G1), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n257), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n260), .A2(new_n430), .A3(G270), .ZN(new_n433));
  INV_X1    g0233(.A(new_n269), .ZN(new_n434));
  INV_X1    g0234(.A(G303), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n434), .A2(new_n379), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G264), .A2(G1698), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n264), .B2(new_n217), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n438), .B2(new_n399), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n432), .B(new_n433), .C1(new_n439), .C2(new_n260), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT84), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT68), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1698), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n445));
  OAI21_X1  g0245(.A(G257), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI22_X1  g0246(.A1(new_n446), .A2(new_n437), .B1(new_n376), .B2(new_n268), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n259), .B1(new_n447), .B2(new_n436), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(KEYINPUT84), .A3(new_n432), .A4(new_n433), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n442), .A2(G200), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n289), .C1(G33), .C2(new_n216), .ZN(new_n452));
  INV_X1    g0252(.A(G116), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G20), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n284), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n452), .A2(KEYINPUT20), .A3(new_n284), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n255), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n317), .A2(new_n459), .A3(new_n229), .A4(new_n283), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n457), .A2(new_n458), .B1(G116), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n318), .A2(new_n453), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n450), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n442), .A2(new_n449), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G190), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n450), .A2(KEYINPUT87), .A3(new_n465), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n275), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n442), .A2(new_n449), .A3(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n440), .A2(new_n279), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n464), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n442), .A2(new_n449), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(KEYINPUT85), .A3(KEYINPUT21), .A4(new_n473), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n442), .A2(new_n449), .A3(KEYINPUT21), .A4(new_n473), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT85), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n472), .A2(new_n477), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n260), .A2(new_n430), .A3(G264), .ZN(new_n485));
  XNOR2_X1  g0285(.A(new_n485), .B(KEYINPUT91), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n399), .A2(G257), .A3(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT90), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G294), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT90), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n399), .A2(new_n490), .A3(G257), .A4(G1698), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n399), .B(G250), .C1(new_n444), .C2(new_n445), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n488), .A2(new_n489), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n486), .B1(new_n493), .B2(new_n259), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(G179), .A3(new_n432), .ZN(new_n495));
  AOI211_X1 g0295(.A(new_n431), .B(new_n486), .C1(new_n493), .C2(new_n259), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n275), .ZN(new_n497));
  INV_X1    g0297(.A(G87), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n498), .A2(G20), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n399), .A2(KEYINPUT22), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n434), .B2(new_n379), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT22), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n289), .B2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT23), .A3(G20), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n501), .A2(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n286), .A2(G116), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n500), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT24), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n500), .A2(new_n507), .A3(new_n511), .A4(new_n508), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n285), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n460), .A2(new_n505), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT88), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(KEYINPUT25), .ZN(new_n517));
  NOR3_X1   g0317(.A1(new_n317), .A2(new_n517), .A3(G107), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(KEYINPUT25), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT89), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT89), .ZN(new_n523));
  NOR4_X1   g0323(.A1(new_n513), .A2(new_n523), .A3(new_n514), .A4(new_n520), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n497), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n484), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n260), .A2(new_n430), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G257), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n264), .A2(new_n221), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT4), .B1(new_n399), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n270), .ZN(new_n532));
  OAI211_X1 g0332(.A(KEYINPUT4), .B(G244), .C1(new_n444), .C2(new_n445), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G250), .A2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n451), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n531), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n432), .B(new_n529), .C1(new_n537), .C2(new_n260), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n533), .A2(new_n534), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n270), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  OAI21_X1  g0342(.A(G244), .B1(new_n444), .B2(new_n445), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n381), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n541), .A2(new_n544), .A3(new_n451), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n259), .B1(G257), .B2(new_n528), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(G190), .A3(new_n432), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n317), .A2(new_n216), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n461), .B2(new_n216), .ZN(new_n549));
  XNOR2_X1  g0349(.A(new_n549), .B(KEYINPUT79), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n216), .A2(new_n505), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n289), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n290), .A2(new_n220), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  AND2_X1   g0359(.A1(new_n390), .A2(new_n391), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n559), .C1(new_n560), .C2(new_n505), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n550), .B1(new_n561), .B2(new_n284), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n539), .A2(new_n547), .A3(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT79), .ZN(new_n564));
  XNOR2_X1  g0364(.A(new_n549), .B(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n505), .B1(new_n390), .B2(new_n391), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n566), .A2(new_n558), .A3(new_n556), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n567), .B2(new_n285), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n545), .A2(new_n259), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(new_n279), .A3(new_n432), .A4(new_n529), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(G169), .B1(new_n546), .B2(new_n432), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT81), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n538), .A2(new_n275), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT81), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n570), .A4(new_n568), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n563), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n399), .A2(new_n289), .A3(G68), .ZN(new_n579));
  NOR3_X1   g0379(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(G33), .B2(G97), .ZN(new_n581));
  OAI21_X1  g0381(.A(KEYINPUT19), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT19), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n263), .A2(new_n583), .A3(new_n289), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n285), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n359), .A2(new_n317), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n578), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n587), .ZN(new_n589));
  AOI21_X1  g0389(.A(G20), .B1(new_n376), .B2(new_n268), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(G68), .B1(new_n582), .B2(new_n584), .ZN(new_n591));
  OAI211_X1 g0391(.A(KEYINPUT82), .B(new_n589), .C1(new_n591), .C2(new_n285), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n429), .A2(G274), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n260), .B(G250), .C1(G1), .C2(new_n428), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n264), .A2(new_n211), .B1(new_n221), .B2(new_n265), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n399), .B1(G33), .B2(G116), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n594), .B(new_n595), .C1(new_n597), .C2(new_n260), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G190), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n461), .A2(G87), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n598), .A2(G200), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n593), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n359), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n460), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NOR3_X1   g0406(.A1(new_n586), .A2(new_n578), .A3(new_n587), .ZN(new_n607));
  AOI211_X1 g0407(.A(G20), .B(new_n210), .C1(new_n376), .C2(new_n268), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n582), .A2(new_n584), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n284), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT82), .B1(new_n610), .B2(new_n589), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n607), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT83), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT83), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n593), .A2(new_n614), .A3(new_n606), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n598), .A2(G179), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n275), .B2(new_n598), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n603), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n494), .A2(new_n432), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G200), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n513), .A2(new_n514), .A3(new_n520), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n305), .C2(new_n620), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n577), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n422), .A2(new_n527), .A3(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n420), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n364), .A3(new_n418), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n302), .B1(new_n307), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n406), .A2(new_n407), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n416), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n414), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n342), .A2(new_n345), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n348), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n422), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT93), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n571), .B2(new_n572), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n574), .A2(KEYINPUT93), .A3(new_n570), .A4(new_n568), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n619), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n614), .B1(new_n593), .B2(new_n606), .ZN(new_n646));
  AOI211_X1 g0446(.A(KEYINPUT83), .B(new_n605), .C1(new_n588), .C2(new_n592), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n618), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n593), .A2(new_n601), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(new_n600), .A3(new_n602), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n648), .A2(new_n573), .A3(new_n651), .A4(new_n576), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n515), .A2(new_n521), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n497), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n480), .A2(new_n481), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n480), .A2(new_n481), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n477), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT92), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n477), .B(KEYINPUT92), .C1(new_n656), .C2(new_n657), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n655), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n577), .A2(new_n619), .A3(new_n623), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n645), .B(new_n653), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n638), .B1(new_n639), .B2(new_n665), .ZN(G369));
  INV_X1    g0466(.A(G13), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(G20), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n255), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n525), .A2(new_n623), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n676), .A2(new_n658), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n677), .B2(new_n655), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n465), .A2(new_n675), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n660), .A2(new_n661), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n679), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n472), .A2(new_n477), .A3(new_n483), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n526), .A2(new_n674), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n674), .B1(new_n522), .B2(new_n524), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n525), .A2(new_n685), .A3(new_n623), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(G330), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n678), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n206), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n580), .A2(new_n453), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n232), .B2(new_n692), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n525), .A2(new_n477), .A3(new_n483), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n619), .A3(new_n577), .A4(new_n623), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n648), .A2(new_n573), .A3(new_n651), .A4(new_n576), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n649), .B1(new_n700), .B2(new_n644), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n643), .A2(new_n619), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT26), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n675), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n664), .A2(new_n707), .A3(new_n675), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n624), .A2(new_n527), .A3(new_n675), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n442), .A2(new_n449), .A3(new_n598), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n620), .A2(new_n710), .A3(new_n279), .A4(new_n538), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n494), .A2(new_n476), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n546), .A2(new_n432), .A3(new_n599), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n712), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT94), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n711), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n713), .A2(new_n714), .A3(new_n712), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT31), .B(new_n674), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n674), .B1(new_n716), .B2(new_n721), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n709), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n706), .A2(new_n708), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n697), .B1(new_n729), .B2(G1), .ZN(G364));
  NOR2_X1   g0530(.A1(new_n532), .A2(new_n690), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G355), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n250), .A2(new_n428), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n399), .A2(new_n690), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G45), .B2(new_n232), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n732), .B1(G116), .B2(new_n206), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n229), .B1(G20), .B2(new_n275), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n255), .B1(new_n668), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n691), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n289), .A2(new_n305), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n279), .A2(new_n303), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n303), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n749), .A2(new_n214), .B1(new_n751), .B2(new_n498), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n279), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n289), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n270), .B1(new_n754), .B2(new_n368), .C1(new_n210), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n750), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n752), .B(new_n757), .C1(G107), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n755), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(new_n764), .B2(G159), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n763), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n289), .B1(new_n762), .B2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n216), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n755), .A2(new_n753), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n760), .B(new_n769), .C1(new_n220), .C2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n532), .B1(new_n763), .B2(new_n772), .C1(new_n773), .C2(new_n754), .ZN(new_n774));
  INV_X1    g0574(.A(new_n767), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G294), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n749), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G326), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n759), .A2(G283), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n751), .A2(new_n435), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n756), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT33), .B(G317), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n771), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n746), .B1(new_n786), .B2(new_n740), .ZN(new_n787));
  INV_X1    g0587(.A(new_n739), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n742), .B(new_n787), .C1(new_n683), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n683), .A2(G330), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n746), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n683), .A2(G330), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n791), .B2(new_n792), .ZN(G396));
  NOR2_X1   g0593(.A1(new_n758), .A2(new_n498), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n505), .A2(new_n751), .B1(new_n754), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(G311), .C2(new_n764), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n532), .B1(new_n749), .B2(new_n435), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n768), .B(new_n798), .C1(G283), .C2(new_n782), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n797), .B(new_n799), .C1(new_n453), .C2(new_n770), .ZN(new_n800));
  INV_X1    g0600(.A(new_n754), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G143), .A2(new_n801), .B1(new_n782), .B2(G150), .ZN(new_n802));
  INV_X1    g0602(.A(G137), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n803), .B2(new_n749), .C1(new_n371), .C2(new_n770), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT34), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n751), .A2(new_n214), .B1(new_n763), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n381), .B(new_n809), .C1(G58), .C2(new_n775), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n758), .A2(new_n210), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n800), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n746), .B1(new_n813), .B2(new_n740), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n740), .A2(new_n737), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n364), .A2(new_n674), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n421), .B1(new_n366), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n627), .A2(new_n674), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT95), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT95), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n421), .A2(new_n675), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n366), .A2(new_n817), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n421), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n814), .B1(G77), .B2(new_n816), .C1(new_n825), .C2(new_n738), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT96), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n652), .A2(KEYINPUT26), .ZN(new_n828));
  AND3_X1   g0628(.A1(new_n645), .A2(new_n828), .A3(new_n648), .ZN(new_n829));
  INV_X1    g0629(.A(new_n655), .ZN(new_n830));
  INV_X1    g0630(.A(new_n661), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT92), .B1(new_n483), .B2(new_n477), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n624), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n674), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT97), .B1(new_n835), .B2(new_n825), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n664), .A2(KEYINPUT97), .A3(new_n675), .A4(new_n825), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n836), .A2(new_n838), .B1(new_n835), .B2(new_n825), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(new_n727), .Z(new_n840));
  AOI21_X1  g0640(.A(new_n827), .B1(new_n840), .B2(new_n746), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G384));
  AND2_X1   g0642(.A1(new_n554), .A2(new_n555), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT35), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n231), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n845), .B(G116), .C1(new_n844), .C2(new_n843), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT36), .ZN(new_n847));
  OAI21_X1  g0647(.A(G77), .B1(new_n368), .B2(new_n210), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n232), .A2(new_n848), .B1(G50), .B2(new_n210), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(G1), .A3(new_n667), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n822), .B1(new_n836), .B2(new_n838), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT98), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n301), .A2(new_n674), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n302), .A2(new_n308), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n301), .B(new_n674), .C1(new_n282), .C2(new_n307), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n662), .A2(new_n663), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n653), .A2(new_n645), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n675), .B(new_n825), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT97), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n819), .B1(new_n862), .B2(new_n837), .ZN(new_n863));
  INV_X1    g0663(.A(new_n856), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT98), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n672), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n410), .B1(new_n413), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n404), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n385), .B1(KEYINPUT16), .B2(new_n384), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n409), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n413), .B2(new_n866), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n868), .B1(new_n873), .B2(new_n404), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n417), .A2(new_n866), .A3(new_n872), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n872), .A2(new_n866), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n629), .B2(new_n632), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n870), .A2(new_n874), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n857), .A2(new_n865), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n632), .A2(new_n866), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n396), .A2(new_n672), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n867), .A2(new_n404), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT37), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n417), .A2(new_n888), .B1(new_n890), .B2(new_n869), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT99), .B1(new_n891), .B2(KEYINPUT38), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT99), .ZN(new_n893));
  INV_X1    g0693(.A(new_n888), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(new_n629), .B2(new_n632), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n868), .B1(new_n867), .B2(new_n404), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n870), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n893), .B(new_n878), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n892), .A2(new_n898), .A3(new_n877), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n887), .B1(new_n886), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n282), .A2(new_n301), .A3(new_n675), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n885), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n884), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT100), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n706), .A2(new_n708), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n422), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n664), .A2(new_n707), .A3(new_n675), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n707), .B1(new_n704), .B2(new_n675), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n905), .B(new_n422), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n638), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n904), .B(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n854), .A2(new_n855), .B1(new_n824), .B2(new_n820), .ZN(new_n914));
  NOR2_X1   g0714(.A1(KEYINPUT101), .A2(KEYINPUT31), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n723), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n723), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n709), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n883), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n918), .A4(new_n914), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND3_X1   g0723(.A1(new_n709), .A2(new_n916), .A3(new_n917), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n639), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n923), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(G330), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n913), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT102), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT102), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n929), .B(new_n930), .C1(new_n913), .C2(new_n927), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n668), .A2(new_n255), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n847), .B(new_n850), .C1(new_n931), .C2(new_n932), .ZN(G367));
  NAND2_X1  g0733(.A1(new_n573), .A2(new_n576), .ZN(new_n934));
  INV_X1    g0734(.A(new_n563), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n568), .A2(new_n674), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(KEYINPUT104), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n574), .A2(new_n570), .A3(new_n568), .A4(new_n674), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT104), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n577), .A2(new_n940), .A3(new_n936), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(new_n688), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n675), .A3(new_n677), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT42), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n942), .A2(new_n526), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n674), .B1(new_n947), .B2(new_n934), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT43), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n650), .A2(new_n675), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT103), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(new_n619), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n649), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n950), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n950), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n946), .C2(new_n948), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n944), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n958), .A2(new_n944), .A3(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT105), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n691), .B(KEYINPUT41), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n658), .A2(new_n675), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n683), .A2(G330), .A3(new_n687), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n687), .B1(new_n683), .B2(G330), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n687), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n790), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(new_n688), .A3(new_n970), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT108), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n908), .A2(new_n909), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n727), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n676), .A2(new_n658), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n674), .B1(new_n982), .B2(new_n830), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n938), .A2(new_n941), .ZN(new_n984));
  XOR2_X1   g0784(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n985));
  NAND3_X1  g0785(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n985), .B1(new_n983), .B2(new_n984), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n972), .A2(KEYINPUT107), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n943), .B2(new_n983), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n990), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n981), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n990), .ZN(new_n997));
  INV_X1    g0797(.A(new_n994), .ZN(new_n998));
  INV_X1    g0798(.A(new_n988), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n986), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n997), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n974), .A2(new_n977), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT108), .B1(new_n1002), .B2(new_n728), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n996), .A2(KEYINPUT109), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1003), .A2(new_n1001), .A3(new_n981), .A4(new_n995), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n969), .B1(new_n1008), .B2(new_n729), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n967), .B1(new_n1009), .B2(new_n744), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n734), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n741), .B1(new_n206), .B2(new_n604), .C1(new_n1011), .C2(new_n242), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n749), .A2(new_n780), .B1(new_n754), .B2(new_n435), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n751), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT46), .B1(new_n1014), .B2(G116), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n770), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1013), .B(new_n1016), .C1(G283), .C2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n381), .B1(new_n795), .B2(new_n756), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1014), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n505), .B2(new_n767), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1019), .B(new_n1021), .C1(G317), .C2(new_n764), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n759), .A2(G97), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1018), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n758), .A2(new_n220), .ZN(new_n1026));
  INV_X1    g0826(.A(G143), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n749), .A2(new_n1027), .B1(new_n763), .B2(new_n803), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(G150), .C2(new_n801), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n270), .B1(new_n770), .B2(new_n214), .C1(new_n368), .C2(new_n751), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G68), .B2(new_n775), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(new_n371), .C2(new_n756), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT47), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n746), .B1(new_n1034), .B2(new_n740), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1012), .B(new_n1035), .C1(new_n956), .C2(new_n788), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1010), .A2(new_n1036), .ZN(G387));
  NAND2_X1  g0837(.A1(new_n729), .A2(new_n978), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1002), .A2(new_n728), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n691), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G311), .A2(new_n782), .B1(new_n801), .B2(G317), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n435), .B2(new_n770), .C1(new_n773), .C2(new_n749), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT48), .ZN(new_n1043));
  INV_X1    g0843(.A(G283), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n767), .C1(new_n795), .C2(new_n751), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT49), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n399), .B1(G326), .B2(new_n764), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1047), .B(new_n1050), .C1(G116), .C2(new_n759), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n381), .B1(G77), .B2(new_n1014), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT112), .B(G150), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1023), .C1(new_n763), .C2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(KEYINPUT113), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(KEYINPUT113), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n749), .A2(new_n371), .B1(new_n754), .B2(new_n214), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n604), .A2(new_n767), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n311), .C2(new_n782), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1056), .B(new_n1061), .C1(G68), .C2(new_n1017), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n740), .B1(new_n1051), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1011), .B1(new_n239), .B2(G45), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n693), .B2(new_n731), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n310), .A2(new_n214), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT50), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT50), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n428), .A4(new_n694), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G68), .B2(G77), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1065), .A2(new_n1070), .B1(G107), .B2(new_n206), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n746), .B1(new_n1071), .B2(new_n741), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT111), .Z(new_n1073));
  OAI211_X1 g0873(.A(new_n1063), .B(new_n1073), .C1(new_n687), .C2(new_n788), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1040), .B(new_n1074), .C1(new_n743), .C2(new_n1002), .ZN(G393));
  NAND2_X1  g0875(.A1(new_n989), .A2(new_n994), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(new_n688), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n744), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n741), .B1(new_n216), .B2(new_n206), .C1(new_n247), .C2(new_n1011), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G150), .A2(new_n777), .B1(new_n801), .B2(G159), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n756), .A2(new_n214), .B1(new_n763), .B2(new_n1027), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1017), .A2(new_n310), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n399), .B1(new_n210), .B2(new_n751), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n767), .A2(new_n220), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1086), .A2(new_n794), .A3(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1082), .A2(new_n1084), .A3(new_n1085), .A4(new_n1088), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G317), .A2(new_n777), .B1(new_n801), .B2(G311), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT52), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n751), .A2(new_n1044), .B1(new_n763), .B2(new_n773), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT115), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1092), .A2(new_n1093), .B1(G107), .B2(new_n759), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n532), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n770), .A2(new_n795), .B1(new_n767), .B2(new_n453), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G303), .B2(new_n782), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT116), .Z(new_n1099));
  OAI21_X1  g0899(.A(new_n1089), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n746), .B1(new_n1100), .B2(new_n740), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1079), .B(new_n1101), .C1(new_n942), .C2(new_n788), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1078), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1077), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1004), .A2(new_n1007), .B1(new_n1104), .B2(new_n1038), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n1105), .B2(new_n691), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G390));
  OAI21_X1  g0907(.A(new_n901), .B1(new_n863), .B2(new_n864), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n900), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n899), .A2(new_n901), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n704), .A2(new_n675), .A3(new_n825), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n822), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1111), .B1(new_n856), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(G330), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n820), .B2(new_n824), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n726), .A2(new_n856), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1110), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1114), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1117), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n924), .A2(new_n864), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n925), .A2(G330), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n638), .B(new_n1125), .C1(new_n907), .C2(new_n911), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT117), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n856), .B1(new_n918), .B2(new_n1117), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1113), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1129), .B2(new_n1118), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1112), .A2(new_n822), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n864), .B1(new_n924), .B2(new_n1122), .ZN(new_n1132));
  AND4_X1   g0932(.A1(new_n1127), .A2(new_n1131), .A3(new_n1132), .A4(new_n1118), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n856), .B1(new_n726), .B2(new_n1117), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n851), .B1(new_n1123), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1126), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n692), .B1(new_n1124), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1124), .B2(new_n1137), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1124), .A2(new_n744), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n311), .A2(new_n816), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1054), .A2(new_n751), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT53), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT54), .B(G143), .Z(new_n1144));
  AOI22_X1  g0944(.A1(new_n1017), .A2(new_n1144), .B1(new_n759), .B2(G50), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n270), .B1(new_n756), .B2(new_n803), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G128), .B2(new_n777), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n808), .B2(new_n754), .C1(new_n371), .C2(new_n767), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1146), .B(new_n1149), .C1(G125), .C2(new_n764), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(G116), .A2(new_n801), .B1(new_n1017), .B2(G97), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n505), .B2(new_n756), .C1(new_n1044), .C2(new_n749), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n532), .B1(new_n763), .B2(new_n795), .C1(new_n498), .C2(new_n751), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1152), .A2(new_n812), .A3(new_n1087), .A4(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n740), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n745), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1141), .B(new_n1156), .C1(new_n1109), .C2(new_n737), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1139), .A2(new_n1140), .A3(new_n1158), .ZN(G378));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT120), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n904), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT55), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n635), .A2(new_n1165), .A3(new_n348), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n348), .ZN(new_n1167));
  OAI21_X1  g0967(.A(KEYINPUT55), .B1(new_n634), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n325), .A2(new_n866), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1166), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1169), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1164), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1172), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n1163), .A3(new_n1170), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n921), .A2(G330), .A3(new_n922), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1176), .B(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1162), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1177), .B(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n904), .A2(new_n1161), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1126), .B1(new_n1124), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1160), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1114), .B(new_n1118), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1137), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1126), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n904), .A2(new_n1178), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1181), .A2(new_n903), .A3(new_n884), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1160), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n692), .B1(new_n1191), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1186), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT121), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1179), .A2(new_n744), .A3(new_n1182), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1176), .A2(new_n737), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n815), .A2(new_n214), .ZN(new_n1200));
  INV_X1    g1000(.A(G128), .ZN(new_n1201));
  INV_X1    g1001(.A(G150), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n754), .A2(new_n1201), .B1(new_n767), .B2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1014), .A2(new_n1144), .B1(new_n1017), .B2(G137), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n808), .B2(new_n756), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(G125), .C2(new_n777), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT59), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G41), .B1(new_n764), .B2(G124), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G33), .B1(new_n759), .B2(G159), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n381), .B1(new_n210), .B2(new_n767), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n424), .B1(new_n220), .B2(new_n751), .C1(new_n604), .C2(new_n770), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(G116), .C2(new_n777), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n758), .A2(new_n368), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT118), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n756), .A2(new_n216), .B1(new_n763), .B2(new_n1044), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1213), .B(new_n1217), .C1(new_n505), .C2(new_n754), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1218), .B(KEYINPUT58), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G41), .B1(new_n380), .B2(G33), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1210), .B(new_n1219), .C1(G50), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n746), .B1(new_n1221), .B2(new_n740), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1199), .A2(new_n1200), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1197), .B1(new_n1198), .B2(new_n1223), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1198), .A2(new_n1197), .A3(new_n1223), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1196), .B1(new_n1224), .B2(new_n1225), .ZN(G375));
  OAI22_X1  g1026(.A1(new_n754), .A2(new_n803), .B1(new_n763), .B2(new_n1201), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1227), .B(new_n1215), .C1(G150), .C2(new_n1017), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n399), .B1(new_n214), .B2(new_n767), .C1(new_n808), .C2(new_n749), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n782), .B2(new_n1144), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n371), .C2(new_n751), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G97), .A2(new_n1014), .B1(new_n764), .B2(G303), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1044), .B2(new_n754), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1233), .A2(new_n1026), .A3(new_n1059), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n749), .A2(new_n795), .B1(new_n770), .B2(new_n505), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G116), .B2(new_n782), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n270), .B1(new_n1236), .B2(KEYINPUT122), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1234), .B(new_n1237), .C1(KEYINPUT122), .C2(new_n1236), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1231), .A2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n746), .B1(new_n1239), .B2(new_n740), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n856), .B2(new_n738), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n210), .B2(new_n815), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1184), .B2(new_n744), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1134), .A2(new_n1126), .A3(new_n1136), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n968), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1245), .B2(new_n1137), .ZN(G381));
  NOR2_X1   g1046(.A1(G375), .A2(G378), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NOR3_X1   g1048(.A1(new_n1248), .A2(G384), .A3(G381), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1010), .A2(new_n1036), .A3(new_n1106), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(G396), .A3(G393), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(G407));
  OAI211_X1 g1052(.A(G407), .B(G213), .C1(G343), .C2(new_n1248), .ZN(G409));
  OAI211_X1 g1053(.A(new_n1196), .B(G378), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n744), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1191), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1256), .B(new_n1223), .C1(new_n1257), .C2(new_n969), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1139), .A2(new_n1140), .A3(new_n1158), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n673), .A2(G213), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1244), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1244), .A2(new_n1264), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1137), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n691), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1243), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n841), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(G384), .A3(new_n1243), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(G2897), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n1262), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1262), .A2(new_n1273), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1270), .A2(new_n1271), .A3(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1263), .A2(new_n1277), .ZN(new_n1278));
  XOR2_X1   g1078(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1279));
  XOR2_X1   g1079(.A(G393), .B(G396), .Z(new_n1280));
  AND3_X1   g1080(.A1(new_n1010), .A2(new_n1036), .A3(new_n1106), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1106), .B1(new_n1010), .B2(new_n1036), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1280), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(G390), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1280), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1250), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1283), .A2(new_n1286), .A3(KEYINPUT125), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1278), .A2(new_n1279), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT62), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1283), .A2(new_n1286), .A3(KEYINPUT125), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT125), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OR3_X1    g1095(.A1(new_n1287), .A2(KEYINPUT61), .A3(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1272), .ZN(new_n1298));
  AND3_X1   g1098(.A1(new_n1254), .A2(KEYINPUT123), .A3(new_n1260), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT123), .B1(new_n1254), .B2(new_n1260), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1298), .B(new_n1262), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1291), .B1(new_n1297), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1261), .A2(new_n1298), .A3(new_n1262), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT61), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1283), .A2(new_n1286), .A3(new_n1305), .A4(KEYINPUT63), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1262), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1307), .B2(new_n1277), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1292), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1304), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(G405));
  AND3_X1   g1111(.A1(new_n904), .A2(new_n1161), .A3(new_n1181), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1181), .B1(new_n904), .B2(new_n1161), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1312), .A2(new_n1313), .A3(new_n743), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1223), .ZN(new_n1315));
  OAI21_X1  g1115(.A(KEYINPUT121), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1198), .A2(new_n1197), .A3(new_n1223), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1318), .A2(G378), .A3(new_n1196), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G378), .B1(new_n1318), .B2(new_n1196), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1272), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(G375), .A2(new_n1259), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1298), .A3(new_n1254), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(KEYINPUT126), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1321), .A2(new_n1323), .A3(KEYINPUT126), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT126), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1328), .A2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1325), .A2(new_n1331), .A3(new_n1332), .A4(new_n1327), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(G402));
endmodule


