

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778;

  NOR2_X1 U371 ( .A1(n655), .A2(n741), .ZN(n657) );
  XNOR2_X1 U372 ( .A(n355), .B(G119), .ZN(n408) );
  NOR2_X1 U373 ( .A1(n728), .A2(n741), .ZN(n426) );
  AND2_X2 U374 ( .A1(n635), .A2(n364), .ZN(n387) );
  NAND2_X1 U375 ( .A1(n351), .A2(n376), .ZN(n413) );
  NAND2_X1 U376 ( .A1(n375), .A2(KEYINPUT79), .ZN(n351) );
  XNOR2_X2 U377 ( .A(n385), .B(n618), .ZN(n481) );
  BUF_X1 U378 ( .A(G107), .Z(n390) );
  AND2_X1 U379 ( .A1(n510), .A2(G472), .ZN(n352) );
  XNOR2_X2 U380 ( .A(G953), .B(KEYINPUT64), .ZN(n536) );
  AND2_X1 U381 ( .A1(n626), .A2(n472), .ZN(n578) );
  XNOR2_X1 U382 ( .A(n614), .B(n613), .ZN(n619) );
  NOR2_X2 U383 ( .A1(n687), .A2(n637), .ZN(n660) );
  NOR2_X2 U384 ( .A1(n619), .A2(n616), .ZN(n385) );
  XNOR2_X2 U385 ( .A(n631), .B(n406), .ZN(n403) );
  AND2_X2 U386 ( .A1(n402), .A2(n400), .ZN(n394) );
  AND2_X2 U387 ( .A1(n714), .A2(n650), .ZN(n414) );
  XNOR2_X2 U388 ( .A(n745), .B(n465), .ZN(n407) );
  NOR2_X1 U389 ( .A1(n625), .A2(n478), .ZN(n638) );
  INV_X1 U390 ( .A(n673), .ZN(n671) );
  BUF_X1 U391 ( .A(n700), .Z(n590) );
  INV_X1 U392 ( .A(n593), .ZN(n454) );
  XNOR2_X1 U393 ( .A(n532), .B(n515), .ZN(n565) );
  INV_X1 U394 ( .A(n759), .ZN(n456) );
  INV_X1 U395 ( .A(G140), .ZN(n359) );
  INV_X1 U396 ( .A(G137), .ZN(n360) );
  INV_X1 U397 ( .A(KEYINPUT75), .ZN(n465) );
  AND2_X1 U398 ( .A1(n433), .A2(n434), .ZN(n391) );
  AND2_X1 U399 ( .A1(n437), .A2(n775), .ZN(n434) );
  XNOR2_X1 U400 ( .A(n386), .B(KEYINPUT108), .ZN(n775) );
  NAND2_X1 U401 ( .A1(n469), .A2(n468), .ZN(n670) );
  NOR2_X1 U402 ( .A1(n602), .A2(n605), .ZN(n562) );
  NAND2_X1 U403 ( .A1(n387), .A2(n590), .ZN(n398) );
  NOR2_X1 U404 ( .A1(n703), .A2(n702), .ZN(n595) );
  AND2_X1 U405 ( .A1(n441), .A2(n444), .ZN(n440) );
  OR2_X1 U406 ( .A1(n510), .A2(n445), .ZN(n441) );
  XNOR2_X1 U407 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U408 ( .A(n462), .B(n460), .ZN(n689) );
  XNOR2_X1 U409 ( .A(n480), .B(n565), .ZN(n493) );
  INV_X1 U410 ( .A(n741), .ZN(n431) );
  XNOR2_X1 U411 ( .A(n497), .B(n479), .ZN(n532) );
  NAND2_X1 U412 ( .A1(n361), .A2(n362), .ZN(n563) );
  INV_X1 U413 ( .A(n427), .ZN(n497) );
  XNOR2_X1 U414 ( .A(G902), .B(KEYINPUT15), .ZN(n542) );
  XNOR2_X1 U415 ( .A(KEYINPUT74), .B(KEYINPUT24), .ZN(n545) );
  XNOR2_X1 U416 ( .A(G143), .B(G128), .ZN(n427) );
  XNOR2_X1 U417 ( .A(KEYINPUT4), .B(KEYINPUT69), .ZN(n762) );
  XOR2_X1 U418 ( .A(G146), .B(G137), .Z(n491) );
  XNOR2_X2 U419 ( .A(n353), .B(n651), .ZN(n764) );
  NAND2_X1 U420 ( .A1(n397), .A2(n681), .ZN(n353) );
  XNOR2_X2 U421 ( .A(n354), .B(KEYINPUT87), .ZN(n397) );
  NAND2_X2 U422 ( .A1(n391), .A2(n435), .ZN(n354) );
  XNOR2_X2 U423 ( .A(G116), .B(KEYINPUT73), .ZN(n355) );
  BUF_X1 U424 ( .A(n764), .Z(n356) );
  NOR2_X1 U425 ( .A1(n737), .A2(n741), .ZN(n425) );
  XNOR2_X1 U426 ( .A(n475), .B(KEYINPUT35), .ZN(n774) );
  XNOR2_X1 U427 ( .A(n484), .B(n506), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n484), .B(n506), .ZN(n725) );
  XNOR2_X2 U429 ( .A(n393), .B(n742), .ZN(n484) );
  BUF_X1 U430 ( .A(n714), .Z(n358) );
  NAND2_X1 U431 ( .A1(G140), .A2(n360), .ZN(n361) );
  NAND2_X1 U432 ( .A1(n359), .A2(G137), .ZN(n362) );
  BUF_X1 U433 ( .A(n777), .Z(n363) );
  XNOR2_X1 U434 ( .A(n459), .B(n592), .ZN(n777) );
  NOR2_X2 U435 ( .A1(n739), .A2(G902), .ZN(n558) );
  INV_X1 U436 ( .A(n596), .ZN(n469) );
  XNOR2_X2 U437 ( .A(n398), .B(KEYINPUT39), .ZN(n648) );
  NAND2_X1 U438 ( .A1(n511), .A2(n449), .ZN(n448) );
  INV_X1 U439 ( .A(G902), .ZN(n449) );
  INV_X1 U440 ( .A(KEYINPUT86), .ZN(n651) );
  NAND2_X1 U441 ( .A1(n415), .A2(n588), .ZN(n601) );
  XOR2_X1 U442 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n544) );
  XNOR2_X1 U443 ( .A(n543), .B(KEYINPUT20), .ZN(n554) );
  NOR2_X1 U444 ( .A1(n601), .A2(KEYINPUT48), .ZN(n438) );
  INV_X1 U445 ( .A(n448), .ZN(n446) );
  NOR2_X1 U446 ( .A1(G902), .A2(G237), .ZN(n507) );
  XNOR2_X1 U447 ( .A(KEYINPUT70), .B(G131), .ZN(n515) );
  XNOR2_X1 U448 ( .A(n762), .B(G101), .ZN(n505) );
  XNOR2_X1 U449 ( .A(G125), .B(G146), .ZN(n516) );
  AND2_X1 U450 ( .A1(n689), .A2(n369), .ZN(n472) );
  NAND2_X1 U451 ( .A1(G214), .A2(n561), .ZN(n699) );
  INV_X1 U452 ( .A(KEYINPUT28), .ZN(n471) );
  NAND2_X1 U453 ( .A1(n383), .A2(n443), .ZN(n579) );
  OR2_X1 U454 ( .A1(n510), .A2(n448), .ZN(n443) );
  NOR2_X1 U455 ( .A1(n352), .A2(n371), .ZN(n383) );
  XNOR2_X1 U456 ( .A(n617), .B(KEYINPUT67), .ZN(n618) );
  INV_X1 U457 ( .A(KEYINPUT22), .ZN(n617) );
  XNOR2_X1 U458 ( .A(n419), .B(n418), .ZN(n417) );
  XNOR2_X1 U459 ( .A(n546), .B(KEYINPUT23), .ZN(n418) );
  XNOR2_X1 U460 ( .A(n563), .B(n545), .ZN(n419) );
  XNOR2_X1 U461 ( .A(KEYINPUT95), .B(KEYINPUT93), .ZN(n546) );
  XNOR2_X1 U462 ( .A(n516), .B(KEYINPUT10), .ZN(n759) );
  INV_X1 U463 ( .A(G134), .ZN(n479) );
  XOR2_X1 U464 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n526) );
  XOR2_X1 U465 ( .A(n390), .B(KEYINPUT9), .Z(n528) );
  XNOR2_X1 U466 ( .A(n530), .B(n529), .ZN(n531) );
  INV_X1 U467 ( .A(KEYINPUT7), .ZN(n529) );
  XNOR2_X1 U468 ( .A(G116), .B(G122), .ZN(n530) );
  XOR2_X1 U469 ( .A(G104), .B(G113), .Z(n514) );
  XNOR2_X1 U470 ( .A(G143), .B(G122), .ZN(n513) );
  INV_X1 U471 ( .A(n542), .ZN(n650) );
  XOR2_X1 U472 ( .A(KEYINPUT89), .B(KEYINPUT18), .Z(n501) );
  XNOR2_X1 U473 ( .A(KEYINPUT17), .B(KEYINPUT80), .ZN(n500) );
  XNOR2_X1 U474 ( .A(G122), .B(KEYINPUT16), .ZN(n485) );
  INV_X1 U475 ( .A(n536), .ZN(n765) );
  INV_X1 U476 ( .A(KEYINPUT66), .ZN(n405) );
  INV_X1 U477 ( .A(KEYINPUT105), .ZN(n406) );
  XNOR2_X1 U478 ( .A(n534), .B(G478), .ZN(n594) );
  OR2_X1 U479 ( .A1(n654), .A2(G902), .ZN(n534) );
  NOR2_X1 U480 ( .A1(n765), .A2(G952), .ZN(n741) );
  XNOR2_X1 U481 ( .A(n716), .B(KEYINPUT85), .ZN(n717) );
  INV_X1 U482 ( .A(KEYINPUT47), .ZN(n467) );
  INV_X1 U483 ( .A(KEYINPUT38), .ZN(n463) );
  XNOR2_X1 U484 ( .A(n544), .B(n461), .ZN(n460) );
  NAND2_X1 U485 ( .A1(n554), .A2(G221), .ZN(n462) );
  INV_X1 U486 ( .A(KEYINPUT21), .ZN(n461) );
  NOR2_X1 U487 ( .A1(n765), .A2(n537), .ZN(n538) );
  XNOR2_X1 U488 ( .A(n452), .B(n451), .ZN(n616) );
  INV_X1 U489 ( .A(KEYINPUT103), .ZN(n451) );
  OR2_X1 U490 ( .A1(n702), .A2(n615), .ZN(n452) );
  XNOR2_X1 U491 ( .A(n489), .B(KEYINPUT5), .ZN(n450) );
  NOR2_X1 U492 ( .A1(G953), .A2(G237), .ZN(n520) );
  XNOR2_X1 U493 ( .A(n565), .B(n564), .ZN(n758) );
  NAND2_X1 U494 ( .A1(G237), .A2(G234), .ZN(n535) );
  NAND2_X1 U495 ( .A1(n454), .A2(n453), .ZN(n702) );
  INV_X1 U496 ( .A(n594), .ZN(n453) );
  NOR2_X1 U497 ( .A1(n447), .A2(n511), .ZN(n439) );
  NAND2_X1 U498 ( .A1(n699), .A2(n371), .ZN(n444) );
  NAND2_X1 U499 ( .A1(n699), .A2(n446), .ZN(n445) );
  INV_X1 U500 ( .A(G104), .ZN(n420) );
  INV_X1 U501 ( .A(KEYINPUT19), .ZN(n486) );
  XNOR2_X1 U502 ( .A(n582), .B(n470), .ZN(n596) );
  INV_X1 U503 ( .A(KEYINPUT109), .ZN(n470) );
  XNOR2_X1 U504 ( .A(n409), .B(n471), .ZN(n581) );
  XNOR2_X1 U505 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U506 ( .A(n417), .B(n759), .ZN(n553) );
  XNOR2_X1 U507 ( .A(n532), .B(n533), .ZN(n654) );
  XNOR2_X1 U508 ( .A(n527), .B(n423), .ZN(n533) );
  XNOR2_X1 U509 ( .A(n531), .B(n528), .ZN(n423) );
  XNOR2_X1 U510 ( .A(n457), .B(n455), .ZN(n734) );
  XNOR2_X1 U511 ( .A(n523), .B(n456), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n458), .B(n522), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n476), .A2(n366), .ZN(n475) );
  XNOR2_X1 U514 ( .A(n629), .B(n373), .ZN(n630) );
  NOR2_X1 U515 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U516 ( .A1(n401), .A2(n688), .ZN(n400) );
  NOR2_X1 U517 ( .A1(n512), .A2(n405), .ZN(n401) );
  NOR2_X2 U518 ( .A1(n594), .A2(n454), .ZN(n673) );
  XNOR2_X1 U519 ( .A(n729), .B(n424), .ZN(n732) );
  XNOR2_X1 U520 ( .A(n388), .B(n730), .ZN(n424) );
  AND2_X1 U521 ( .A1(n723), .A2(n422), .ZN(n724) );
  AND2_X1 U522 ( .A1(n722), .A2(n753), .ZN(n422) );
  XNOR2_X1 U523 ( .A(n630), .B(n404), .ZN(G21) );
  INV_X1 U524 ( .A(G119), .ZN(n404) );
  AND2_X1 U525 ( .A1(n389), .A2(n369), .ZN(n364) );
  AND2_X1 U526 ( .A1(n512), .A2(n405), .ZN(n365) );
  XNOR2_X1 U527 ( .A(KEYINPUT81), .B(n623), .ZN(n366) );
  XOR2_X1 U528 ( .A(KEYINPUT82), .B(n649), .Z(n367) );
  AND2_X1 U529 ( .A1(n632), .A2(n699), .ZN(n368) );
  OR2_X1 U530 ( .A1(n541), .A2(n540), .ZN(n369) );
  OR2_X1 U531 ( .A1(n647), .A2(KEYINPUT44), .ZN(n370) );
  AND2_X1 U532 ( .A1(G472), .A2(G902), .ZN(n371) );
  AND2_X1 U533 ( .A1(n394), .A2(n395), .ZN(n372) );
  XOR2_X1 U534 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n373) );
  XOR2_X1 U535 ( .A(n510), .B(n496), .Z(n374) );
  INV_X1 U536 ( .A(KEYINPUT79), .ZN(n382) );
  INV_X1 U537 ( .A(G953), .ZN(n753) );
  NAND2_X1 U538 ( .A1(n394), .A2(n395), .ZN(n473) );
  INV_X1 U539 ( .A(n612), .ZN(n468) );
  NAND2_X1 U540 ( .A1(n764), .A2(n382), .ZN(n376) );
  INV_X1 U541 ( .A(n764), .ZN(n375) );
  OR2_X1 U542 ( .A1(n403), .A2(n405), .ZN(n395) );
  AND2_X1 U543 ( .A1(n414), .A2(n410), .ZN(n378) );
  AND2_X2 U544 ( .A1(n410), .A2(n414), .ZN(n396) );
  NAND2_X1 U545 ( .A1(n412), .A2(n411), .ZN(n410) );
  BUF_X1 U546 ( .A(n392), .Z(n379) );
  INV_X1 U547 ( .A(n639), .ZN(n380) );
  BUF_X1 U548 ( .A(n720), .Z(n381) );
  XNOR2_X1 U549 ( .A(n595), .B(KEYINPUT41), .ZN(n720) );
  INV_X1 U550 ( .A(KEYINPUT2), .ZN(n411) );
  XNOR2_X1 U551 ( .A(n646), .B(n483), .ZN(n384) );
  NAND2_X1 U552 ( .A1(n384), .A2(n370), .ZN(n482) );
  NAND2_X1 U553 ( .A1(n606), .A2(n605), .ZN(n386) );
  XNOR2_X1 U554 ( .A(n602), .B(KEYINPUT107), .ZN(n603) );
  NAND2_X1 U555 ( .A1(n560), .A2(n368), .ZN(n602) );
  XNOR2_X1 U556 ( .A(n525), .B(n524), .ZN(n593) );
  XNOR2_X1 U557 ( .A(n399), .B(n758), .ZN(n731) );
  XNOR2_X1 U558 ( .A(n589), .B(n463), .ZN(n700) );
  NOR2_X1 U559 ( .A1(n774), .A2(n630), .ZN(n474) );
  BUF_X1 U560 ( .A(n731), .Z(n388) );
  NAND2_X1 U561 ( .A1(n638), .A2(n632), .ZN(n477) );
  XNOR2_X1 U562 ( .A(n477), .B(n620), .ZN(n719) );
  XNOR2_X1 U563 ( .A(n575), .B(KEYINPUT30), .ZN(n389) );
  NAND2_X1 U564 ( .A1(n647), .A2(KEYINPUT44), .ZN(n645) );
  NAND2_X1 U565 ( .A1(n473), .A2(n474), .ZN(n647) );
  NAND2_X1 U566 ( .A1(n392), .A2(n428), .ZN(n714) );
  XNOR2_X1 U567 ( .A(n466), .B(n526), .ZN(n547) );
  NAND2_X1 U568 ( .A1(n392), .A2(n356), .ZN(n713) );
  NAND2_X1 U569 ( .A1(n379), .A2(n753), .ZN(n754) );
  NAND2_X1 U570 ( .A1(n413), .A2(n392), .ZN(n412) );
  XNOR2_X2 U571 ( .A(n482), .B(KEYINPUT45), .ZN(n392) );
  XNOR2_X1 U572 ( .A(n393), .B(n569), .ZN(n399) );
  XNOR2_X2 U573 ( .A(n407), .B(n505), .ZN(n393) );
  NAND2_X1 U574 ( .A1(n396), .A2(G478), .ZN(n653) );
  NAND2_X1 U575 ( .A1(n396), .A2(G210), .ZN(n727) );
  NAND2_X1 U576 ( .A1(n396), .A2(G475), .ZN(n736) );
  NAND2_X1 U577 ( .A1(n378), .A2(G472), .ZN(n652) );
  NAND2_X1 U578 ( .A1(n378), .A2(G217), .ZN(n738) );
  NAND2_X1 U579 ( .A1(n378), .A2(G469), .ZN(n729) );
  AND2_X1 U580 ( .A1(n397), .A2(n367), .ZN(n428) );
  NAND2_X1 U581 ( .A1(n648), .A2(n673), .ZN(n459) );
  NAND2_X1 U582 ( .A1(n403), .A2(n365), .ZN(n402) );
  XNOR2_X2 U583 ( .A(n504), .B(n485), .ZN(n742) );
  XNOR2_X2 U584 ( .A(n408), .B(n490), .ZN(n504) );
  XNOR2_X2 U585 ( .A(n421), .B(n420), .ZN(n745) );
  INV_X1 U586 ( .A(n536), .ZN(n566) );
  NAND2_X1 U587 ( .A1(n579), .A2(n578), .ZN(n409) );
  XNOR2_X2 U588 ( .A(n558), .B(n557), .ZN(n626) );
  NAND2_X1 U589 ( .A1(n601), .A2(KEYINPUT48), .ZN(n437) );
  NAND2_X1 U590 ( .A1(n416), .A2(n587), .ZN(n415) );
  XNOR2_X1 U591 ( .A(n586), .B(n467), .ZN(n416) );
  XNOR2_X2 U592 ( .A(G110), .B(G107), .ZN(n421) );
  XNOR2_X1 U593 ( .A(n519), .B(n521), .ZN(n458) );
  NAND2_X1 U594 ( .A1(n432), .A2(n431), .ZN(n430) );
  NOR2_X2 U595 ( .A1(n615), .A2(n626), .ZN(n684) );
  NOR2_X2 U596 ( .A1(n670), .A2(n704), .ZN(n586) );
  XNOR2_X1 U597 ( .A(n425), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U598 ( .A(n426), .B(KEYINPUT56), .ZN(G51) );
  BUF_X1 U599 ( .A(n589), .Z(n429) );
  INV_X2 U600 ( .A(n579), .ZN(n512) );
  XNOR2_X1 U601 ( .A(n652), .B(n374), .ZN(n432) );
  NOR2_X2 U602 ( .A1(n777), .A2(n776), .ZN(n599) );
  XNOR2_X1 U603 ( .A(n430), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U604 ( .A1(n364), .A2(n635), .ZN(n591) );
  XNOR2_X2 U605 ( .A(n576), .B(KEYINPUT99), .ZN(n635) );
  NAND2_X1 U606 ( .A1(n600), .A2(KEYINPUT48), .ZN(n433) );
  NAND2_X1 U607 ( .A1(n436), .A2(n438), .ZN(n435) );
  INV_X1 U608 ( .A(n600), .ZN(n436) );
  XNOR2_X2 U609 ( .A(n493), .B(n492), .ZN(n510) );
  NAND2_X1 U610 ( .A1(n510), .A2(n439), .ZN(n442) );
  NAND2_X1 U611 ( .A1(n442), .A2(n440), .ZN(n575) );
  INV_X1 U612 ( .A(n699), .ZN(n447) );
  XNOR2_X1 U613 ( .A(n505), .B(n450), .ZN(n480) );
  XNOR2_X2 U614 ( .A(n464), .B(n509), .ZN(n589) );
  NAND2_X1 U615 ( .A1(n725), .A2(n542), .ZN(n464) );
  NAND2_X1 U616 ( .A1(n547), .A2(G221), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n566), .A2(G234), .ZN(n466) );
  INV_X1 U618 ( .A(n624), .ZN(n476) );
  INV_X1 U619 ( .A(n512), .ZN(n687) );
  INV_X1 U620 ( .A(n625), .ZN(n683) );
  XNOR2_X2 U621 ( .A(n512), .B(KEYINPUT6), .ZN(n632) );
  INV_X1 U622 ( .A(n684), .ZN(n478) );
  AND2_X2 U623 ( .A1(n481), .A2(n625), .ZN(n631) );
  NAND2_X1 U624 ( .A1(n481), .A2(n626), .ZN(n627) );
  INV_X1 U625 ( .A(KEYINPUT88), .ZN(n483) );
  NOR2_X2 U626 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X2 U627 ( .A(n487), .B(n486), .ZN(n612) );
  NAND2_X1 U628 ( .A1(n589), .A2(n699), .ZN(n487) );
  XNOR2_X1 U629 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n488) );
  INV_X1 U630 ( .A(KEYINPUT46), .ZN(n598) );
  NOR2_X1 U631 ( .A1(n671), .A2(n559), .ZN(n560) );
  XNOR2_X1 U632 ( .A(n504), .B(n491), .ZN(n492) );
  XNOR2_X1 U633 ( .A(n570), .B(G469), .ZN(n571) );
  INV_X1 U634 ( .A(KEYINPUT25), .ZN(n555) );
  XNOR2_X1 U635 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U636 ( .A(n508), .B(KEYINPUT91), .ZN(n509) );
  XNOR2_X1 U637 ( .A(n552), .B(n553), .ZN(n739) );
  XNOR2_X1 U638 ( .A(n727), .B(n726), .ZN(n728) );
  INV_X1 U639 ( .A(KEYINPUT119), .ZN(n656) );
  AND2_X1 U640 ( .A1(n520), .A2(G210), .ZN(n489) );
  XNOR2_X1 U641 ( .A(KEYINPUT3), .B(G113), .ZN(n490) );
  XOR2_X1 U642 ( .A(KEYINPUT111), .B(KEYINPUT90), .Z(n495) );
  XNOR2_X1 U643 ( .A(KEYINPUT110), .B(KEYINPUT62), .ZN(n494) );
  XNOR2_X1 U644 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U645 ( .A(n497), .B(n516), .ZN(n499) );
  NAND2_X1 U646 ( .A1(G224), .A2(n765), .ZN(n498) );
  XNOR2_X1 U647 ( .A(n499), .B(n498), .ZN(n503) );
  XNOR2_X1 U648 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U649 ( .A(n503), .B(n502), .Z(n506) );
  XOR2_X1 U650 ( .A(KEYINPUT78), .B(n507), .Z(n561) );
  NAND2_X1 U651 ( .A1(G210), .A2(n561), .ZN(n508) );
  INV_X1 U652 ( .A(n429), .ZN(n605) );
  INV_X1 U653 ( .A(G472), .ZN(n511) );
  XNOR2_X1 U654 ( .A(n514), .B(n513), .ZN(n523) );
  XOR2_X1 U655 ( .A(n515), .B(KEYINPUT102), .Z(n522) );
  XOR2_X1 U656 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n518) );
  XNOR2_X1 U657 ( .A(G140), .B(KEYINPUT101), .ZN(n517) );
  XNOR2_X1 U658 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U659 ( .A1(n520), .A2(G214), .ZN(n521) );
  NOR2_X1 U660 ( .A1(G902), .A2(n734), .ZN(n525) );
  XNOR2_X1 U661 ( .A(KEYINPUT13), .B(G475), .ZN(n524) );
  NAND2_X1 U662 ( .A1(G217), .A2(n547), .ZN(n527) );
  NAND2_X1 U663 ( .A1(G952), .A2(n753), .ZN(n607) );
  XOR2_X1 U664 ( .A(n535), .B(KEYINPUT14), .Z(n610) );
  NOR2_X1 U665 ( .A1(n607), .A2(n610), .ZN(n541) );
  INV_X1 U666 ( .A(n610), .ZN(n682) );
  NAND2_X1 U667 ( .A1(G902), .A2(n682), .ZN(n537) );
  XOR2_X1 U668 ( .A(KEYINPUT106), .B(n538), .Z(n539) );
  NOR2_X1 U669 ( .A1(G900), .A2(n539), .ZN(n540) );
  NAND2_X1 U670 ( .A1(G234), .A2(n542), .ZN(n543) );
  XOR2_X1 U671 ( .A(KEYINPUT94), .B(G110), .Z(n549) );
  XNOR2_X1 U672 ( .A(G128), .B(G119), .ZN(n548) );
  XNOR2_X1 U673 ( .A(n549), .B(n548), .ZN(n550) );
  NAND2_X1 U674 ( .A1(G217), .A2(n554), .ZN(n556) );
  INV_X1 U675 ( .A(n578), .ZN(n559) );
  XNOR2_X1 U676 ( .A(n562), .B(KEYINPUT36), .ZN(n574) );
  INV_X1 U677 ( .A(n563), .ZN(n564) );
  XOR2_X1 U678 ( .A(G146), .B(KEYINPUT92), .Z(n568) );
  NAND2_X1 U679 ( .A1(G227), .A2(n765), .ZN(n567) );
  XNOR2_X1 U680 ( .A(n568), .B(n567), .ZN(n569) );
  NOR2_X2 U681 ( .A1(G902), .A2(n731), .ZN(n572) );
  XNOR2_X1 U682 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n570) );
  XNOR2_X2 U683 ( .A(n572), .B(n571), .ZN(n580) );
  XOR2_X1 U684 ( .A(KEYINPUT1), .B(KEYINPUT68), .Z(n573) );
  XNOR2_X1 U685 ( .A(n580), .B(n573), .ZN(n625) );
  NAND2_X1 U686 ( .A1(n574), .A2(n683), .ZN(n680) );
  NAND2_X1 U687 ( .A1(n594), .A2(n593), .ZN(n623) );
  XOR2_X1 U688 ( .A(KEYINPUT98), .B(n689), .Z(n615) );
  NAND2_X1 U689 ( .A1(n580), .A2(n684), .ZN(n576) );
  NOR2_X1 U690 ( .A1(n623), .A2(n591), .ZN(n577) );
  NAND2_X1 U691 ( .A1(n429), .A2(n577), .ZN(n668) );
  NAND2_X1 U692 ( .A1(n680), .A2(n668), .ZN(n585) );
  NAND2_X1 U693 ( .A1(n454), .A2(n594), .ZN(n664) );
  INV_X1 U694 ( .A(n664), .ZN(n676) );
  NOR2_X1 U695 ( .A1(n673), .A2(n676), .ZN(n704) );
  NAND2_X1 U696 ( .A1(n704), .A2(KEYINPUT83), .ZN(n583) );
  NAND2_X1 U697 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U698 ( .A1(n583), .A2(n670), .ZN(n584) );
  NOR2_X1 U699 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U700 ( .A1(n586), .A2(KEYINPUT83), .ZN(n587) );
  INV_X1 U701 ( .A(KEYINPUT40), .ZN(n592) );
  NAND2_X1 U702 ( .A1(n700), .A2(n699), .ZN(n703) );
  NOR2_X1 U703 ( .A1(n596), .A2(n720), .ZN(n597) );
  XNOR2_X1 U704 ( .A(n597), .B(KEYINPUT42), .ZN(n776) );
  XNOR2_X1 U705 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U706 ( .A1(n603), .A2(n625), .ZN(n604) );
  XNOR2_X1 U707 ( .A(n604), .B(KEYINPUT43), .ZN(n606) );
  NOR2_X1 U708 ( .A1(G898), .A2(n753), .ZN(n747) );
  NAND2_X1 U709 ( .A1(n747), .A2(G902), .ZN(n608) );
  AND2_X1 U710 ( .A1(n608), .A2(n607), .ZN(n609) );
  OR2_X1 U711 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U712 ( .A(KEYINPUT0), .ZN(n613) );
  INV_X1 U713 ( .A(n626), .ZN(n688) );
  XNOR2_X1 U714 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n622) );
  XOR2_X1 U715 ( .A(KEYINPUT33), .B(KEYINPUT76), .Z(n620) );
  NOR2_X1 U716 ( .A1(n380), .A2(n719), .ZN(n621) );
  XNOR2_X1 U717 ( .A(n622), .B(n621), .ZN(n624) );
  OR2_X1 U718 ( .A1(n625), .A2(n632), .ZN(n628) );
  NAND2_X1 U719 ( .A1(n631), .A2(n688), .ZN(n633) );
  NOR2_X1 U720 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U721 ( .A(n634), .B(KEYINPUT104), .ZN(n778) );
  XOR2_X1 U722 ( .A(n704), .B(KEYINPUT83), .Z(n642) );
  INV_X1 U723 ( .A(n619), .ZN(n639) );
  AND2_X1 U724 ( .A1(n639), .A2(n635), .ZN(n636) );
  XOR2_X1 U725 ( .A(KEYINPUT100), .B(n636), .Z(n637) );
  AND2_X1 U726 ( .A1(n687), .A2(n638), .ZN(n695) );
  NAND2_X1 U727 ( .A1(n639), .A2(n695), .ZN(n640) );
  XNOR2_X1 U728 ( .A(n640), .B(KEYINPUT31), .ZN(n677) );
  NOR2_X1 U729 ( .A1(n660), .A2(n677), .ZN(n641) );
  NOR2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U731 ( .A1(n778), .A2(n643), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n676), .A2(n648), .ZN(n681) );
  NAND2_X1 U734 ( .A1(KEYINPUT2), .A2(n681), .ZN(n649) );
  XNOR2_X1 U735 ( .A(n653), .B(n654), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n657), .B(n656), .ZN(G63) );
  NAND2_X1 U737 ( .A1(n660), .A2(n673), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(KEYINPUT112), .ZN(n659) );
  XNOR2_X1 U739 ( .A(G104), .B(n659), .ZN(G6) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n662) );
  NAND2_X1 U741 ( .A1(n660), .A2(n676), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U743 ( .A(n390), .B(n663), .ZN(G9) );
  XOR2_X1 U744 ( .A(G110), .B(n372), .Z(G12) );
  NOR2_X1 U745 ( .A1(n664), .A2(n670), .ZN(n666) );
  XNOR2_X1 U746 ( .A(KEYINPUT29), .B(KEYINPUT113), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U748 ( .A(G128), .B(n667), .Z(G30) );
  XNOR2_X1 U749 ( .A(G143), .B(KEYINPUT114), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(n668), .ZN(G45) );
  NOR2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U752 ( .A(G146), .B(n672), .Z(G48) );
  XOR2_X1 U753 ( .A(G113), .B(KEYINPUT115), .Z(n675) );
  NAND2_X1 U754 ( .A1(n677), .A2(n673), .ZN(n674) );
  XNOR2_X1 U755 ( .A(n675), .B(n674), .ZN(G15) );
  NAND2_X1 U756 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n678), .B(G116), .ZN(G18) );
  XOR2_X1 U758 ( .A(G125), .B(KEYINPUT37), .Z(n679) );
  XNOR2_X1 U759 ( .A(n680), .B(n679), .ZN(G27) );
  XNOR2_X1 U760 ( .A(G134), .B(n681), .ZN(G36) );
  NAND2_X1 U761 ( .A1(G952), .A2(n682), .ZN(n712) );
  NOR2_X1 U762 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U763 ( .A(n685), .B(KEYINPUT50), .ZN(n686) );
  NOR2_X1 U764 ( .A1(n687), .A2(n686), .ZN(n692) );
  NOR2_X1 U765 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U766 ( .A(n690), .B(KEYINPUT49), .ZN(n691) );
  NAND2_X1 U767 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U768 ( .A(KEYINPUT116), .B(n693), .Z(n694) );
  NOR2_X1 U769 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U770 ( .A(n696), .B(KEYINPUT51), .ZN(n697) );
  XNOR2_X1 U771 ( .A(KEYINPUT117), .B(n697), .ZN(n698) );
  NOR2_X1 U772 ( .A1(n381), .A2(n698), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n590), .A2(n699), .ZN(n701) );
  NOR2_X1 U774 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U775 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U777 ( .A1(n719), .A2(n707), .ZN(n708) );
  NOR2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U779 ( .A(n710), .B(KEYINPUT52), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U781 ( .A1(n713), .A2(n411), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n715), .A2(n358), .ZN(n716) );
  NOR2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n723) );
  NOR2_X1 U784 ( .A1(n381), .A2(n719), .ZN(n721) );
  XOR2_X1 U785 ( .A(KEYINPUT118), .B(n721), .Z(n722) );
  XNOR2_X1 U786 ( .A(n724), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U787 ( .A(n357), .B(n488), .ZN(n726) );
  XOR2_X1 U788 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n730) );
  NOR2_X1 U789 ( .A1(n741), .A2(n732), .ZN(G54) );
  INV_X1 U790 ( .A(KEYINPUT59), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U792 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U793 ( .A1(n741), .A2(n740), .ZN(G66) );
  XNOR2_X1 U794 ( .A(n742), .B(G101), .ZN(n743) );
  XNOR2_X1 U795 ( .A(n743), .B(KEYINPUT123), .ZN(n744) );
  XOR2_X1 U796 ( .A(n745), .B(n744), .Z(n746) );
  NOR2_X1 U797 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U798 ( .A(KEYINPUT122), .B(n748), .Z(n757) );
  XOR2_X1 U799 ( .A(KEYINPUT61), .B(KEYINPUT121), .Z(n750) );
  NAND2_X1 U800 ( .A1(G224), .A2(G953), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n750), .B(n749), .ZN(n751) );
  XNOR2_X1 U802 ( .A(KEYINPUT120), .B(n751), .ZN(n752) );
  NAND2_X1 U803 ( .A1(n752), .A2(G898), .ZN(n755) );
  NAND2_X1 U804 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U805 ( .A(n757), .B(n756), .Z(G69) );
  XOR2_X1 U806 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n761) );
  XNOR2_X1 U807 ( .A(n759), .B(n758), .ZN(n760) );
  XNOR2_X1 U808 ( .A(n761), .B(n760), .ZN(n763) );
  XOR2_X1 U809 ( .A(n762), .B(n763), .Z(n769) );
  XNOR2_X1 U810 ( .A(n356), .B(n769), .ZN(n766) );
  NAND2_X1 U811 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U812 ( .A(n767), .B(KEYINPUT126), .ZN(n773) );
  XNOR2_X1 U813 ( .A(G227), .B(KEYINPUT127), .ZN(n768) );
  XNOR2_X1 U814 ( .A(n769), .B(n768), .ZN(n770) );
  NAND2_X1 U815 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U816 ( .A1(n771), .A2(G953), .ZN(n772) );
  NAND2_X1 U817 ( .A1(n773), .A2(n772), .ZN(G72) );
  XOR2_X1 U818 ( .A(G122), .B(n774), .Z(G24) );
  XNOR2_X1 U819 ( .A(G140), .B(n775), .ZN(G42) );
  XOR2_X1 U820 ( .A(n776), .B(G137), .Z(G39) );
  XOR2_X1 U821 ( .A(n363), .B(G131), .Z(G33) );
  XOR2_X1 U822 ( .A(G101), .B(n778), .Z(G3) );
endmodule

