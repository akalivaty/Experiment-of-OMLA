

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(KEYINPUT98), .ZN(n753) );
  NOR2_X2 U550 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XNOR2_X1 U551 ( .A(KEYINPUT23), .B(n518), .ZN(n515) );
  AND2_X1 U552 ( .A1(n521), .A2(n520), .ZN(n516) );
  AND2_X1 U553 ( .A1(n724), .A2(n723), .ZN(n727) );
  INV_X1 U554 ( .A(KEYINPUT96), .ZN(n725) );
  INV_X1 U555 ( .A(n728), .ZN(n759) );
  NOR2_X1 U556 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U557 ( .A1(n808), .A2(n807), .ZN(n809) );
  INV_X1 U558 ( .A(KEYINPUT67), .ZN(n523) );
  XNOR2_X1 U559 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U560 ( .A(G2105), .ZN(n519) );
  AND2_X1 U561 ( .A1(G2104), .A2(n519), .ZN(n517) );
  XNOR2_X2 U562 ( .A(n517), .B(KEYINPUT66), .ZN(n882) );
  NAND2_X1 U563 ( .A1(n882), .A2(G101), .ZN(n518) );
  AND2_X1 U564 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U565 ( .A1(G113), .A2(n885), .ZN(n521) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n519), .ZN(n886) );
  NAND2_X1 U567 ( .A1(G125), .A2(n886), .ZN(n520) );
  XOR2_X2 U568 ( .A(KEYINPUT17), .B(n522), .Z(n881) );
  NAND2_X1 U569 ( .A1(G137), .A2(n881), .ZN(n524) );
  NAND2_X1 U570 ( .A1(n516), .A2(n525), .ZN(n526) );
  NOR2_X2 U571 ( .A1(n515), .A2(n526), .ZN(G160) );
  XOR2_X1 U572 ( .A(G2443), .B(G2446), .Z(n528) );
  XNOR2_X1 U573 ( .A(G2427), .B(G2451), .ZN(n527) );
  XNOR2_X1 U574 ( .A(n528), .B(n527), .ZN(n534) );
  XOR2_X1 U575 ( .A(G2430), .B(G2454), .Z(n530) );
  XNOR2_X1 U576 ( .A(G1348), .B(G1341), .ZN(n529) );
  XNOR2_X1 U577 ( .A(n530), .B(n529), .ZN(n532) );
  XOR2_X1 U578 ( .A(G2435), .B(G2438), .Z(n531) );
  XNOR2_X1 U579 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U580 ( .A(n534), .B(n533), .Z(n535) );
  AND2_X1 U581 ( .A1(G14), .A2(n535), .ZN(G401) );
  AND2_X1 U582 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U583 ( .A(G57), .ZN(G237) );
  INV_X1 U584 ( .A(G132), .ZN(G219) );
  INV_X1 U585 ( .A(G82), .ZN(G220) );
  NOR2_X1 U586 ( .A1(G543), .A2(G651), .ZN(n536) );
  XOR2_X1 U587 ( .A(KEYINPUT65), .B(n536), .Z(n645) );
  NAND2_X1 U588 ( .A1(G88), .A2(n645), .ZN(n539) );
  INV_X1 U589 ( .A(G651), .ZN(n540) );
  XOR2_X1 U590 ( .A(G543), .B(KEYINPUT0), .Z(n642) );
  OR2_X1 U591 ( .A1(n540), .A2(n642), .ZN(n537) );
  XOR2_X1 U592 ( .A(KEYINPUT68), .B(n537), .Z(n653) );
  NAND2_X1 U593 ( .A1(G75), .A2(n653), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n546) );
  NOR2_X1 U595 ( .A1(G651), .A2(n642), .ZN(n646) );
  NAND2_X1 U596 ( .A1(G50), .A2(n646), .ZN(n544) );
  NOR2_X1 U597 ( .A1(G543), .A2(n540), .ZN(n542) );
  XNOR2_X1 U598 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n542), .B(n541), .ZN(n649) );
  NAND2_X1 U600 ( .A1(G62), .A2(n649), .ZN(n543) );
  NAND2_X1 U601 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U602 ( .A1(n546), .A2(n545), .ZN(G166) );
  NAND2_X1 U603 ( .A1(n649), .A2(G64), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT71), .B(n547), .Z(n549) );
  NAND2_X1 U605 ( .A1(n646), .A2(G52), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U607 ( .A(KEYINPUT72), .B(n550), .ZN(n556) );
  NAND2_X1 U608 ( .A1(G77), .A2(n653), .ZN(n551) );
  XOR2_X1 U609 ( .A(KEYINPUT73), .B(n551), .Z(n553) );
  NAND2_X1 U610 ( .A1(n645), .A2(G90), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U613 ( .A1(n556), .A2(n555), .ZN(G171) );
  INV_X1 U614 ( .A(G171), .ZN(G301) );
  NAND2_X1 U615 ( .A1(G89), .A2(n645), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n557), .B(KEYINPUT4), .ZN(n558) );
  XNOR2_X1 U617 ( .A(KEYINPUT80), .B(n558), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G76), .A2(n653), .ZN(n559) );
  XOR2_X1 U619 ( .A(KEYINPUT81), .B(n559), .Z(n560) );
  NAND2_X1 U620 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n562), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G51), .A2(n646), .ZN(n564) );
  NAND2_X1 U623 ( .A1(G63), .A2(n649), .ZN(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U625 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U626 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U628 ( .A(G168), .B(KEYINPUT8), .Z(n569) );
  XNOR2_X1 U629 ( .A(KEYINPUT82), .B(n569), .ZN(G286) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n572) );
  INV_X1 U633 ( .A(G223), .ZN(n829) );
  NAND2_X1 U634 ( .A1(G567), .A2(n829), .ZN(n571) );
  XNOR2_X1 U635 ( .A(n572), .B(n571), .ZN(G234) );
  XOR2_X1 U636 ( .A(KEYINPUT12), .B(KEYINPUT76), .Z(n574) );
  NAND2_X1 U637 ( .A1(G81), .A2(n645), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT75), .B(n575), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G68), .A2(n653), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT13), .B(n578), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G43), .A2(n646), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT77), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G56), .A2(n649), .ZN(n580) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n580), .Z(n581) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n974) );
  INV_X1 U649 ( .A(G860), .ZN(n605) );
  OR2_X1 U650 ( .A1(n974), .A2(n605), .ZN(G153) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U652 ( .A1(G92), .A2(n645), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G66), .A2(n649), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U655 ( .A(KEYINPUT78), .B(n587), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G54), .A2(n646), .ZN(n588) );
  XNOR2_X1 U657 ( .A(KEYINPUT79), .B(n588), .ZN(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G79), .A2(n653), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U661 ( .A(KEYINPUT15), .B(n593), .ZN(n958) );
  OR2_X1 U662 ( .A1(n958), .A2(G868), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U664 ( .A1(G53), .A2(n646), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G65), .A2(n649), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G91), .A2(n645), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G78), .A2(n653), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n968) );
  INV_X1 U671 ( .A(n968), .ZN(G299) );
  INV_X1 U672 ( .A(G868), .ZN(n664) );
  NOR2_X1 U673 ( .A1(G286), .A2(n664), .ZN(n602) );
  XOR2_X1 U674 ( .A(KEYINPUT83), .B(n602), .Z(n604) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n603) );
  NOR2_X1 U676 ( .A1(n604), .A2(n603), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n605), .A2(G559), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n606), .A2(n958), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n974), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G868), .A2(n958), .ZN(n608) );
  NOR2_X1 U682 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G99), .A2(n882), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G111), .A2(n885), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G135), .A2(n881), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n886), .A2(G123), .ZN(n613) );
  XOR2_X1 U689 ( .A(KEYINPUT18), .B(n613), .Z(n614) );
  NOR2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U692 ( .A(KEYINPUT84), .B(n618), .Z(n938) );
  XOR2_X1 U693 ( .A(G2096), .B(n938), .Z(n619) );
  NOR2_X1 U694 ( .A1(G2100), .A2(n619), .ZN(n620) );
  XNOR2_X1 U695 ( .A(KEYINPUT85), .B(n620), .ZN(G156) );
  NAND2_X1 U696 ( .A1(G55), .A2(n646), .ZN(n622) );
  NAND2_X1 U697 ( .A1(G80), .A2(n653), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U699 ( .A1(n645), .A2(G93), .ZN(n623) );
  XOR2_X1 U700 ( .A(KEYINPUT86), .B(n623), .Z(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n649), .A2(G67), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n665) );
  NAND2_X1 U704 ( .A1(n958), .A2(G559), .ZN(n662) );
  XNOR2_X1 U705 ( .A(n974), .B(n662), .ZN(n628) );
  NOR2_X1 U706 ( .A1(G860), .A2(n628), .ZN(n629) );
  XOR2_X1 U707 ( .A(n665), .B(n629), .Z(G145) );
  NAND2_X1 U708 ( .A1(G73), .A2(n653), .ZN(n631) );
  XNOR2_X1 U709 ( .A(KEYINPUT88), .B(KEYINPUT2), .ZN(n630) );
  XNOR2_X1 U710 ( .A(n631), .B(n630), .ZN(n638) );
  NAND2_X1 U711 ( .A1(G48), .A2(n646), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G61), .A2(n649), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G86), .A2(n645), .ZN(n634) );
  XNOR2_X1 U715 ( .A(KEYINPUT87), .B(n634), .ZN(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G49), .A2(n646), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U721 ( .A1(n649), .A2(n641), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n642), .A2(G87), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U724 ( .A1(G85), .A2(n645), .ZN(n648) );
  NAND2_X1 U725 ( .A1(G47), .A2(n646), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G60), .A2(n649), .ZN(n650) );
  XOR2_X1 U728 ( .A(KEYINPUT70), .B(n650), .Z(n651) );
  NOR2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n655) );
  NAND2_X1 U730 ( .A1(G72), .A2(n653), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(G290) );
  XNOR2_X1 U732 ( .A(KEYINPUT19), .B(G305), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n656), .B(G288), .ZN(n657) );
  XNOR2_X1 U734 ( .A(G166), .B(n657), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n974), .B(n968), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n660), .B(G290), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n661), .B(n665), .ZN(n898) );
  XOR2_X1 U739 ( .A(n898), .B(n662), .Z(n663) );
  NAND2_X1 U740 ( .A1(G868), .A2(n663), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U748 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n672) );
  XNOR2_X1 U750 ( .A(KEYINPUT22), .B(n672), .ZN(n673) );
  NAND2_X1 U751 ( .A1(n673), .A2(G96), .ZN(n674) );
  NOR2_X1 U752 ( .A1(n674), .A2(G218), .ZN(n675) );
  XNOR2_X1 U753 ( .A(n675), .B(KEYINPUT89), .ZN(n834) );
  NAND2_X1 U754 ( .A1(n834), .A2(G2106), .ZN(n680) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n676) );
  NOR2_X1 U756 ( .A1(G237), .A2(n676), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G108), .A2(n677), .ZN(n833) );
  NAND2_X1 U758 ( .A1(G567), .A2(n833), .ZN(n678) );
  XNOR2_X1 U759 ( .A(KEYINPUT90), .B(n678), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n680), .A2(n679), .ZN(n835) );
  NAND2_X1 U761 ( .A1(G661), .A2(G483), .ZN(n681) );
  NOR2_X1 U762 ( .A1(n835), .A2(n681), .ZN(n832) );
  NAND2_X1 U763 ( .A1(n832), .A2(G36), .ZN(n682) );
  XOR2_X1 U764 ( .A(KEYINPUT91), .B(n682), .Z(G176) );
  NAND2_X1 U765 ( .A1(n885), .A2(G114), .ZN(n683) );
  XNOR2_X1 U766 ( .A(n683), .B(KEYINPUT92), .ZN(n685) );
  NAND2_X1 U767 ( .A1(G138), .A2(n881), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U769 ( .A1(n886), .A2(G126), .ZN(n687) );
  NAND2_X1 U770 ( .A1(G102), .A2(n882), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U772 ( .A1(n689), .A2(n688), .ZN(G164) );
  INV_X1 U773 ( .A(G166), .ZN(G303) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n716) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n714) );
  NOR2_X1 U776 ( .A1(n716), .A2(n714), .ZN(n824) );
  NAND2_X1 U777 ( .A1(n882), .A2(G105), .ZN(n690) );
  XNOR2_X1 U778 ( .A(n690), .B(KEYINPUT38), .ZN(n697) );
  NAND2_X1 U779 ( .A1(G141), .A2(n881), .ZN(n692) );
  NAND2_X1 U780 ( .A1(G129), .A2(n886), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U782 ( .A1(G117), .A2(n885), .ZN(n693) );
  XNOR2_X1 U783 ( .A(KEYINPUT93), .B(n693), .ZN(n694) );
  NOR2_X1 U784 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n869) );
  AND2_X1 U786 ( .A1(n869), .A2(G1996), .ZN(n945) );
  NAND2_X1 U787 ( .A1(G107), .A2(n885), .ZN(n699) );
  NAND2_X1 U788 ( .A1(G131), .A2(n881), .ZN(n698) );
  NAND2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n886), .A2(G119), .ZN(n701) );
  NAND2_X1 U791 ( .A1(G95), .A2(n882), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n702) );
  OR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n866) );
  AND2_X1 U794 ( .A1(n866), .A2(G1991), .ZN(n939) );
  OR2_X1 U795 ( .A1(n945), .A2(n939), .ZN(n704) );
  NAND2_X1 U796 ( .A1(n824), .A2(n704), .ZN(n811) );
  NAND2_X1 U797 ( .A1(G140), .A2(n881), .ZN(n706) );
  NAND2_X1 U798 ( .A1(G104), .A2(n882), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U800 ( .A(KEYINPUT34), .B(n707), .ZN(n712) );
  NAND2_X1 U801 ( .A1(G116), .A2(n885), .ZN(n709) );
  NAND2_X1 U802 ( .A1(G128), .A2(n886), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U804 ( .A(KEYINPUT35), .B(n710), .Z(n711) );
  NOR2_X1 U805 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U806 ( .A(KEYINPUT36), .B(n713), .ZN(n894) );
  XNOR2_X1 U807 ( .A(KEYINPUT37), .B(G2067), .ZN(n822) );
  NOR2_X1 U808 ( .A1(n894), .A2(n822), .ZN(n931) );
  NAND2_X1 U809 ( .A1(n824), .A2(n931), .ZN(n820) );
  AND2_X1 U810 ( .A1(n811), .A2(n820), .ZN(n810) );
  XNOR2_X1 U811 ( .A(G1981), .B(G305), .ZN(n960) );
  INV_X1 U812 ( .A(KEYINPUT33), .ZN(n785) );
  XOR2_X1 U813 ( .A(KEYINPUT94), .B(n714), .Z(n715) );
  NAND2_X1 U814 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n721), .A2(G8), .ZN(n802) );
  INV_X1 U816 ( .A(n802), .ZN(n796) );
  NOR2_X1 U817 ( .A1(G1976), .A2(G288), .ZN(n971) );
  NAND2_X1 U818 ( .A1(n796), .A2(n971), .ZN(n717) );
  NOR2_X1 U819 ( .A1(n785), .A2(n717), .ZN(n718) );
  XOR2_X1 U820 ( .A(n718), .B(KEYINPUT102), .Z(n793) );
  INV_X1 U821 ( .A(n721), .ZN(n728) );
  AND2_X1 U822 ( .A1(n728), .A2(G1996), .ZN(n720) );
  XOR2_X1 U823 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n719) );
  XNOR2_X1 U824 ( .A(n720), .B(n719), .ZN(n724) );
  AND2_X1 U825 ( .A1(n721), .A2(G1341), .ZN(n722) );
  NOR2_X1 U826 ( .A1(n722), .A2(n974), .ZN(n723) );
  NOR2_X1 U827 ( .A1(n727), .A2(n958), .ZN(n726) );
  XNOR2_X1 U828 ( .A(n726), .B(n725), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n727), .A2(n958), .ZN(n732) );
  NOR2_X1 U830 ( .A1(n728), .A2(G1348), .ZN(n730) );
  NOR2_X1 U831 ( .A1(G2067), .A2(n759), .ZN(n729) );
  NOR2_X1 U832 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U833 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U834 ( .A1(n734), .A2(n733), .ZN(n739) );
  NAND2_X1 U835 ( .A1(n728), .A2(G2072), .ZN(n735) );
  XNOR2_X1 U836 ( .A(n735), .B(KEYINPUT27), .ZN(n737) );
  INV_X1 U837 ( .A(G1956), .ZN(n969) );
  NOR2_X1 U838 ( .A1(n969), .A2(n728), .ZN(n736) );
  NOR2_X1 U839 ( .A1(n737), .A2(n736), .ZN(n740) );
  NAND2_X1 U840 ( .A1(n968), .A2(n740), .ZN(n738) );
  NAND2_X1 U841 ( .A1(n739), .A2(n738), .ZN(n743) );
  NOR2_X1 U842 ( .A1(n968), .A2(n740), .ZN(n741) );
  XOR2_X1 U843 ( .A(n741), .B(KEYINPUT28), .Z(n742) );
  NAND2_X1 U844 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U845 ( .A(n744), .B(KEYINPUT29), .ZN(n748) );
  NAND2_X1 U846 ( .A1(G1961), .A2(n759), .ZN(n746) );
  XOR2_X1 U847 ( .A(G2078), .B(KEYINPUT25), .Z(n917) );
  NAND2_X1 U848 ( .A1(n728), .A2(n917), .ZN(n745) );
  NAND2_X1 U849 ( .A1(n746), .A2(n745), .ZN(n755) );
  NOR2_X1 U850 ( .A1(G301), .A2(n755), .ZN(n747) );
  XNOR2_X1 U851 ( .A(n749), .B(KEYINPUT97), .ZN(n775) );
  NOR2_X1 U852 ( .A1(G1966), .A2(n802), .ZN(n778) );
  NOR2_X1 U853 ( .A1(G2084), .A2(n759), .ZN(n776) );
  NOR2_X1 U854 ( .A1(n778), .A2(n776), .ZN(n750) );
  NAND2_X1 U855 ( .A1(G8), .A2(n750), .ZN(n751) );
  XNOR2_X1 U856 ( .A(KEYINPUT30), .B(n751), .ZN(n752) );
  NOR2_X1 U857 ( .A1(G168), .A2(n752), .ZN(n754) );
  XNOR2_X1 U858 ( .A(n754), .B(n753), .ZN(n757) );
  NAND2_X1 U859 ( .A1(G301), .A2(n755), .ZN(n756) );
  NAND2_X1 U860 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U861 ( .A(KEYINPUT31), .B(n758), .ZN(n774) );
  INV_X1 U862 ( .A(G8), .ZN(n766) );
  NOR2_X1 U863 ( .A1(G1971), .A2(n802), .ZN(n761) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n759), .ZN(n760) );
  NOR2_X1 U865 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U866 ( .A(n762), .B(KEYINPUT99), .ZN(n763) );
  NOR2_X1 U867 ( .A1(G166), .A2(n763), .ZN(n764) );
  XOR2_X1 U868 ( .A(KEYINPUT100), .B(n764), .Z(n765) );
  OR2_X1 U869 ( .A1(n766), .A2(n765), .ZN(n768) );
  AND2_X1 U870 ( .A1(n774), .A2(n768), .ZN(n767) );
  NAND2_X1 U871 ( .A1(n775), .A2(n767), .ZN(n772) );
  INV_X1 U872 ( .A(n768), .ZN(n770) );
  AND2_X1 U873 ( .A1(G286), .A2(G8), .ZN(n769) );
  OR2_X1 U874 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U875 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U876 ( .A(n773), .B(KEYINPUT32), .ZN(n783) );
  AND2_X1 U877 ( .A1(n775), .A2(n774), .ZN(n781) );
  NAND2_X1 U878 ( .A1(G8), .A2(n776), .ZN(n777) );
  XNOR2_X1 U879 ( .A(KEYINPUT95), .B(n777), .ZN(n779) );
  OR2_X1 U880 ( .A1(n779), .A2(n778), .ZN(n780) );
  OR2_X1 U881 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U882 ( .A1(n783), .A2(n782), .ZN(n800) );
  NOR2_X1 U883 ( .A1(G1971), .A2(G303), .ZN(n784) );
  NOR2_X1 U884 ( .A1(n971), .A2(n784), .ZN(n786) );
  AND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U886 ( .A1(n800), .A2(n787), .ZN(n791) );
  NAND2_X1 U887 ( .A1(G288), .A2(G1976), .ZN(n788) );
  XNOR2_X1 U888 ( .A(n788), .B(KEYINPUT101), .ZN(n967) );
  NOR2_X1 U889 ( .A1(n967), .A2(n802), .ZN(n789) );
  OR2_X1 U890 ( .A1(KEYINPUT33), .A2(n789), .ZN(n790) );
  AND2_X1 U891 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U892 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U893 ( .A1(n960), .A2(n794), .ZN(n806) );
  NOR2_X1 U894 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XNOR2_X1 U895 ( .A(KEYINPUT24), .B(n795), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n804) );
  NOR2_X1 U897 ( .A1(G2090), .A2(G303), .ZN(n798) );
  NAND2_X1 U898 ( .A1(G8), .A2(n798), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n808) );
  XNOR2_X1 U903 ( .A(G1986), .B(G290), .ZN(n980) );
  AND2_X1 U904 ( .A1(n980), .A2(n824), .ZN(n807) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n827) );
  XOR2_X1 U906 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n819) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n869), .ZN(n946) );
  INV_X1 U908 ( .A(n811), .ZN(n815) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n866), .ZN(n812) );
  XOR2_X1 U910 ( .A(KEYINPUT103), .B(n812), .Z(n941) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n813) );
  NOR2_X1 U912 ( .A1(n941), .A2(n813), .ZN(n814) );
  NOR2_X1 U913 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U914 ( .A(n816), .B(KEYINPUT104), .ZN(n817) );
  NOR2_X1 U915 ( .A1(n946), .A2(n817), .ZN(n818) );
  XNOR2_X1 U916 ( .A(n819), .B(n818), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n894), .A2(n822), .ZN(n930) );
  NAND2_X1 U919 ( .A1(n823), .A2(n930), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n828), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n829), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U925 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U927 ( .A1(n832), .A2(n831), .ZN(G188) );
  NOR2_X1 U928 ( .A1(n834), .A2(n833), .ZN(G325) );
  XOR2_X1 U929 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  INV_X1 U934 ( .A(n835), .ZN(G319) );
  XOR2_X1 U935 ( .A(KEYINPUT109), .B(G1976), .Z(n837) );
  XNOR2_X1 U936 ( .A(G1986), .B(G1961), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U938 ( .A(n838), .B(KEYINPUT41), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U941 ( .A(G1981), .B(G1971), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1966), .B(G1956), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U945 ( .A(KEYINPUT110), .B(G2474), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(G229) );
  XOR2_X1 U947 ( .A(G2678), .B(KEYINPUT43), .Z(n848) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(KEYINPUT107), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U950 ( .A(KEYINPUT108), .B(G2090), .Z(n850) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U954 ( .A(G2096), .B(G2100), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n856) );
  XOR2_X1 U956 ( .A(G2078), .B(G2084), .Z(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G112), .A2(n885), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G100), .A2(n882), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U961 ( .A1(n886), .A2(G124), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G136), .A2(n881), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U965 ( .A(KEYINPUT111), .B(n862), .Z(n863) );
  NOR2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U967 ( .A(KEYINPUT112), .B(n865), .ZN(G162) );
  XOR2_X1 U968 ( .A(n866), .B(KEYINPUT46), .Z(n867) );
  XNOR2_X1 U969 ( .A(n867), .B(KEYINPUT48), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n938), .B(n868), .ZN(n871) );
  XOR2_X1 U971 ( .A(G160), .B(n869), .Z(n870) );
  XNOR2_X1 U972 ( .A(n871), .B(n870), .ZN(n880) );
  NAND2_X1 U973 ( .A1(G118), .A2(n885), .ZN(n873) );
  NAND2_X1 U974 ( .A1(G130), .A2(n886), .ZN(n872) );
  NAND2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G142), .A2(n881), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G106), .A2(n882), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  NOR2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(n880), .B(n879), .Z(n893) );
  NAND2_X1 U982 ( .A1(G139), .A2(n881), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G103), .A2(n882), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n891) );
  NAND2_X1 U985 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U987 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n933) );
  XNOR2_X1 U990 ( .A(G164), .B(n933), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n895) );
  XOR2_X1 U992 ( .A(n895), .B(n894), .Z(n896) );
  XNOR2_X1 U993 ( .A(G162), .B(n896), .ZN(n897) );
  NOR2_X1 U994 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U995 ( .A(KEYINPUT113), .B(n898), .Z(n900) );
  XNOR2_X1 U996 ( .A(G171), .B(n958), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(G286), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G397) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n903) );
  XOR2_X1 U1001 ( .A(KEYINPUT49), .B(n903), .Z(n904) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n904), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n905), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT114), .B(n906), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1009 ( .A(G1996), .B(G32), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(G33), .B(G2072), .ZN(n909) );
  NOR2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n916) );
  XOR2_X1 U1012 ( .A(G2067), .B(G26), .Z(n911) );
  NAND2_X1 U1013 ( .A1(n911), .A2(G28), .ZN(n914) );
  XNOR2_X1 U1014 ( .A(G25), .B(G1991), .ZN(n912) );
  XNOR2_X1 U1015 ( .A(KEYINPUT116), .B(n912), .ZN(n913) );
  NOR2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(G27), .B(n917), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1020 ( .A(KEYINPUT53), .B(n920), .Z(n923) );
  XOR2_X1 U1021 ( .A(KEYINPUT54), .B(G34), .Z(n921) );
  XNOR2_X1 U1022 ( .A(G2084), .B(n921), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(G35), .B(G2090), .ZN(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1026 ( .A(KEYINPUT117), .B(n926), .Z(n927) );
  NOR2_X1 U1027 ( .A1(G29), .A2(n927), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(KEYINPUT55), .B(n928), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n929), .A2(G11), .ZN(n988) );
  INV_X1 U1030 ( .A(n930), .ZN(n932) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n954) );
  XNOR2_X1 U1032 ( .A(G164), .B(G2078), .ZN(n936) );
  XOR2_X1 U1033 ( .A(G2072), .B(n933), .Z(n934) );
  XNOR2_X1 U1034 ( .A(KEYINPUT115), .B(n934), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(n937), .B(KEYINPUT50), .ZN(n952) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n943) );
  XOR2_X1 U1038 ( .A(G160), .B(G2084), .Z(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n950) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n947) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1044 ( .A(KEYINPUT51), .B(n948), .Z(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(n955), .B(KEYINPUT52), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n956), .A2(G29), .ZN(n986) );
  XNOR2_X1 U1050 ( .A(G16), .B(KEYINPUT56), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT118), .ZN(n984) );
  XNOR2_X1 U1052 ( .A(G1348), .B(n958), .ZN(n963) );
  XOR2_X1 U1053 ( .A(G168), .B(G1966), .Z(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1055 ( .A(KEYINPUT57), .B(n961), .Z(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G1961), .B(G301), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n982) );
  XOR2_X1 U1059 ( .A(G1971), .B(G166), .Z(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n978) );
  XNOR2_X1 U1061 ( .A(n969), .B(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n970), .B(KEYINPUT119), .ZN(n973) );
  XOR2_X1 U1063 ( .A(n971), .B(KEYINPUT120), .Z(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(G1341), .B(n974), .ZN(n975) );
  NOR2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1069 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1071 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1072 ( .A1(n988), .A2(n987), .ZN(n1017) );
  XOR2_X1 U1073 ( .A(G1961), .B(G5), .Z(n1004) );
  XOR2_X1 U1074 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n999) );
  XOR2_X1 U1075 ( .A(KEYINPUT122), .B(G4), .Z(n990) );
  XNOR2_X1 U1076 ( .A(G1348), .B(KEYINPUT59), .ZN(n989) );
  XNOR2_X1 U1077 ( .A(n990), .B(n989), .ZN(n993) );
  XOR2_X1 U1078 ( .A(KEYINPUT121), .B(G1956), .Z(n991) );
  XNOR2_X1 U1079 ( .A(G20), .B(n991), .ZN(n992) );
  NOR2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n997) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(G1981), .B(G6), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(n999), .B(n998), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G21), .B(G1966), .ZN(n1000) );
  NOR2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(KEYINPUT124), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1011) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G22), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G23), .B(G1976), .ZN(n1005) );
  NOR2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XOR2_X1 U1093 ( .A(G1986), .B(G24), .Z(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(n1012), .B(KEYINPUT61), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(n1013), .B(KEYINPUT125), .ZN(n1014) );
  NOR2_X1 U1099 ( .A1(G16), .A2(n1014), .ZN(n1015) );
  XOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1015), .Z(n1016) );
  NAND2_X1 U1101 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

