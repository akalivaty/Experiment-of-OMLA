

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765;

  XNOR2_X1 U373 ( .A(n608), .B(n416), .ZN(n721) );
  NOR2_X1 U374 ( .A1(n607), .A2(n675), .ZN(n608) );
  NOR2_X2 U375 ( .A1(G953), .A2(G237), .ZN(n494) );
  NOR2_X1 U376 ( .A1(n681), .A2(n682), .ZN(n394) );
  INV_X1 U377 ( .A(G953), .ZN(n757) );
  XNOR2_X2 U378 ( .A(n404), .B(n403), .ZN(n764) );
  NOR2_X2 U379 ( .A1(n702), .A2(n355), .ZN(n703) );
  XNOR2_X2 U380 ( .A(KEYINPUT67), .B(KEYINPUT4), .ZN(n393) );
  NOR2_X1 U381 ( .A1(n406), .A2(n726), .ZN(n584) );
  INV_X1 U382 ( .A(KEYINPUT101), .ZN(n410) );
  AND2_X1 U383 ( .A1(n632), .A2(n436), .ZN(n384) );
  XNOR2_X1 U384 ( .A(n617), .B(KEYINPUT103), .ZN(n618) );
  NAND2_X1 U385 ( .A1(n616), .A2(n706), .ZN(n617) );
  XNOR2_X1 U386 ( .A(n411), .B(n410), .ZN(n616) );
  AND2_X1 U387 ( .A1(n369), .A2(n368), .ZN(n367) );
  OR2_X1 U388 ( .A1(n553), .A2(n696), .ZN(n404) );
  XNOR2_X1 U389 ( .A(n400), .B(n399), .ZN(n697) );
  XNOR2_X1 U390 ( .A(n468), .B(KEYINPUT100), .ZN(n562) );
  AND2_X1 U391 ( .A1(n431), .A2(n429), .ZN(n428) );
  XNOR2_X1 U392 ( .A(G119), .B(G116), .ZN(n482) );
  XNOR2_X1 U393 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n473) );
  NAND2_X2 U394 ( .A1(n426), .A2(n390), .ZN(n351) );
  BUF_X1 U395 ( .A(n409), .Z(n352) );
  NAND2_X1 U396 ( .A1(n426), .A2(n390), .ZN(n728) );
  XNOR2_X1 U397 ( .A(n370), .B(n402), .ZN(n409) );
  XNOR2_X1 U398 ( .A(n375), .B(KEYINPUT0), .ZN(n598) );
  XNOR2_X2 U399 ( .A(n499), .B(n438), .ZN(n741) );
  INV_X1 U400 ( .A(G902), .ZN(n534) );
  XNOR2_X1 U401 ( .A(n606), .B(KEYINPUT104), .ZN(n595) );
  NOR2_X1 U402 ( .A1(n422), .A2(n420), .ZN(n408) );
  NAND2_X1 U403 ( .A1(n421), .A2(n571), .ZN(n420) );
  NAND2_X1 U404 ( .A1(n424), .A2(n423), .ZN(n422) );
  NAND2_X1 U405 ( .A1(n676), .A2(n353), .ZN(n682) );
  XNOR2_X1 U406 ( .A(n425), .B(n503), .ZN(n606) );
  XNOR2_X1 U407 ( .A(n612), .B(n396), .ZN(n395) );
  INV_X1 U408 ( .A(KEYINPUT78), .ZN(n396) );
  XNOR2_X1 U409 ( .A(KEYINPUT48), .B(KEYINPUT68), .ZN(n573) );
  XNOR2_X1 U410 ( .A(G143), .B(G128), .ZN(n470) );
  XNOR2_X1 U411 ( .A(n551), .B(n552), .ZN(n666) );
  NOR2_X1 U412 ( .A1(n430), .A2(n492), .ZN(n429) );
  XNOR2_X1 U413 ( .A(n519), .B(n518), .ZN(n676) );
  INV_X1 U414 ( .A(KEYINPUT83), .ZN(n483) );
  XNOR2_X1 U415 ( .A(G122), .B(G134), .ZN(n445) );
  XNOR2_X1 U416 ( .A(n405), .B(KEYINPUT41), .ZN(n696) );
  NOR2_X1 U417 ( .A1(n670), .A2(n669), .ZN(n405) );
  XNOR2_X1 U418 ( .A(n600), .B(n599), .ZN(n373) );
  OR2_X1 U419 ( .A1(n697), .A2(n607), .ZN(n600) );
  NOR2_X1 U420 ( .A1(n681), .A2(n398), .ZN(n397) );
  INV_X1 U421 ( .A(n611), .ZN(n398) );
  XNOR2_X1 U422 ( .A(n554), .B(n386), .ZN(n385) );
  XNOR2_X1 U423 ( .A(n679), .B(n541), .ZN(n612) );
  NAND2_X1 U424 ( .A1(n351), .A2(G475), .ZN(n379) );
  NAND2_X1 U425 ( .A1(n366), .A2(n365), .ZN(n364) );
  NOR2_X1 U426 ( .A1(n417), .A2(KEYINPUT105), .ZN(n365) );
  NAND2_X1 U427 ( .A1(n763), .A2(KEYINPUT46), .ZN(n421) );
  INV_X1 U428 ( .A(n721), .ZN(n415) );
  NAND2_X1 U429 ( .A1(G234), .A2(G237), .ZN(n504) );
  INV_X1 U430 ( .A(G237), .ZN(n488) );
  NAND2_X1 U431 ( .A1(n490), .A2(n436), .ZN(n434) );
  NAND2_X1 U432 ( .A1(n433), .A2(n633), .ZN(n432) );
  INV_X1 U433 ( .A(n490), .ZN(n433) );
  NAND2_X1 U434 ( .A1(n584), .A2(n761), .ZN(n660) );
  XNOR2_X1 U435 ( .A(n393), .B(KEYINPUT64), .ZN(n392) );
  INV_X1 U436 ( .A(G146), .ZN(n452) );
  XNOR2_X1 U437 ( .A(n441), .B(n387), .ZN(n508) );
  INV_X1 U438 ( .A(KEYINPUT8), .ZN(n387) );
  XOR2_X1 U439 ( .A(KEYINPUT93), .B(KEYINPUT12), .Z(n455) );
  XNOR2_X1 U440 ( .A(G113), .B(G122), .ZN(n457) );
  XOR2_X1 U441 ( .A(KEYINPUT94), .B(G131), .Z(n458) );
  XOR2_X1 U442 ( .A(G143), .B(G104), .Z(n459) );
  XNOR2_X1 U443 ( .A(n401), .B(n493), .ZN(n529) );
  INV_X1 U444 ( .A(G131), .ZN(n493) );
  XNOR2_X1 U445 ( .A(G137), .B(G134), .ZN(n401) );
  XNOR2_X1 U446 ( .A(KEYINPUT18), .B(KEYINPUT85), .ZN(n478) );
  XNOR2_X1 U447 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n479) );
  AND2_X1 U448 ( .A1(n584), .A2(n583), .ZN(n661) );
  INV_X1 U449 ( .A(KEYINPUT30), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n466), .B(n465), .ZN(n565) );
  BUF_X1 U451 ( .A(n660), .Z(n755) );
  XNOR2_X1 U452 ( .A(G104), .B(G110), .ZN(n472) );
  NAND2_X1 U453 ( .A1(n508), .A2(G221), .ZN(n510) );
  XNOR2_X1 U454 ( .A(G128), .B(G110), .ZN(n511) );
  XOR2_X1 U455 ( .A(G146), .B(G140), .Z(n527) );
  XNOR2_X1 U456 ( .A(n529), .B(KEYINPUT90), .ZN(n750) );
  INV_X1 U457 ( .A(KEYINPUT33), .ZN(n399) );
  NAND2_X1 U458 ( .A1(n394), .A2(n612), .ZN(n400) );
  NAND2_X1 U459 ( .A1(n662), .A2(n661), .ZN(n380) );
  INV_X1 U460 ( .A(KEYINPUT39), .ZN(n560) );
  XNOR2_X1 U461 ( .A(n544), .B(KEYINPUT107), .ZN(n574) );
  AND2_X1 U462 ( .A1(n542), .A2(n612), .ZN(n543) );
  INV_X1 U463 ( .A(n551), .ZN(n578) );
  NAND2_X1 U464 ( .A1(n597), .A2(n611), .ZN(n417) );
  NAND2_X1 U465 ( .A1(n417), .A2(KEYINPUT105), .ZN(n368) );
  INV_X1 U466 ( .A(n555), .ZN(n389) );
  BUF_X1 U467 ( .A(n606), .Z(n679) );
  XOR2_X1 U468 ( .A(KEYINPUT16), .B(G122), .Z(n438) );
  XNOR2_X1 U469 ( .A(n449), .B(n448), .ZN(n729) );
  XNOR2_X1 U470 ( .A(n447), .B(n439), .ZN(n448) );
  INV_X1 U471 ( .A(KEYINPUT42), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n372), .B(n604), .ZN(n762) );
  INV_X1 U473 ( .A(KEYINPUT32), .ZN(n402) );
  INV_X1 U474 ( .A(KEYINPUT60), .ZN(n376) );
  NAND2_X1 U475 ( .A1(n378), .A2(n644), .ZN(n377) );
  XNOR2_X1 U476 ( .A(n379), .B(n359), .ZN(n378) );
  INV_X1 U477 ( .A(KEYINPUT56), .ZN(n381) );
  INV_X1 U478 ( .A(G110), .ZN(n362) );
  XOR2_X1 U479 ( .A(n522), .B(n521), .Z(n353) );
  NAND2_X1 U480 ( .A1(n593), .A2(n353), .ZN(n354) );
  AND2_X1 U481 ( .A1(n380), .A2(KEYINPUT2), .ZN(n355) );
  NAND2_X1 U482 ( .A1(n397), .A2(n395), .ZN(n356) );
  XOR2_X1 U483 ( .A(n594), .B(KEYINPUT22), .Z(n357) );
  XNOR2_X1 U484 ( .A(KEYINPUT15), .B(G902), .ZN(n633) );
  XOR2_X1 U485 ( .A(n642), .B(n641), .Z(n358) );
  XOR2_X1 U486 ( .A(n655), .B(n654), .Z(n359) );
  XOR2_X1 U487 ( .A(n657), .B(n658), .Z(n360) );
  AND2_X1 U488 ( .A1(n436), .A2(KEYINPUT2), .ZN(n361) );
  INV_X1 U489 ( .A(n363), .ZN(n371) );
  XNOR2_X1 U490 ( .A(n363), .B(n362), .ZN(G12) );
  NAND2_X1 U491 ( .A1(n367), .A2(n364), .ZN(n363) );
  INV_X1 U492 ( .A(n615), .ZN(n366) );
  NAND2_X1 U493 ( .A1(n615), .A2(KEYINPUT105), .ZN(n369) );
  NAND2_X1 U494 ( .A1(n371), .A2(n409), .ZN(n374) );
  NOR2_X2 U495 ( .A1(n615), .A2(n356), .ZN(n370) );
  XNOR2_X1 U496 ( .A(n377), .B(n376), .ZN(G60) );
  OR2_X2 U497 ( .A1(n623), .A2(n762), .ZN(n605) );
  NAND2_X1 U498 ( .A1(n373), .A2(n602), .ZN(n372) );
  XNOR2_X1 U499 ( .A(n374), .B(KEYINPUT82), .ZN(n623) );
  NAND2_X1 U500 ( .A1(n592), .A2(n591), .ZN(n375) );
  XNOR2_X2 U501 ( .A(n545), .B(KEYINPUT19), .ZN(n592) );
  NAND2_X2 U502 ( .A1(n428), .A2(n435), .ZN(n545) );
  NAND2_X1 U503 ( .A1(n380), .A2(n361), .ZN(n426) );
  XNOR2_X1 U504 ( .A(n382), .B(n381), .ZN(G51) );
  NAND2_X1 U505 ( .A1(n383), .A2(n644), .ZN(n382) );
  XNOR2_X1 U506 ( .A(n659), .B(n360), .ZN(n383) );
  XNOR2_X1 U507 ( .A(n501), .B(n502), .ZN(n649) );
  NAND2_X1 U508 ( .A1(n384), .A2(n631), .ZN(n390) );
  XNOR2_X1 U509 ( .A(n407), .B(n573), .ZN(n406) );
  NOR2_X1 U510 ( .A1(n567), .A2(n559), .ZN(n561) );
  NAND2_X1 U511 ( .A1(n557), .A2(n385), .ZN(n558) );
  NAND2_X1 U512 ( .A1(n389), .A2(n388), .ZN(n609) );
  INV_X1 U513 ( .A(n682), .ZN(n388) );
  NOR2_X1 U514 ( .A1(n734), .A2(n661), .ZN(n631) );
  XNOR2_X2 U515 ( .A(n630), .B(n629), .ZN(n734) );
  XNOR2_X2 U516 ( .A(n391), .B(n357), .ZN(n615) );
  NOR2_X2 U517 ( .A1(n598), .A2(n354), .ZN(n391) );
  XNOR2_X2 U518 ( .A(n392), .B(n470), .ZN(n749) );
  NAND2_X1 U519 ( .A1(n394), .A2(n679), .ZN(n675) );
  XNOR2_X2 U520 ( .A(n555), .B(KEYINPUT1), .ZN(n681) );
  XNOR2_X1 U521 ( .A(n352), .B(G119), .ZN(G21) );
  NAND2_X1 U522 ( .A1(n572), .A2(n408), .ZN(n407) );
  NAND2_X1 U523 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U524 ( .A(n671), .ZN(n412) );
  NAND2_X1 U525 ( .A1(n415), .A2(n414), .ZN(n413) );
  INV_X1 U526 ( .A(n709), .ZN(n414) );
  INV_X1 U527 ( .A(KEYINPUT31), .ZN(n416) );
  NAND2_X1 U528 ( .A1(n419), .A2(n418), .ZN(n424) );
  NOR2_X1 U529 ( .A1(n764), .A2(KEYINPUT46), .ZN(n418) );
  INV_X1 U530 ( .A(n763), .ZN(n419) );
  XNOR2_X2 U531 ( .A(n564), .B(n563), .ZN(n763) );
  NAND2_X1 U532 ( .A1(n764), .A2(KEYINPUT46), .ZN(n423) );
  NAND2_X1 U533 ( .A1(n595), .A2(n665), .ZN(n554) );
  NAND2_X1 U534 ( .A1(n649), .A2(n534), .ZN(n425) );
  NAND2_X1 U535 ( .A1(n427), .A2(n435), .ZN(n551) );
  AND2_X1 U536 ( .A1(n431), .A2(n434), .ZN(n427) );
  INV_X1 U537 ( .A(n434), .ZN(n430) );
  OR2_X2 U538 ( .A1(n656), .A2(n432), .ZN(n431) );
  NAND2_X1 U539 ( .A1(n656), .A2(n490), .ZN(n435) );
  INV_X1 U540 ( .A(n633), .ZN(n436) );
  XNOR2_X1 U541 ( .A(KEYINPUT110), .B(KEYINPUT36), .ZN(n437) );
  XOR2_X1 U542 ( .A(n446), .B(n445), .Z(n439) );
  NAND2_X1 U543 ( .A1(n707), .A2(n543), .ZN(n544) );
  INV_X1 U544 ( .A(n733), .ZN(n644) );
  INV_X1 U545 ( .A(KEYINPUT124), .ZN(n638) );
  XOR2_X1 U546 ( .A(KEYINPUT7), .B(KEYINPUT98), .Z(n443) );
  INV_X1 U547 ( .A(G953), .ZN(n440) );
  NAND2_X1 U548 ( .A1(G234), .A2(n440), .ZN(n441) );
  NAND2_X1 U549 ( .A1(G217), .A2(n508), .ZN(n442) );
  XNOR2_X1 U550 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U551 ( .A(n444), .B(G116), .Z(n449) );
  XOR2_X1 U552 ( .A(G107), .B(n470), .Z(n447) );
  XOR2_X1 U553 ( .A(KEYINPUT9), .B(KEYINPUT97), .Z(n446) );
  NOR2_X1 U554 ( .A1(G902), .A2(n729), .ZN(n451) );
  XNOR2_X1 U555 ( .A(KEYINPUT99), .B(G478), .ZN(n450) );
  XNOR2_X1 U556 ( .A(n451), .B(n450), .ZN(n566) );
  XNOR2_X1 U557 ( .A(n452), .B(G125), .ZN(n477) );
  XNOR2_X1 U558 ( .A(n477), .B(G140), .ZN(n453) );
  XNOR2_X1 U559 ( .A(n453), .B(KEYINPUT10), .ZN(n748) );
  NAND2_X1 U560 ( .A1(n494), .A2(G214), .ZN(n454) );
  XNOR2_X1 U561 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U562 ( .A(n456), .B(KEYINPUT11), .Z(n462) );
  XNOR2_X1 U563 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U564 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U565 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U566 ( .A(n463), .B(n748), .ZN(n655) );
  NAND2_X1 U567 ( .A1(n655), .A2(n534), .ZN(n466) );
  XOR2_X1 U568 ( .A(G475), .B(KEYINPUT95), .Z(n464) );
  XOR2_X1 U569 ( .A(KEYINPUT13), .B(n464), .Z(n465) );
  XOR2_X1 U570 ( .A(n565), .B(KEYINPUT96), .Z(n467) );
  AND2_X1 U571 ( .A1(n566), .A2(n467), .ZN(n720) );
  NOR2_X1 U572 ( .A1(n467), .A2(n566), .ZN(n468) );
  NOR2_X1 U573 ( .A1(n720), .A2(n562), .ZN(n671) );
  NAND2_X1 U574 ( .A1(n671), .A2(KEYINPUT47), .ZN(n469) );
  XNOR2_X1 U575 ( .A(n469), .B(KEYINPUT80), .ZN(n540) );
  INV_X1 U576 ( .A(G101), .ZN(n471) );
  XNOR2_X2 U577 ( .A(n749), .B(n471), .ZN(n501) );
  XNOR2_X1 U578 ( .A(n472), .B(G107), .ZN(n742) );
  XNOR2_X1 U579 ( .A(n742), .B(n473), .ZN(n474) );
  XNOR2_X2 U580 ( .A(n501), .B(n474), .ZN(n533) );
  NAND2_X1 U581 ( .A1(n757), .A2(G224), .ZN(n475) );
  XNOR2_X1 U582 ( .A(n475), .B(KEYINPUT76), .ZN(n476) );
  XNOR2_X1 U583 ( .A(n477), .B(n476), .ZN(n481) );
  XNOR2_X1 U584 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n481), .B(n480), .ZN(n486) );
  XNOR2_X1 U586 ( .A(n482), .B(KEYINPUT3), .ZN(n485) );
  XNOR2_X1 U587 ( .A(n483), .B(G113), .ZN(n484) );
  XNOR2_X2 U588 ( .A(n485), .B(n484), .ZN(n499) );
  XNOR2_X1 U589 ( .A(n486), .B(n741), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n533), .B(n487), .ZN(n656) );
  NAND2_X1 U591 ( .A1(n534), .A2(n488), .ZN(n491) );
  NAND2_X1 U592 ( .A1(n491), .A2(G210), .ZN(n489) );
  XNOR2_X1 U593 ( .A(n489), .B(KEYINPUT86), .ZN(n490) );
  NAND2_X1 U594 ( .A1(n491), .A2(G214), .ZN(n665) );
  INV_X1 U595 ( .A(n665), .ZN(n492) );
  XOR2_X1 U596 ( .A(KEYINPUT108), .B(KEYINPUT28), .Z(n525) );
  INV_X1 U597 ( .A(n529), .ZN(n498) );
  XOR2_X1 U598 ( .A(G146), .B(KEYINPUT5), .Z(n496) );
  NAND2_X1 U599 ( .A1(n494), .A2(G210), .ZN(n495) );
  XNOR2_X1 U600 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U602 ( .A(n500), .B(n499), .ZN(n502) );
  XNOR2_X1 U603 ( .A(KEYINPUT92), .B(G472), .ZN(n503) );
  XNOR2_X1 U604 ( .A(n504), .B(KEYINPUT14), .ZN(n505) );
  AND2_X1 U605 ( .A1(n505), .A2(G952), .ZN(n694) );
  AND2_X1 U606 ( .A1(n694), .A2(n757), .ZN(n589) );
  NAND2_X1 U607 ( .A1(G902), .A2(n505), .ZN(n586) );
  OR2_X1 U608 ( .A1(n757), .A2(n586), .ZN(n506) );
  NOR2_X1 U609 ( .A1(G900), .A2(n506), .ZN(n507) );
  NOR2_X1 U610 ( .A1(n589), .A2(n507), .ZN(n556) );
  XOR2_X1 U611 ( .A(G137), .B(KEYINPUT24), .Z(n509) );
  XNOR2_X1 U612 ( .A(n510), .B(n509), .ZN(n514) );
  XOR2_X1 U613 ( .A(KEYINPUT23), .B(G119), .Z(n512) );
  XNOR2_X1 U614 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U615 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U616 ( .A(n515), .B(n748), .ZN(n634) );
  NAND2_X1 U617 ( .A1(n634), .A2(n534), .ZN(n519) );
  NAND2_X1 U618 ( .A1(G234), .A2(n633), .ZN(n516) );
  XNOR2_X1 U619 ( .A(KEYINPUT20), .B(n516), .ZN(n520) );
  AND2_X1 U620 ( .A1(G217), .A2(n520), .ZN(n517) );
  XNOR2_X1 U621 ( .A(KEYINPUT25), .B(n517), .ZN(n518) );
  NOR2_X1 U622 ( .A1(n556), .A2(n676), .ZN(n523) );
  AND2_X1 U623 ( .A1(n520), .A2(G221), .ZN(n522) );
  INV_X1 U624 ( .A(KEYINPUT21), .ZN(n521) );
  AND2_X1 U625 ( .A1(n523), .A2(n353), .ZN(n542) );
  NAND2_X1 U626 ( .A1(n595), .A2(n542), .ZN(n524) );
  XOR2_X1 U627 ( .A(n525), .B(n524), .Z(n537) );
  NAND2_X1 U628 ( .A1(G227), .A2(n757), .ZN(n526) );
  XNOR2_X1 U629 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U630 ( .A(n528), .B(KEYINPUT91), .Z(n531) );
  XNOR2_X1 U631 ( .A(n750), .B(KEYINPUT75), .ZN(n530) );
  XNOR2_X1 U632 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U633 ( .A(n533), .B(n532), .ZN(n642) );
  NAND2_X1 U634 ( .A1(n642), .A2(n534), .ZN(n536) );
  XNOR2_X1 U635 ( .A(KEYINPUT69), .B(G469), .ZN(n535) );
  XNOR2_X2 U636 ( .A(n536), .B(n535), .ZN(n555) );
  NOR2_X1 U637 ( .A1(n537), .A2(n555), .ZN(n550) );
  AND2_X1 U638 ( .A1(n592), .A2(n550), .ZN(n716) );
  INV_X1 U639 ( .A(n716), .ZN(n538) );
  NAND2_X1 U640 ( .A1(n538), .A2(KEYINPUT47), .ZN(n539) );
  NAND2_X1 U641 ( .A1(n540), .A2(n539), .ZN(n549) );
  XNOR2_X1 U642 ( .A(n562), .B(KEYINPUT106), .ZN(n707) );
  XOR2_X1 U643 ( .A(KEYINPUT102), .B(KEYINPUT6), .Z(n541) );
  INV_X1 U644 ( .A(n545), .ZN(n546) );
  NAND2_X1 U645 ( .A1(n574), .A2(n546), .ZN(n547) );
  XNOR2_X1 U646 ( .A(n547), .B(n437), .ZN(n548) );
  NOR2_X1 U647 ( .A1(n548), .A2(n681), .ZN(n724) );
  NOR2_X1 U648 ( .A1(n549), .A2(n724), .ZN(n572) );
  INV_X1 U649 ( .A(n550), .ZN(n553) );
  OR2_X1 U650 ( .A1(n566), .A2(n565), .ZN(n669) );
  XNOR2_X1 U651 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n552) );
  NAND2_X1 U652 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U653 ( .A1(n609), .A2(n556), .ZN(n557) );
  XNOR2_X1 U654 ( .A(n558), .B(KEYINPUT74), .ZN(n567) );
  INV_X1 U655 ( .A(n666), .ZN(n559) );
  XNOR2_X1 U656 ( .A(n561), .B(n560), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n580), .A2(n562), .ZN(n564) );
  XNOR2_X1 U658 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n563) );
  NAND2_X1 U659 ( .A1(n566), .A2(n565), .ZN(n601) );
  NOR2_X1 U660 ( .A1(n567), .A2(n601), .ZN(n568) );
  NAND2_X1 U661 ( .A1(n568), .A2(n578), .ZN(n647) );
  NOR2_X1 U662 ( .A1(KEYINPUT47), .A2(n671), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n716), .A2(n569), .ZN(n570) );
  AND2_X1 U664 ( .A1(n647), .A2(n570), .ZN(n571) );
  INV_X1 U665 ( .A(n681), .ZN(n576) );
  NAND2_X1 U666 ( .A1(n574), .A2(n665), .ZN(n575) );
  NOR2_X1 U667 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U668 ( .A(n577), .B(KEYINPUT43), .ZN(n579) );
  NOR2_X1 U669 ( .A1(n579), .A2(n578), .ZN(n726) );
  AND2_X1 U670 ( .A1(n720), .A2(n580), .ZN(n581) );
  XNOR2_X1 U671 ( .A(n581), .B(KEYINPUT111), .ZN(n761) );
  XNOR2_X1 U672 ( .A(n660), .B(KEYINPUT73), .ZN(n632) );
  NAND2_X1 U673 ( .A1(n761), .A2(KEYINPUT2), .ZN(n582) );
  XNOR2_X1 U674 ( .A(n582), .B(KEYINPUT79), .ZN(n583) );
  NOR2_X1 U675 ( .A1(G898), .A2(n757), .ZN(n585) );
  XNOR2_X1 U676 ( .A(KEYINPUT87), .B(n585), .ZN(n744) );
  NOR2_X1 U677 ( .A1(n586), .A2(n744), .ZN(n587) );
  XNOR2_X1 U678 ( .A(n587), .B(KEYINPUT88), .ZN(n588) );
  NOR2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U680 ( .A(n590), .B(KEYINPUT89), .ZN(n591) );
  INV_X1 U681 ( .A(n669), .ZN(n593) );
  INV_X1 U682 ( .A(KEYINPUT65), .ZN(n594) );
  INV_X1 U683 ( .A(n595), .ZN(n596) );
  AND2_X1 U684 ( .A1(n681), .A2(n596), .ZN(n597) );
  INV_X1 U685 ( .A(n676), .ZN(n611) );
  BUF_X1 U686 ( .A(n598), .Z(n607) );
  INV_X1 U687 ( .A(KEYINPUT34), .ZN(n599) );
  INV_X1 U688 ( .A(n601), .ZN(n602) );
  INV_X1 U689 ( .A(KEYINPUT77), .ZN(n603) );
  XNOR2_X1 U690 ( .A(n603), .B(KEYINPUT35), .ZN(n604) );
  NAND2_X1 U691 ( .A1(n605), .A2(KEYINPUT44), .ZN(n619) );
  OR2_X1 U692 ( .A1(n609), .A2(n679), .ZN(n610) );
  NOR2_X1 U693 ( .A1(n607), .A2(n610), .ZN(n709) );
  NOR2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U695 ( .A1(n681), .A2(n613), .ZN(n614) );
  OR2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n706) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U698 ( .A(n620), .B(KEYINPUT81), .ZN(n628) );
  OR2_X1 U699 ( .A1(n762), .A2(KEYINPUT44), .ZN(n622) );
  INV_X1 U700 ( .A(KEYINPUT66), .ZN(n621) );
  XNOR2_X1 U701 ( .A(n622), .B(n621), .ZN(n626) );
  BUF_X1 U702 ( .A(n623), .Z(n624) );
  INV_X1 U703 ( .A(n624), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n630) );
  INV_X1 U706 ( .A(KEYINPUT45), .ZN(n629) );
  INV_X1 U707 ( .A(n734), .ZN(n662) );
  NAND2_X1 U708 ( .A1(n728), .A2(G217), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n634), .B(n635), .ZN(n637) );
  INV_X1 U710 ( .A(G952), .ZN(n636) );
  AND2_X1 U711 ( .A1(n636), .A2(G953), .ZN(n733) );
  NAND2_X1 U712 ( .A1(n637), .A2(n644), .ZN(n639) );
  XNOR2_X1 U713 ( .A(n639), .B(n638), .ZN(G66) );
  NAND2_X1 U714 ( .A1(n351), .A2(G469), .ZN(n643) );
  XNOR2_X1 U715 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n640), .B(KEYINPUT58), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n643), .B(n358), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n646), .B(KEYINPUT121), .ZN(G54) );
  XNOR2_X1 U720 ( .A(n647), .B(G143), .ZN(G45) );
  NAND2_X1 U721 ( .A1(n728), .A2(G472), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U725 ( .A1(n652), .A2(n644), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n653), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U727 ( .A(KEYINPUT122), .B(KEYINPUT59), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n351), .A2(G210), .ZN(n659) );
  BUF_X1 U729 ( .A(n656), .Z(n657) );
  XOR2_X1 U730 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n658) );
  NOR2_X1 U731 ( .A1(n661), .A2(n755), .ZN(n664) );
  BUF_X1 U732 ( .A(n662), .Z(n663) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n701) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT118), .ZN(n668) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U739 ( .A1(n697), .A2(n674), .ZN(n692) );
  INV_X1 U740 ( .A(n675), .ZN(n687) );
  NOR2_X1 U741 ( .A1(n353), .A2(n676), .ZN(n677) );
  XOR2_X1 U742 ( .A(KEYINPUT49), .B(n677), .Z(n678) );
  NOR2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U744 ( .A(KEYINPUT116), .B(n680), .Z(n685) );
  AND2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U746 ( .A(KEYINPUT50), .B(n683), .ZN(n684) );
  NOR2_X1 U747 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U749 ( .A(KEYINPUT51), .B(n688), .Z(n689) );
  NOR2_X1 U750 ( .A1(n696), .A2(n689), .ZN(n690) );
  XOR2_X1 U751 ( .A(KEYINPUT117), .B(n690), .Z(n691) );
  NOR2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U753 ( .A(KEYINPUT52), .B(n693), .Z(n695) );
  AND2_X1 U754 ( .A1(n695), .A2(n694), .ZN(n699) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U757 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U758 ( .A(n703), .B(KEYINPUT119), .ZN(n704) );
  NOR2_X1 U759 ( .A1(n704), .A2(G953), .ZN(n705) );
  XNOR2_X1 U760 ( .A(n705), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U761 ( .A(G101), .B(n706), .ZN(G3) );
  BUF_X1 U762 ( .A(n707), .Z(n718) );
  NAND2_X1 U763 ( .A1(n718), .A2(n709), .ZN(n708) );
  XNOR2_X1 U764 ( .A(n708), .B(G104), .ZN(G6) );
  XOR2_X1 U765 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n711) );
  NAND2_X1 U766 ( .A1(n709), .A2(n720), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U768 ( .A(G107), .B(n712), .ZN(G9) );
  XOR2_X1 U769 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n714) );
  NAND2_X1 U770 ( .A1(n716), .A2(n720), .ZN(n713) );
  XNOR2_X1 U771 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U772 ( .A(G128), .B(n715), .Z(G30) );
  NAND2_X1 U773 ( .A1(n718), .A2(n716), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n717), .B(G146), .ZN(G48) );
  NAND2_X1 U775 ( .A1(n721), .A2(n718), .ZN(n719) );
  XNOR2_X1 U776 ( .A(n719), .B(G113), .ZN(G15) );
  NAND2_X1 U777 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n722), .B(KEYINPUT114), .ZN(n723) );
  XNOR2_X1 U779 ( .A(G116), .B(n723), .ZN(G18) );
  XNOR2_X1 U780 ( .A(n724), .B(G125), .ZN(n725) );
  XNOR2_X1 U781 ( .A(n725), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U782 ( .A(n726), .B(G140), .ZN(n727) );
  XNOR2_X1 U783 ( .A(n727), .B(KEYINPUT115), .ZN(G42) );
  NAND2_X1 U784 ( .A1(n351), .A2(G478), .ZN(n731) );
  XOR2_X1 U785 ( .A(n729), .B(KEYINPUT123), .Z(n730) );
  XNOR2_X1 U786 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U787 ( .A1(n733), .A2(n732), .ZN(G63) );
  BUF_X1 U788 ( .A(n734), .Z(n735) );
  NOR2_X1 U789 ( .A1(n735), .A2(G953), .ZN(n736) );
  XNOR2_X1 U790 ( .A(n736), .B(KEYINPUT125), .ZN(n740) );
  NAND2_X1 U791 ( .A1(G953), .A2(G224), .ZN(n737) );
  XNOR2_X1 U792 ( .A(KEYINPUT61), .B(n737), .ZN(n738) );
  NAND2_X1 U793 ( .A1(n738), .A2(G898), .ZN(n739) );
  NAND2_X1 U794 ( .A1(n740), .A2(n739), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n742), .B(G101), .ZN(n743) );
  XNOR2_X1 U796 ( .A(n741), .B(n743), .ZN(n745) );
  NAND2_X1 U797 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U798 ( .A(n747), .B(n746), .Z(G69) );
  XOR2_X1 U799 ( .A(KEYINPUT126), .B(n748), .Z(n752) );
  XNOR2_X1 U800 ( .A(n749), .B(n750), .ZN(n751) );
  XOR2_X1 U801 ( .A(n752), .B(n751), .Z(n756) );
  XNOR2_X1 U802 ( .A(G227), .B(n756), .ZN(n753) );
  NAND2_X1 U803 ( .A1(G900), .A2(n753), .ZN(n754) );
  NAND2_X1 U804 ( .A1(n754), .A2(G953), .ZN(n760) );
  XNOR2_X1 U805 ( .A(n756), .B(n755), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n760), .A2(n759), .ZN(G72) );
  XNOR2_X1 U808 ( .A(G134), .B(n761), .ZN(G36) );
  XOR2_X1 U809 ( .A(G122), .B(n762), .Z(G24) );
  XOR2_X1 U810 ( .A(n763), .B(G131), .Z(G33) );
  XNOR2_X1 U811 ( .A(G137), .B(KEYINPUT127), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n765), .B(n764), .ZN(G39) );
endmodule

