//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n449, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g035(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G101), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n462), .A2(G137), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n473), .B(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(new_n467), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n462), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n460), .A2(new_n461), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI221_X1 g059(.A(new_n479), .B1(new_n480), .B2(new_n481), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n467), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n484), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n471), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT3), .B1(KEYINPUT69), .B2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(KEYINPUT72), .B(new_n493), .C1(new_n496), .C2(new_n497), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n495), .B1(new_n502), .B2(KEYINPUT73), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT4), .A4(new_n501), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n490), .B1(new_n503), .B2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT74), .B(G651), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(G543), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n509), .B2(new_n510), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n518), .A2(new_n507), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n513), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n516), .A2(G89), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n512), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n514), .B(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(G63), .A3(G651), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n522), .A2(new_n523), .A3(new_n525), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  NAND2_X1  g105(.A1(new_n527), .A2(G64), .ZN(new_n531));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n507), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n511), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n514), .B(KEYINPUT75), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n507), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT76), .ZN(new_n544));
  AOI22_X1  g119(.A1(G43), .A2(new_n512), .B1(new_n516), .B2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(KEYINPUT76), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n511), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n511), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(KEYINPUT77), .A2(G78), .A3(G543), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n514), .A2(G65), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G651), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n562), .B2(new_n563), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n516), .A2(G91), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n557), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  NAND2_X1  g144(.A1(new_n520), .A2(KEYINPUT79), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT79), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n513), .A2(new_n517), .A3(new_n571), .A4(new_n519), .ZN(new_n572));
  AND2_X1   g147(.A1(new_n570), .A2(new_n572), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n574));
  OAI211_X1 g149(.A(G49), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n575));
  INV_X1    g150(.A(G87), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n515), .ZN(G288));
  OAI211_X1 g152(.A(G48), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n578));
  OAI211_X1 g153(.A(G86), .B(new_n514), .C1(new_n509), .C2(new_n510), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n514), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(new_n585), .A3(new_n542), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT80), .B1(new_n587), .B2(new_n507), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n580), .A2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n527), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n507), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n593), .A2(new_n511), .B1(new_n515), .B2(new_n594), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n592), .A2(KEYINPUT81), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT81), .B1(new_n592), .B2(new_n595), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n516), .A2(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n582), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n512), .A2(G54), .B1(G651), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n599), .B1(new_n608), .B2(G868), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  INV_X1    g186(.A(G299), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n608), .B1(new_n615), .B2(G860), .ZN(G148));
  OR3_X1    g191(.A1(new_n607), .A2(KEYINPUT82), .A3(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT82), .B1(new_n607), .B2(G559), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  OR3_X1    g195(.A1(new_n619), .A2(KEYINPUT83), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT83), .B1(new_n619), .B2(new_n620), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n621), .B(new_n622), .C1(G868), .C2(new_n548), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n462), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n467), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(G123), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n625), .B1(new_n626), .B2(new_n627), .C1(new_n628), .C2(new_n484), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT85), .Z(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n471), .A2(new_n464), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2100), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n630), .A2(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n648), .A2(new_n651), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT87), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n659), .B(KEYINPUT17), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n660), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n663), .B(new_n664), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n659), .A2(new_n656), .A3(new_n660), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n656), .A3(new_n667), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1961), .B(G1966), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(G229));
  NOR2_X1   g270(.A1(G6), .A2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G305), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT32), .ZN(new_n699));
  INV_X1    g274(.A(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G23), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT91), .Z(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(G288), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT33), .ZN(new_n706));
  INV_X1    g281(.A(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(G22), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT92), .Z(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G166), .B2(new_n704), .ZN(new_n711));
  INV_X1    g286(.A(G1971), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n701), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n714), .A2(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n704), .A2(G24), .ZN(new_n716));
  INV_X1    g291(.A(G290), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(new_n704), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(G1986), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(G1986), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n462), .A2(G131), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n467), .A2(G107), .ZN(new_n722));
  OAI21_X1  g297(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n723));
  INV_X1    g298(.A(G119), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n721), .B1(new_n722), .B2(new_n723), .C1(new_n724), .C2(new_n484), .ZN(new_n725));
  MUX2_X1   g300(.A(G25), .B(new_n725), .S(G29), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n719), .A2(new_n720), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n714), .A2(KEYINPUT93), .A3(KEYINPUT34), .ZN(new_n731));
  AOI21_X1  g306(.A(KEYINPUT93), .B1(new_n714), .B2(KEYINPUT34), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT36), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(KEYINPUT94), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n730), .B(new_n735), .C1(new_n731), .C2(new_n732), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n704), .A2(G20), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT23), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G299), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1956), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G35), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G162), .B2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT29), .B(G2090), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n548), .A2(new_n704), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n704), .B2(G19), .ZN(new_n750));
  INV_X1    g325(.A(G1341), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n744), .B(new_n752), .C1(new_n751), .C2(new_n750), .ZN(new_n753));
  OAI21_X1  g328(.A(KEYINPUT101), .B1(G29), .B2(G32), .ZN(new_n754));
  INV_X1    g329(.A(new_n484), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G129), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n462), .A2(G141), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n464), .ZN(new_n762));
  AND3_X1   g337(.A1(new_n756), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  MUX2_X1   g339(.A(KEYINPUT101), .B(new_n754), .S(new_n764), .Z(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT31), .B(G11), .Z(new_n768));
  INV_X1    g343(.A(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n769), .B2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  INV_X1    g348(.A(G29), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(G33), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT100), .B(KEYINPUT25), .Z(new_n776));
  NAND3_X1  g351(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n462), .A2(G139), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n778), .B(new_n779), .C1(new_n467), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(G29), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n767), .B(new_n772), .C1(new_n773), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n704), .A2(G5), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G171), .B2(new_n704), .ZN(new_n785));
  INV_X1    g360(.A(G1961), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n766), .B2(new_n765), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n704), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G168), .B2(new_n704), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1966), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n774), .B1(KEYINPUT24), .B2(G34), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(KEYINPUT24), .B2(G34), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n477), .B2(G29), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n782), .A2(new_n773), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n796), .B1(new_n792), .B2(new_n795), .C1(new_n774), .C2(new_n630), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n783), .A2(new_n788), .A3(new_n791), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n774), .A2(G27), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT102), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n801));
  AOI21_X1  g376(.A(KEYINPUT72), .B1(new_n483), .B2(new_n493), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT73), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n803), .A2(new_n505), .A3(new_n494), .ZN(new_n804));
  INV_X1    g379(.A(new_n490), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(G29), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2078), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n798), .A2(KEYINPUT103), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G4), .A2(G16), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n608), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT95), .ZN(new_n812));
  INV_X1    g387(.A(G1348), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n774), .A2(G26), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT28), .ZN(new_n816));
  NOR2_X1   g391(.A1(G104), .A2(G2105), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT96), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G116), .C2(new_n467), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT97), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n755), .A2(G128), .B1(G140), .B2(new_n462), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(KEYINPUT98), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n825), .A2(KEYINPUT99), .A3(G29), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT99), .B1(new_n825), .B2(G29), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n816), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(G2067), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n753), .A2(new_n809), .A3(new_n814), .A4(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT103), .B1(new_n798), .B2(new_n808), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n738), .A2(new_n739), .A3(new_n833), .ZN(G150));
  INV_X1    g409(.A(G150), .ZN(G311));
  NAND2_X1  g410(.A1(new_n608), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n527), .A2(G67), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n507), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n841), .A2(new_n511), .B1(new_n515), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n548), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n546), .B2(new_n547), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n837), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n844), .A2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(G145));
  INV_X1    g433(.A(new_n763), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n806), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n462), .A2(G142), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n467), .A2(KEYINPUT107), .A3(G118), .ZN(new_n862));
  OAI21_X1  g437(.A(KEYINPUT107), .B1(new_n467), .B2(G118), .ZN(new_n863));
  OR2_X1    g438(.A1(G106), .A2(G2105), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(G2104), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  OAI221_X1 g441(.A(new_n861), .B1(new_n862), .B2(new_n865), .C1(new_n866), .C2(new_n484), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n860), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n781), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT105), .Z(new_n872));
  OR2_X1    g447(.A1(new_n825), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n825), .A2(new_n872), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n725), .B(new_n634), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n873), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n873), .B2(new_n874), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n869), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n868), .A3(new_n877), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n630), .B(new_n477), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G162), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n884), .B1(new_n880), .B2(new_n882), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n888), .A2(KEYINPUT108), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n890));
  AOI211_X1 g465(.A(new_n890), .B(new_n884), .C1(new_n880), .C2(new_n882), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g468(.A1(new_n619), .A2(new_n849), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n849), .A2(new_n618), .A3(new_n617), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n607), .A2(G299), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n612), .A2(new_n602), .A3(new_n606), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(new_n898), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n894), .B2(new_n895), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT110), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n697), .B(new_n520), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n911));
  INV_X1    g486(.A(G288), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n717), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G290), .A2(G288), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(KEYINPUT109), .A3(new_n910), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(KEYINPUT109), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n911), .A2(new_n913), .A3(new_n917), .A4(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT42), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n905), .A2(new_n908), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT110), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n909), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NOR3_X1   g500(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n846), .A2(new_n620), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(G331));
  OAI21_X1  g505(.A(G286), .B1(G171), .B2(KEYINPUT111), .ZN(new_n931));
  NAND2_X1  g506(.A1(G171), .A2(KEYINPUT111), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n845), .A2(new_n847), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n845), .B2(new_n847), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n935), .ZN(new_n937));
  INV_X1    g512(.A(new_n931), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n933), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n936), .A2(new_n939), .A3(new_n907), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n903), .B1(new_n936), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n919), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n919), .B1(new_n940), .B2(new_n941), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT43), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n936), .A2(new_n939), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n904), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n936), .A2(new_n939), .A3(new_n907), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n901), .A2(KEYINPUT112), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT112), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n902), .B1(new_n952), .B2(new_n900), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n936), .A2(new_n939), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n919), .B1(new_n940), .B2(new_n954), .ZN(new_n955));
  AND4_X1   g530(.A1(KEYINPUT43), .A2(new_n950), .A3(new_n955), .A4(new_n886), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n946), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT43), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n944), .B2(new_n945), .ZN(new_n960));
  AND4_X1   g535(.A1(new_n959), .A2(new_n950), .A3(new_n955), .A4(new_n886), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(new_n962), .ZN(G397));
  AOI21_X1  g538(.A(KEYINPUT57), .B1(new_n557), .B2(KEYINPUT120), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(G299), .ZN(new_n965));
  OAI211_X1 g540(.A(G40), .B(new_n470), .C1(new_n476), .C2(new_n467), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(G1384), .B1(new_n804), .B2(new_n805), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(KEYINPUT45), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  XNOR2_X1  g545(.A(KEYINPUT113), .B(G1384), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n970), .B(new_n971), .C1(new_n804), .C2(new_n805), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT56), .B(G2072), .Z(new_n973));
  NOR3_X1   g548(.A1(new_n969), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n806), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n978), .A3(new_n967), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n974), .A2(KEYINPUT121), .B1(new_n743), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n970), .B1(G164), .B2(G1384), .ZN(new_n981));
  INV_X1    g556(.A(new_n971), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n806), .A2(KEYINPUT45), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n973), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n981), .A2(new_n967), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT121), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n965), .B1(new_n980), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n806), .A2(new_n977), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n966), .B1(new_n989), .B2(new_n970), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n990), .A2(KEYINPUT121), .A3(new_n983), .A4(new_n984), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n979), .A2(new_n743), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n965), .A2(new_n987), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n967), .B1(new_n968), .B2(new_n976), .ZN(new_n994));
  AOI211_X1 g569(.A(KEYINPUT50), .B(G1384), .C1(new_n804), .C2(new_n805), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n813), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g571(.A(G1384), .B(new_n966), .C1(new_n804), .C2(new_n805), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n829), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n607), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n988), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT61), .ZN(new_n1001));
  INV_X1    g576(.A(new_n993), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n988), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n987), .A2(new_n991), .A3(new_n992), .ZN(new_n1004));
  INV_X1    g579(.A(new_n965), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1006), .A2(KEYINPUT123), .A3(KEYINPUT61), .A4(new_n993), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n996), .A2(new_n998), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n607), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n996), .A2(new_n608), .A3(new_n998), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(KEYINPUT60), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1996), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n981), .A2(new_n1012), .A3(new_n967), .A4(new_n983), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT58), .B(G1341), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT122), .B1(new_n997), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n806), .A2(new_n977), .A3(new_n967), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT122), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1014), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1013), .A2(new_n1015), .A3(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1020), .A2(KEYINPUT59), .A3(new_n548), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT59), .B1(new_n1020), .B2(new_n548), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT60), .ZN(new_n1023));
  AND4_X1   g598(.A1(new_n1023), .A2(new_n996), .A3(new_n608), .A4(new_n998), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1003), .A2(new_n1007), .A3(new_n1011), .A4(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n988), .A2(new_n1002), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT123), .B1(new_n1027), .B2(KEYINPUT61), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1000), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n975), .A2(new_n792), .A3(new_n978), .A4(new_n967), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT118), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n966), .B1(new_n989), .B2(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n792), .A4(new_n978), .ZN(new_n1034));
  INV_X1    g609(.A(G1966), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n989), .A2(new_n970), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n969), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G8), .ZN(new_n1039));
  INV_X1    g614(.A(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G168), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT124), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1039), .B(new_n1042), .C1(new_n1043), .C2(KEYINPUT51), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT51), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1045));
  OAI211_X1 g620(.A(G8), .B(new_n1045), .C1(new_n1038), .C2(G286), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT49), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n580), .A2(new_n589), .A3(new_n700), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n700), .B1(new_n580), .B2(new_n589), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G305), .A2(G1981), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n580), .A2(new_n589), .A3(new_n700), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(KEYINPUT49), .A3(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1052), .A2(new_n1055), .A3(G8), .A4(new_n1016), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1016), .A2(G8), .ZN(new_n1057));
  NOR2_X1   g632(.A1(G288), .A2(new_n707), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT52), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1058), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n707), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(G8), .A4(new_n1016), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1056), .A2(new_n1059), .A3(KEYINPUT117), .A4(new_n1062), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n570), .A2(new_n572), .A3(G8), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G2090), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1032), .A2(new_n1070), .A3(new_n978), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n712), .B1(new_n969), .B2(new_n972), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1040), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1065), .A2(new_n1066), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G2078), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n981), .A2(new_n1075), .A3(new_n967), .A4(new_n983), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n470), .A2(KEYINPUT53), .A3(G40), .A4(new_n1075), .ZN(new_n1079));
  INV_X1    g654(.A(new_n476), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1080), .A2(KEYINPUT125), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n467), .B1(new_n1080), .B2(KEYINPUT125), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n983), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT45), .B1(new_n806), .B2(new_n982), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n979), .A2(new_n786), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1078), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G171), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1077), .A2(new_n1076), .B1(new_n979), .B2(new_n786), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1036), .A2(new_n969), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT53), .A3(new_n1075), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1092), .A3(G301), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(KEYINPUT54), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1069), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1071), .A2(new_n1096), .A3(new_n1072), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1096), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1074), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1088), .A2(G171), .ZN(new_n1103));
  AOI21_X1  g678(.A(G301), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT126), .B(new_n1102), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1101), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1029), .A2(new_n1048), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1048), .A2(KEYINPUT62), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1044), .A2(new_n1112), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1074), .A2(new_n1100), .A3(new_n1104), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1073), .A2(new_n1069), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G288), .A2(G1976), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1050), .B1(new_n1056), .B2(new_n1117), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1116), .A2(new_n1063), .B1(new_n1057), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1038), .A2(G8), .A3(G168), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT119), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1074), .A2(new_n1100), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1120), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1063), .A2(new_n1120), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(new_n1116), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT119), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1129));
  OAI221_X1 g704(.A(new_n1126), .B1(new_n1069), .B2(new_n1073), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1119), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1110), .A2(new_n1115), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1085), .A2(new_n967), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(G1996), .A3(new_n859), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT114), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n825), .B(new_n829), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(G1996), .B2(new_n859), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1136), .B1(new_n1138), .B2(new_n1134), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n725), .B(new_n727), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n1133), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(G290), .B(G1986), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1141), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1132), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1133), .B1(new_n1137), .B2(new_n763), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT46), .B1(new_n1133), .B2(G1996), .ZN(new_n1146));
  OR3_X1    g721(.A1(new_n1133), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT47), .ZN(new_n1149));
  NOR3_X1   g724(.A1(G290), .A2(new_n1133), .A3(G1986), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1151));
  XNOR2_X1  g726(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1141), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n727), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n725), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1139), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n823), .A2(new_n829), .A3(new_n824), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1133), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1149), .A2(new_n1153), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1144), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g735(.A(G319), .B1(new_n653), .B2(new_n654), .ZN(new_n1162));
  OR2_X1    g736(.A1(G227), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g737(.A(new_n1163), .B1(new_n693), .B2(new_n694), .ZN(new_n1164));
  OAI211_X1 g738(.A(new_n892), .B(new_n1164), .C1(new_n960), .C2(new_n961), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


