//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XOR2_X1   g001(.A(G15gat), .B(G43gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT28), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT27), .B1(new_n209), .B2(KEYINPUT69), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR3_X1   g011(.A1(new_n209), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n208), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT28), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221));
  OAI22_X1  g020(.A1(new_n220), .A2(new_n221), .B1(new_n209), .B2(new_n211), .ZN(new_n222));
  AND2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT26), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(G183gat), .A3(G190gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(G183gat), .B(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(new_n229), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n223), .B1(KEYINPUT23), .B2(new_n224), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT64), .B1(new_n220), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT64), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n224), .A2(new_n236), .A3(KEYINPUT23), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n232), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI211_X1 g039(.A(KEYINPUT65), .B(new_n233), .C1(new_n235), .C2(new_n237), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT25), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n209), .A2(G190gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n211), .A2(G183gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n229), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n230), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n249), .B(new_n230), .C1(new_n231), .C2(new_n229), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n220), .A2(KEYINPUT64), .A3(new_n234), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n236), .B1(new_n224), .B2(KEYINPUT23), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT23), .ZN(new_n256));
  NAND2_X1  g055(.A1(G169gat), .A2(G176gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n255), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n251), .A2(new_n262), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n242), .A2(new_n243), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n232), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n258), .B1(new_n254), .B2(new_n253), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(KEYINPUT65), .ZN(new_n267));
  INV_X1    g066(.A(new_n241), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n252), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n248), .A2(new_n250), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n255), .A2(new_n260), .A3(new_n261), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT68), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n228), .B1(new_n264), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G113gat), .ZN(new_n275));
  INV_X1    g074(.A(G120gat), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n275), .B2(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G127gat), .ZN(new_n280));
  INV_X1    g079(.A(G127gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G134gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n283), .B1(new_n280), .B2(new_n282), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n278), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n280), .A2(new_n282), .ZN(new_n287));
  XOR2_X1   g086(.A(KEYINPUT71), .B(G120gat), .Z(new_n288));
  OAI211_X1 g087(.A(new_n287), .B(new_n277), .C1(new_n288), .C2(new_n275), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n207), .B1(new_n274), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n243), .B1(new_n242), .B2(new_n263), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n269), .A2(KEYINPUT68), .A3(new_n272), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n227), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n286), .A4(new_n289), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n274), .A2(new_n290), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n291), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT33), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n206), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n303), .B1(new_n297), .B2(new_n299), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  AOI221_X4 g105(.A(new_n303), .B1(KEYINPUT33), .B2(new_n205), .C1(new_n297), .C2(new_n299), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n291), .A2(new_n296), .ZN(new_n309));
  NAND2_X1  g108(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n309), .A2(new_n298), .A3(new_n295), .A4(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(KEYINPUT73), .A2(KEYINPUT34), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n313), .B(new_n310), .C1(new_n297), .C2(new_n299), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n306), .A2(new_n308), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n306), .B2(new_n308), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n202), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n315), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT33), .B1(new_n297), .B2(new_n299), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n304), .A2(new_n321), .A3(new_n206), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n322), .B2(new_n307), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT36), .A3(new_n316), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT82), .ZN(new_n326));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT80), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G148gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT77), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G148gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n333), .A3(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(G141gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G148gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(G155gat), .ZN(new_n339));
  INV_X1    g138(.A(G162gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n338), .B1(new_n341), .B2(KEYINPUT2), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT76), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(G155gat), .B2(G162gat), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n343), .A2(new_n345), .A3(new_n338), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n330), .A2(G141gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n335), .A2(G148gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n337), .A2(new_n342), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(new_n286), .A3(new_n289), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT4), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT77), .B(G148gat), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n348), .B1(new_n354), .B2(G141gat), .ZN(new_n355));
  AND2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n356), .B1(new_n347), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n330), .A2(G141gat), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT2), .B1(new_n336), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n345), .A3(new_n338), .ZN(new_n361));
  OAI22_X1  g160(.A1(new_n355), .A2(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n362), .A2(KEYINPUT3), .B1(new_n286), .B2(new_n289), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT78), .B1(new_n351), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n337), .A2(new_n342), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n356), .B1(new_n341), .B2(new_n344), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n343), .A3(new_n367), .ZN(new_n368));
  AND4_X1   g167(.A1(KEYINPUT78), .A2(new_n366), .A3(new_n364), .A4(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT79), .B(new_n363), .C1(new_n365), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT78), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n372), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n366), .A2(new_n368), .A3(KEYINPUT78), .A4(new_n364), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT79), .B1(new_n375), .B2(new_n363), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n329), .B(new_n353), .C1(new_n371), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n290), .A2(new_n362), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n352), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n378), .B(KEYINPUT5), .C1(new_n380), .C2(new_n329), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n329), .B1(new_n352), .B2(new_n379), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT81), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n326), .B1(new_n377), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n376), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n370), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n388), .A2(new_n383), .A3(new_n329), .A4(new_n353), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT0), .ZN(new_n392));
  XNOR2_X1  g191(.A(G57gat), .B(G85gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n385), .A3(new_n326), .ZN(new_n396));
  AND4_X1   g195(.A1(KEYINPUT6), .A2(new_n390), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n377), .A2(new_n326), .A3(new_n385), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n389), .B2(new_n386), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT6), .B1(new_n399), .B2(new_n395), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n395), .B1(new_n390), .B2(new_n396), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT30), .ZN(new_n404));
  XNOR2_X1  g203(.A(G197gat), .B(G204gat), .ZN(new_n405));
  INV_X1    g204(.A(G211gat), .ZN(new_n406));
  INV_X1    g205(.A(G218gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(KEYINPUT22), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n410), .B(new_n405), .C1(KEYINPUT22), .C2(new_n408), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT74), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n238), .A2(new_n239), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n241), .A3(new_n265), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n418), .A2(new_n252), .B1(new_n271), .B2(new_n270), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(new_n227), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n269), .A2(new_n272), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(KEYINPUT74), .A3(new_n228), .ZN(new_n422));
  AND2_X1   g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n423), .A2(KEYINPUT29), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n423), .B(new_n228), .C1(new_n264), .C2(new_n273), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n415), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n422), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n423), .A2(new_n428), .B1(new_n274), .B2(new_n424), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(new_n415), .ZN(new_n430));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(G64gat), .B(G92gat), .ZN(new_n432));
  XOR2_X1   g231(.A(new_n431), .B(new_n432), .Z(new_n433));
  AOI21_X1  g232(.A(new_n404), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n425), .A2(new_n426), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n414), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n274), .A2(new_n424), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT74), .B1(new_n421), .B2(new_n228), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n416), .B(new_n227), .C1(new_n269), .C2(new_n272), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n423), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n440), .A3(new_n415), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n436), .A2(new_n441), .A3(new_n433), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(KEYINPUT30), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n436), .A2(new_n441), .ZN(new_n444));
  INV_X1    g243(.A(new_n433), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT75), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT75), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n447), .B(new_n433), .C1(new_n436), .C2(new_n441), .ZN(new_n448));
  OAI22_X1  g247(.A1(new_n434), .A2(new_n443), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT83), .B1(new_n403), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n444), .A2(new_n445), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n447), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n433), .B1(new_n436), .B2(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT75), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n430), .A2(new_n404), .A3(new_n433), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n442), .A2(KEYINPUT30), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n452), .A2(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n390), .A2(new_n395), .A3(new_n396), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n458), .B1(new_n461), .B2(new_n401), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n457), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n450), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT31), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(G50gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT29), .B1(new_n412), .B2(new_n413), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n364), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI211_X1 g271(.A(KEYINPUT86), .B(KEYINPUT29), .C1(new_n412), .C2(new_n413), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n362), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT29), .B1(new_n373), .B2(new_n374), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n474), .B(new_n476), .C1(new_n414), .C2(new_n477), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n414), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT29), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n409), .A2(KEYINPUT85), .A3(new_n411), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n480), .B(new_n481), .C1(new_n414), .C2(KEYINPUT85), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n351), .B1(new_n482), .B2(new_n364), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(new_n475), .B(KEYINPUT84), .Z(new_n485));
  OAI21_X1  g284(.A(new_n478), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G22gat), .ZN(new_n487));
  INV_X1    g286(.A(G22gat), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n478), .B(new_n488), .C1(new_n484), .C2(new_n485), .ZN(new_n489));
  AOI211_X1 g288(.A(KEYINPUT87), .B(new_n469), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n487), .A2(new_n489), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n468), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(KEYINPUT87), .A3(new_n489), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n462), .A2(KEYINPUT93), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n397), .A2(KEYINPUT93), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT91), .B1(new_n429), .B2(new_n415), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n414), .B2(new_n435), .ZN(new_n501));
  INV_X1    g300(.A(new_n429), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n414), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT37), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT92), .B(KEYINPUT38), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n451), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n508), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT37), .ZN(new_n512));
  OAI22_X1  g311(.A1(new_n453), .A2(new_n511), .B1(new_n430), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n513), .A2(new_n507), .B1(new_n430), .B2(new_n433), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n499), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n388), .A2(new_n353), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT88), .B(KEYINPUT39), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n328), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n352), .A2(new_n379), .A3(new_n329), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT39), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n520), .B2(new_n519), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n352), .B(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n387), .B2(new_n370), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n522), .B1(new_n525), .B2(new_n329), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n518), .A2(new_n394), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT90), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT40), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(KEYINPUT90), .A3(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n529), .A2(new_n459), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n496), .B1(new_n532), .B2(new_n449), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n465), .A2(new_n496), .B1(new_n515), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n323), .A2(new_n316), .A3(new_n495), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT35), .B1(new_n465), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n498), .B1(new_n462), .B2(KEYINPUT93), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT35), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n457), .A2(new_n538), .A3(new_n495), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n323), .A2(KEYINPUT94), .A3(new_n316), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT94), .B1(new_n323), .B2(new_n316), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n325), .A2(new_n534), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G71gat), .A2(G78gat), .ZN(new_n546));
  OR2_X1    g345(.A1(G71gat), .A2(G78gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT101), .B1(new_n550), .B2(G57gat), .ZN(new_n551));
  INV_X1    g350(.A(G57gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(G64gat), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n550), .A2(KEYINPUT101), .A3(G57gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n550), .A2(G57gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n552), .A2(G64gat), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT9), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(new_n546), .A3(new_n547), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT21), .ZN(new_n561));
  AND2_X1   g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n281), .ZN(new_n564));
  XNOR2_X1  g363(.A(G15gat), .B(G22gat), .ZN(new_n565));
  INV_X1    g364(.A(G1gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT16), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(KEYINPUT99), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n565), .A2(G1gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(KEYINPUT99), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT100), .B(G8gat), .Z(new_n573));
  NAND4_X1  g372(.A1(new_n569), .A2(new_n571), .A3(new_n572), .A4(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(G8gat), .B1(new_n568), .B2(new_n570), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(KEYINPUT21), .B2(new_n560), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n564), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n339), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n564), .A2(new_n577), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n564), .A2(new_n577), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n586), .A3(new_n582), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(KEYINPUT97), .B(G29gat), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(G36gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G43gat), .A2(G50gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(G43gat), .A2(G50gat), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT15), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n595));
  INV_X1    g394(.A(G36gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT98), .B(G50gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G43gat), .ZN(new_n603));
  AOI211_X1 g402(.A(KEYINPUT15), .B(new_n592), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n598), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT96), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n597), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n595), .A2(KEYINPUT96), .A3(new_n596), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n608), .B1(G36gat), .B2(new_n589), .ZN(new_n609));
  OAI22_X1  g408(.A1(new_n600), .A2(new_n604), .B1(new_n609), .B2(new_n594), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT17), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n614));
  INV_X1    g413(.A(G85gat), .ZN(new_n615));
  INV_X1    g414(.A(G92gat), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G99gat), .B(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n612), .A2(new_n613), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n621), .B(new_n622), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n626), .A2(new_n610), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G190gat), .B(G218gat), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G134gat), .B(G162gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n588), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n560), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n624), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(G230gat), .A3(G233gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(KEYINPUT10), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n560), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT105), .Z(new_n651));
  OAI21_X1  g450(.A(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(G120gat), .B(G148gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT104), .ZN(new_n654));
  XNOR2_X1  g453(.A(G176gat), .B(G204gat), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n654), .B(new_n655), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n658));
  INV_X1    g457(.A(new_n656), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n645), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n576), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n612), .A2(new_n663), .A3(new_n613), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n576), .A2(new_n610), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G229gat), .A2(G233gat), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT18), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n576), .B(new_n610), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n667), .B(KEYINPUT13), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G113gat), .B(G141gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G169gat), .B(G197gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT95), .B(KEYINPUT11), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT12), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n669), .A2(new_n670), .A3(new_n673), .A4(new_n680), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n640), .A2(new_n662), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n545), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n462), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n566), .ZN(G1324gat));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n457), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT106), .Z(new_n694));
  INV_X1    g493(.A(G8gat), .ZN(new_n695));
  OAI221_X1 g494(.A(new_n694), .B1(new_n692), .B2(new_n691), .C1(new_n695), .C2(new_n689), .ZN(G1325gat));
  INV_X1    g495(.A(new_n686), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT94), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n317), .B2(new_n318), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n323), .A2(KEYINPUT94), .A3(new_n316), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(G15gat), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT107), .ZN(new_n703));
  INV_X1    g502(.A(new_n325), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n704), .A2(G15gat), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n697), .B2(new_n705), .ZN(G1326gat));
  NOR2_X1   g505(.A1(new_n686), .A2(new_n495), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT108), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NOR2_X1   g509(.A1(new_n544), .A2(new_n638), .ZN(new_n711));
  INV_X1    g510(.A(new_n684), .ZN(new_n712));
  INV_X1    g511(.A(new_n588), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n713), .A3(new_n661), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n462), .A3(new_n589), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT45), .Z(new_n717));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n711), .A2(new_n718), .A3(KEYINPUT44), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n536), .A2(new_n543), .ZN(new_n720));
  INV_X1    g519(.A(new_n464), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n463), .B1(new_n457), .B2(new_n462), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n496), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n515), .A2(new_n533), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n325), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n718), .B(new_n639), .C1(new_n720), .C2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n714), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n589), .B1(new_n730), .B2(new_n462), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n717), .A2(new_n731), .ZN(G1328gat));
  OAI21_X1  g531(.A(G36gat), .B1(new_n730), .B2(new_n457), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n715), .A2(G36gat), .A3(new_n457), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n701), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n603), .B1(new_n715), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n704), .A2(G43gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n730), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g540(.A(new_n601), .B1(new_n730), .B2(new_n495), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n495), .A2(new_n601), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT110), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n715), .B2(new_n744), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT48), .Z(G1331gat));
  AND3_X1   g545(.A1(new_n712), .A2(new_n640), .A3(new_n661), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n545), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n462), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(new_n552), .ZN(G1332gat));
  NOR2_X1   g549(.A1(new_n748), .A2(new_n457), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  NOR3_X1   g554(.A1(new_n748), .A2(G71gat), .A3(new_n737), .ZN(new_n756));
  INV_X1    g555(.A(new_n748), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n704), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(G71gat), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n496), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g561(.A1(new_n713), .A2(new_n684), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n662), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n729), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766), .B2(new_n462), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n544), .B2(new_n638), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT111), .B(new_n639), .C1(new_n720), .C2(new_n725), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT112), .A4(new_n772), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n769), .A2(new_n770), .A3(new_n763), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n775), .A2(new_n776), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n661), .A2(new_n403), .A3(new_n615), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n767), .B1(new_n778), .B2(new_n779), .ZN(G1336gat));
  NAND3_X1  g579(.A1(new_n729), .A2(new_n449), .A3(new_n765), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n661), .A2(new_n616), .A3(new_n449), .ZN(new_n784));
  XOR2_X1   g583(.A(new_n784), .B(KEYINPUT113), .Z(new_n785));
  OAI211_X1 g584(.A(new_n782), .B(new_n783), .C1(new_n778), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n777), .A2(new_n771), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n787), .A2(new_n773), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n782), .B1(new_n788), .B2(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n790), .A3(KEYINPUT52), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n789), .B2(KEYINPUT52), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n786), .B1(new_n792), .B2(new_n793), .ZN(G1337gat));
  XOR2_X1   g593(.A(KEYINPUT115), .B(G99gat), .Z(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n766), .B2(new_n325), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n737), .A2(new_n662), .A3(new_n795), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n778), .B2(new_n797), .ZN(G1338gat));
  NAND4_X1  g597(.A1(new_n719), .A2(new_n728), .A3(new_n496), .A4(new_n765), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(G106gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n662), .A2(G106gat), .A3(new_n495), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT116), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n802), .B1(new_n787), .B2(new_n773), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n799), .B2(G106gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n775), .A2(new_n776), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n802), .B1(new_n806), .B2(new_n787), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n778), .A2(KEYINPUT117), .A3(new_n802), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT118), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n804), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1339gat));
  INV_X1    g614(.A(new_n651), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT54), .B(new_n658), .C1(new_n648), .C2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n648), .A2(new_n818), .A3(new_n816), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n817), .A2(KEYINPUT55), .A3(new_n656), .A4(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(new_n660), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n656), .A3(new_n819), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n684), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n666), .A2(new_n667), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n671), .A2(new_n672), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n679), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n683), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n661), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n639), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n638), .B1(new_n822), .B2(new_n823), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n821), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n588), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n712), .A2(new_n640), .A3(new_n662), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT119), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n712), .A2(new_n640), .A3(new_n662), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n841), .A2(new_n737), .A3(new_n496), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n449), .A2(new_n462), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n275), .A3(new_n712), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n841), .A2(new_n462), .A3(new_n449), .A4(new_n535), .ZN(new_n846));
  AOI21_X1  g645(.A(G113gat), .B1(new_n846), .B2(new_n684), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n845), .A2(new_n847), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n844), .B2(new_n662), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n846), .A2(new_n288), .A3(new_n661), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1341gat));
  OAI21_X1  g650(.A(G127gat), .B1(new_n844), .B2(new_n588), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n846), .A2(new_n281), .A3(new_n713), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1342gat));
  OAI21_X1  g653(.A(G134gat), .B1(new_n844), .B2(new_n638), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT120), .Z(new_n856));
  NAND3_X1  g655(.A1(new_n846), .A2(new_n279), .A3(new_n639), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT56), .Z(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1343gat));
  NAND2_X1  g658(.A1(new_n325), .A2(new_n843), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n840), .B2(new_n496), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n863), .B(new_n495), .C1(new_n834), .C2(new_n839), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(new_n712), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G141gat), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n841), .A2(new_n495), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n861), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(G141gat), .A3(new_n712), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n865), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT121), .B(new_n861), .C1(new_n862), .C2(new_n864), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n684), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n871), .B1(new_n879), .B2(G141gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n873), .B1(new_n880), .B2(new_n868), .ZN(G1344gat));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n875), .A2(new_n661), .A3(new_n876), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n354), .A2(KEYINPUT59), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n840), .A2(KEYINPUT57), .A3(new_n496), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n821), .A2(KEYINPUT123), .A3(new_n832), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n829), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT123), .B1(new_n821), .B2(new_n832), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n588), .B1(new_n890), .B2(new_n831), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n495), .B1(new_n891), .B2(new_n835), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n886), .B1(new_n892), .B2(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n861), .A2(KEYINPUT122), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n861), .A2(KEYINPUT122), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n893), .A2(new_n661), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G148gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT59), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(KEYINPUT124), .A3(KEYINPUT59), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n885), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n870), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n354), .A3(new_n661), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n882), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT124), .B1(new_n897), .B2(KEYINPUT59), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n899), .B(new_n908), .C1(new_n896), .C2(G148gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT125), .B(new_n904), .C1(new_n910), .C2(new_n885), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n906), .A2(new_n911), .ZN(G1345gat));
  OAI21_X1  g711(.A(G155gat), .B1(new_n877), .B2(new_n588), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n903), .A2(new_n339), .A3(new_n713), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  AOI21_X1  g714(.A(G162gat), .B1(new_n903), .B2(new_n639), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n638), .A2(new_n340), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n878), .B2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n403), .A2(new_n457), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT126), .Z(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n842), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n218), .A3(new_n712), .ZN(new_n923));
  NOR4_X1   g722(.A1(new_n841), .A2(new_n403), .A3(new_n457), .A4(new_n535), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n684), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n923), .A2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(G176gat), .B1(new_n922), .B2(new_n662), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n924), .A2(new_n219), .A3(new_n661), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(G1349gat));
  OAI21_X1  g728(.A(G183gat), .B1(new_n922), .B2(new_n588), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n924), .A2(new_n215), .A3(new_n713), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g732(.A(new_n211), .B1(KEYINPUT127), .B2(KEYINPUT61), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n934), .B1(new_n922), .B2(new_n638), .ZN(new_n935));
  NOR2_X1   g734(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n935), .B(new_n936), .Z(new_n937));
  NAND3_X1  g736(.A1(new_n924), .A2(new_n211), .A3(new_n639), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1351gat));
  NAND3_X1  g738(.A1(new_n869), .A2(new_n325), .A3(new_n919), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n684), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n893), .A2(new_n325), .A3(new_n921), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n684), .A2(G197gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(G1352gat));
  NOR3_X1   g744(.A1(new_n940), .A2(G204gat), .A3(new_n662), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT62), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n893), .A2(new_n661), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n921), .A2(new_n325), .ZN(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n941), .A2(new_n406), .A3(new_n713), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n943), .A2(new_n713), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n407), .A3(new_n639), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n943), .A2(new_n639), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n407), .ZN(G1355gat));
endmodule


