//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1219, new_n1220, new_n1221;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n460), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n468), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  NAND2_X1  g048(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n475), .B1(new_n464), .B2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n464), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n480), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n481), .A2(G124), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  XNOR2_X1  g062(.A(KEYINPUT3), .B(G2104), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .A3(G138), .A4(new_n480), .ZN(new_n489));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT69), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AND4_X1   g066(.A1(KEYINPUT69), .A2(new_n461), .A3(new_n463), .A4(new_n490), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n480), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AND4_X1   g072(.A1(G138), .A2(new_n461), .A3(new_n463), .A4(new_n480), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT70), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n461), .A2(new_n463), .A3(new_n490), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n461), .A2(new_n463), .A3(new_n490), .A4(KEYINPUT69), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n480), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n506), .A2(new_n507), .B1(new_n494), .B2(new_n496), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n505), .A2(new_n508), .A3(new_n509), .A4(new_n489), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n500), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT72), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT5), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n513), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(KEYINPUT71), .B1(new_n524), .B2(KEYINPUT6), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n526), .A2(new_n527), .A3(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n524), .A2(KEYINPUT6), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(new_n519), .ZN(new_n532));
  INV_X1    g107(.A(G88), .ZN(new_n533));
  INV_X1    g108(.A(G50), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(G543), .ZN(new_n535));
  OAI221_X1 g110(.A(new_n523), .B1(new_n532), .B2(new_n533), .C1(new_n534), .C2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT73), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n529), .A2(new_n530), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n514), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G51), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n520), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G89), .ZN(new_n545));
  AND2_X1   g120(.A1(G63), .A2(G651), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n519), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n540), .A2(new_n543), .A3(new_n545), .A4(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n524), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n542), .A2(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n544), .A2(G90), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(G301));
  INV_X1    g129(.A(G301), .ZN(G171));
  AOI22_X1  g130(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n524), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n542), .A2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n544), .A2(G81), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  XOR2_X1   g139(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n565));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G188));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n535), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n542), .A2(new_n571), .A3(G53), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n520), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(G91), .A2(new_n544), .B1(new_n576), .B2(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n544), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n542), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  AND2_X1   g157(.A1(new_n519), .A2(G61), .ZN(new_n583));
  AND2_X1   g158(.A1(G73), .A2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n529), .A2(new_n519), .A3(G86), .A4(new_n530), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n529), .A2(G48), .A3(G543), .A4(new_n530), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n542), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT75), .B(G85), .Z(new_n591));
  OAI221_X1 g166(.A(new_n589), .B1(new_n524), .B2(new_n590), .C1(new_n532), .C2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NOR2_X1   g172(.A1(G301), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n532), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT77), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n520), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(G54), .A2(new_n542), .B1(new_n607), .B2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n598), .B1(new_n611), .B2(new_n597), .ZN(G284));
  XOR2_X1   g187(.A(G284), .B(KEYINPUT79), .Z(G321));
  NAND2_X1  g188(.A1(G299), .A2(new_n597), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(new_n597), .B2(G168), .ZN(G297));
  OAI21_X1  g190(.A(new_n614), .B1(new_n597), .B2(G168), .ZN(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n560), .A2(new_n597), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n609), .B(KEYINPUT78), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n620), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n621), .B2(new_n597), .ZN(G323));
  XOR2_X1   g197(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n623));
  XNOR2_X1  g198(.A(G323), .B(new_n623), .ZN(G282));
  NAND2_X1  g199(.A1(new_n478), .A2(G135), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n480), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n481), .A2(G123), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT82), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND2_X1  g207(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n465), .A2(G2104), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT12), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  NOR2_X1   g211(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n632), .B(new_n638), .C1(new_n636), .C2(new_n633), .ZN(G156));
  INV_X1    g214(.A(G14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n640), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n652), .A2(KEYINPUT83), .A3(new_n654), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT83), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n651), .B2(new_n653), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n664), .B(KEYINPUT17), .Z(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n661), .B2(new_n662), .ZN(new_n669));
  INV_X1    g244(.A(new_n661), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(new_n664), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n663), .B1(new_n671), .B2(new_n662), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n667), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n683), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n679), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(KEYINPUT86), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT86), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n679), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n687), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n703), .A3(new_n701), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  NAND2_X1  g283(.A1(new_n481), .A2(G119), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n480), .A2(G107), .ZN(new_n710));
  OAI21_X1  g285(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n711));
  INV_X1    g286(.A(G131), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n709), .B1(new_n710), .B2(new_n711), .C1(new_n477), .C2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G25), .B(new_n713), .S(G29), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(G16), .A2(G24), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(G290), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT89), .B(G1986), .Z(new_n720));
  OAI21_X1  g295(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(G22), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G166), .B2(new_n718), .ZN(new_n724));
  INV_X1    g299(.A(G1971), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G23), .B(G288), .S(G16), .Z(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT33), .B(G1976), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G6), .A2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G305), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G16), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT32), .B(G1981), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n726), .A2(new_n729), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT34), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT34), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n726), .A2(new_n737), .A3(new_n729), .A4(new_n734), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n722), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT36), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(G115), .A2(G2104), .ZN(new_n742));
  INV_X1    g317(.A(G127), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n464), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT25), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n744), .A2(G2105), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G139), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n477), .B2(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G33), .B(new_n751), .S(G29), .Z(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2072), .Z(new_n753));
  AND3_X1   g328(.A1(new_n474), .A2(G141), .A3(new_n476), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT26), .Z(new_n756));
  NAND3_X1  g331(.A1(new_n480), .A2(G105), .A3(G2104), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT93), .ZN(new_n758));
  INV_X1    g333(.A(G129), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n488), .A2(G2105), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n756), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n763), .B2(G32), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT27), .B(G1996), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT94), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(G34), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n768), .B2(G34), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G160), .B2(G29), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n765), .A2(new_n767), .B1(G2084), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n753), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT95), .ZN(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  AOI211_X1 g352(.A(G29), .B(new_n777), .C1(KEYINPUT30), .C2(new_n775), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT31), .B(G11), .Z(new_n779));
  AOI211_X1 g354(.A(new_n778), .B(new_n779), .C1(new_n630), .C2(G29), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n780), .B1(G2084), .B2(new_n771), .C1(new_n767), .C2(new_n765), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n718), .A2(G21), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G168), .B2(new_n718), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n783), .A2(G1966), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(G1966), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n781), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n763), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n763), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(G2078), .Z(new_n789));
  NAND2_X1  g364(.A1(new_n718), .A2(G5), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G171), .B2(new_n718), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT97), .B(G1961), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n774), .A2(new_n786), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(KEYINPUT98), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT98), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n774), .A2(new_n797), .A3(new_n786), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n763), .A2(G26), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT28), .Z(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n801));
  INV_X1    g376(.A(G116), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G2105), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n481), .A2(new_n804), .A3(G128), .ZN(new_n805));
  INV_X1    g380(.A(G128), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT91), .B1(new_n760), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n803), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n474), .A2(G140), .A3(new_n476), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n800), .B1(new_n810), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT92), .ZN(new_n812));
  INV_X1    g387(.A(G2067), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n718), .A2(G20), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT23), .Z(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G299), .B2(G16), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1956), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n763), .A2(G35), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G162), .B2(new_n763), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT29), .B(G2090), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n718), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n561), .B2(new_n718), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1341), .Z(new_n825));
  NAND4_X1  g400(.A1(new_n814), .A2(new_n818), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G4), .A2(G16), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT90), .Z(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n620), .B2(new_n718), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n796), .A2(new_n798), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n741), .A2(new_n833), .ZN(G311));
  OAI21_X1  g409(.A(KEYINPUT99), .B1(new_n741), .B2(new_n833), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n739), .B(KEYINPUT36), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT99), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n798), .A2(new_n832), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n796), .A4(new_n838), .ZN(new_n839));
  AND2_X1   g414(.A1(new_n835), .A2(new_n839), .ZN(G150));
  NAND2_X1  g415(.A1(new_n611), .A2(G559), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(new_n524), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n531), .A2(G93), .A3(new_n519), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n529), .A2(G55), .A3(G543), .A4(new_n530), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(KEYINPUT100), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(KEYINPUT100), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n560), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n846), .A2(new_n847), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(new_n848), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n561), .A3(new_n845), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n843), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n843), .A2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n851), .A2(G860), .ZN(new_n868));
  XOR2_X1   g443(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT102), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(G145));
  NAND3_X1  g450(.A1(new_n488), .A2(G130), .A3(G2105), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(G106), .A2(G2105), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n879), .B(G2104), .C1(G118), .C2(new_n480), .ZN(new_n880));
  INV_X1    g455(.A(G142), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n878), .B(new_n880), .C1(new_n881), .C2(new_n477), .ZN(new_n882));
  OAI211_X1 g457(.A(KEYINPUT103), .B(new_n749), .C1(new_n477), .C2(new_n750), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n882), .B(new_n883), .Z(new_n884));
  NOR2_X1   g459(.A1(new_n493), .A2(new_n499), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n810), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n808), .A3(new_n809), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n762), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n751), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n762), .B1(new_n887), .B2(new_n888), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n884), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n713), .B(new_n635), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n888), .ZN(new_n896));
  INV_X1    g471(.A(new_n762), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n882), .B(new_n883), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n889), .A4(new_n891), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n894), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n895), .B1(new_n894), .B2(new_n900), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n630), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n894), .A2(new_n900), .ZN(new_n906));
  INV_X1    g481(.A(new_n895), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n630), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n908), .A2(new_n902), .A3(new_n909), .A4(new_n901), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n486), .B(G160), .ZN(new_n912));
  AOI21_X1  g487(.A(G37), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n905), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g492(.A(G303), .B(G288), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n594), .A2(G305), .A3(new_n595), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G305), .B1(new_n594), .B2(new_n595), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(G290), .A2(new_n731), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n918), .A3(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT41), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n609), .A2(G299), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n609), .A2(G299), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n609), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n573), .A3(new_n577), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(KEYINPUT41), .A3(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n621), .A2(new_n858), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n611), .A2(new_n617), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(new_n859), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n935), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n621), .A2(new_n858), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n937), .A2(new_n859), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n933), .A2(new_n928), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n940), .A3(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n939), .B2(new_n944), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n926), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n939), .A2(new_n944), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  INV_X1    g525(.A(new_n926), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n945), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n597), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n851), .A2(new_n597), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT106), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n946), .A2(new_n926), .A3(new_n947), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n951), .B1(new_n950), .B2(new_n945), .ZN(new_n958));
  OAI21_X1  g533(.A(G868), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n954), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n961), .ZN(G295));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n954), .ZN(G331));
  NAND2_X1  g538(.A1(G168), .A2(G171), .ZN(new_n964));
  NAND2_X1  g539(.A1(G286), .A2(G301), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n851), .A2(new_n560), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n561), .B1(new_n856), .B2(new_n845), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n852), .A2(new_n857), .A3(new_n965), .A4(new_n964), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n928), .A4(new_n933), .ZN(new_n971));
  INV_X1    g546(.A(new_n970), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n858), .A2(KEYINPUT107), .A3(new_n966), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n926), .B(new_n971), .C1(new_n976), .C2(new_n935), .ZN(new_n977));
  INV_X1    g552(.A(G37), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n943), .B(new_n972), .C1(new_n974), .C2(new_n975), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n935), .B1(new_n970), .B2(new_n969), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n951), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n980), .A2(KEYINPUT43), .A3(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n858), .A2(KEYINPUT107), .A3(new_n966), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT107), .B1(new_n858), .B2(new_n966), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n970), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n935), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n926), .B1(new_n989), .B2(new_n971), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT43), .B1(new_n980), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT44), .B1(new_n984), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT43), .B1(new_n979), .B2(new_n990), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n983), .A2(new_n977), .A3(new_n995), .A4(new_n978), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n993), .B1(KEYINPUT44), .B2(new_n997), .ZN(G397));
  AOI22_X1  g573(.A1(new_n503), .A2(new_n504), .B1(new_n498), .B2(KEYINPUT4), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n999), .B2(new_n508), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1000), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n762), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n810), .B(new_n813), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n1003), .B2(new_n762), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n1006), .B(new_n1007), .C1(new_n1002), .C2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1002), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n713), .B(new_n715), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1013), .B1(new_n1002), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n467), .A2(G40), .A3(new_n471), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1000), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1017), .B(G8), .C1(new_n1018), .C2(G288), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT52), .ZN(new_n1020));
  INV_X1    g595(.A(G1384), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(new_n493), .B2(new_n499), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(new_n1001), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1025), .B(new_n1026), .C1(new_n1018), .C2(G288), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n584), .B1(new_n519), .B2(G61), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n524), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n586), .A2(new_n587), .ZN(new_n1030));
  OAI21_X1  g605(.A(G1981), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(KEYINPUT111), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT110), .B(G1981), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n1031), .A3(KEYINPUT111), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1025), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1033), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1020), .B(new_n1027), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G303), .A2(G8), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT55), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT45), .B(new_n1021), .C1(new_n493), .C2(new_n499), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1384), .B1(new_n500), .B2(new_n510), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1016), .B(new_n1044), .C1(new_n1045), .C2(KEYINPUT45), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n725), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1001), .B1(new_n1000), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT109), .B(G2090), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1049), .B(new_n1050), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1024), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1040), .B1(new_n1043), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n509), .B1(new_n999), .B2(new_n508), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n509), .A2(new_n505), .A3(new_n508), .A4(new_n489), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1048), .B(new_n1021), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1001), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n1050), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1044), .A2(new_n1016), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1021), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1058), .B1(new_n1062), .B2(G1971), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1024), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1047), .A2(KEYINPUT114), .A3(new_n1058), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1043), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1053), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT115), .B(new_n1043), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1048), .B1(new_n511), .B2(new_n1021), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1016), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT116), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1961), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1049), .B(new_n1076), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT122), .B(KEYINPUT53), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1079), .B1(new_n1046), .B2(G2078), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1016), .B1(new_n1000), .B2(KEYINPUT45), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1081), .A2(new_n1082), .A3(G2078), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n1061), .B2(new_n1060), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1078), .A2(new_n1080), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1044), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1078), .A2(new_n1080), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(G171), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n1090));
  INV_X1    g665(.A(G1966), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1061), .B(G1384), .C1(new_n500), .C2(new_n510), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n1081), .ZN(new_n1093));
  INV_X1    g668(.A(G2084), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1049), .B(new_n1094), .C1(new_n1045), .C2(new_n1048), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(G168), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G8), .ZN(new_n1097));
  AOI21_X1  g672(.A(G168), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT51), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1100), .A3(G8), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1089), .A2(new_n1090), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1090), .B1(new_n1088), .B2(G171), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(G171), .B2(new_n1085), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1071), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1074), .A2(new_n830), .A3(new_n1077), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1023), .A2(new_n813), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT60), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1106), .A2(KEYINPUT120), .A3(KEYINPUT60), .A4(new_n1107), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1110), .A2(new_n932), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n609), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT121), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1110), .A2(new_n932), .A3(new_n1111), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1113), .A4(new_n1116), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT58), .B(G1341), .Z(new_n1122));
  AOI22_X1  g697(.A1(new_n1062), .A2(new_n1003), .B1(new_n1017), .B2(new_n1122), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1123), .A2(new_n560), .B1(KEYINPUT118), .B2(KEYINPUT59), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1017), .A2(new_n1122), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n1046), .B2(G1996), .ZN(new_n1126));
  NOR2_X1   g701(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n561), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1124), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g705(.A(KEYINPUT56), .B(G2072), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1046), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1956), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT57), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n573), .B2(new_n577), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1133), .A2(new_n1134), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1137), .A2(new_n1136), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1134), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1062), .A2(new_n1131), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1140), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1138), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1139), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1130), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g723(.A(KEYINPUT119), .B(new_n1130), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1118), .A2(new_n1121), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n609), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1138), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1143), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1105), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1052), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n1042), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT112), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1040), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1040), .A2(new_n1159), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1035), .ZN(new_n1163));
  OR2_X1    g738(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1164));
  NOR2_X1   g739(.A1(G288), .A2(G1976), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT113), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1025), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1162), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1099), .A2(new_n1171), .A3(new_n1101), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1086), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1170), .B1(new_n1176), .B2(new_n1071), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1179), .A2(G8), .A3(G168), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1158), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1157), .A2(new_n1042), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1181), .B(new_n1182), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1183));
  NOR3_X1   g758(.A1(new_n1069), .A2(new_n1070), .A3(new_n1180), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1183), .B1(new_n1184), .B2(KEYINPUT63), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1177), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1015), .B1(new_n1156), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1188));
  NAND2_X1  g763(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1188), .B(new_n1189), .Z(new_n1190));
  AND2_X1   g765(.A1(new_n1008), .A2(new_n762), .ZN(new_n1191));
  OAI221_X1 g766(.A(new_n1190), .B1(KEYINPUT124), .B2(KEYINPUT46), .C1(new_n1011), .C2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g767(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  NOR3_X1   g769(.A1(G290), .A2(G1986), .A3(new_n1011), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1195), .B(KEYINPUT48), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1194), .B1(new_n1013), .B2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n810), .A2(G2067), .ZN(new_n1198));
  INV_X1    g773(.A(new_n715), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n713), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1198), .B1(new_n1010), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT123), .ZN(new_n1202));
  OR2_X1    g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1011), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1197), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1187), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n994), .A2(new_n996), .ZN(new_n1209));
  INV_X1    g783(.A(G319), .ZN(new_n1210));
  NOR2_X1   g784(.A1(G227), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g785(.A(new_n1211), .B(KEYINPUT126), .ZN(new_n1212));
  NAND3_X1  g786(.A1(new_n707), .A2(new_n659), .A3(new_n1212), .ZN(new_n1213));
  INV_X1    g787(.A(new_n1213), .ZN(new_n1214));
  AND4_X1   g788(.A1(new_n1208), .A2(new_n1209), .A3(new_n916), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1213), .B1(new_n913), .B2(new_n915), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1208), .B1(new_n1216), .B2(new_n1209), .ZN(new_n1217));
  NOR2_X1   g791(.A1(new_n1215), .A2(new_n1217), .ZN(G308));
  NAND2_X1  g792(.A1(new_n916), .A2(new_n1214), .ZN(new_n1219));
  OAI21_X1  g793(.A(KEYINPUT127), .B1(new_n1219), .B2(new_n997), .ZN(new_n1220));
  NAND3_X1  g794(.A1(new_n1216), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1220), .A2(new_n1221), .ZN(G225));
endmodule


