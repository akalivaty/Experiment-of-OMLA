//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G87), .B(G97), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT65), .ZN(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  XNOR2_X1  g0046(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n247));
  INV_X1    g0047(.A(G232), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n253), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  AOI21_X1  g0055(.A(G1698), .B1(new_n251), .B2(new_n252), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(G226), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  OAI211_X1 g0060(.A(G226), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n254), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(KEYINPUT68), .A3(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n265), .A2(KEYINPUT66), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G33), .A3(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(new_n264), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G41), .A2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n276), .A2(G1), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n278), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n281), .A2(new_n282), .B1(new_n284), .B2(G238), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n247), .B1(new_n271), .B2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n268), .A2(new_n269), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n251), .A2(new_n252), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n289), .A2(new_n255), .A3(G226), .A4(new_n258), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n287), .B1(new_n291), .B2(new_n254), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n275), .A2(G238), .A3(new_n283), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n278), .ZN(new_n294));
  AOI21_X1  g0094(.A(KEYINPUT67), .B1(new_n275), .B2(new_n278), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n247), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n292), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(G169), .B1(new_n286), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT14), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT14), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(G169), .C1(new_n286), .C2(new_n298), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n271), .A2(new_n247), .A3(new_n285), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT13), .B1(new_n292), .B2(new_n296), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(new_n304), .A3(G179), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n305), .A2(KEYINPUT74), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(KEYINPUT74), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n300), .B(new_n302), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n214), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n206), .A2(G33), .ZN(new_n311));
  INV_X1    g0111(.A(G77), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n311), .A2(new_n312), .B1(new_n206), .B2(G68), .ZN(new_n313));
  INV_X1    g0113(.A(G50), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G20), .A2(G33), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n313), .A2(KEYINPUT73), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n313), .A2(KEYINPUT73), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT11), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT12), .B1(new_n322), .B2(G68), .ZN(new_n323));
  OR3_X1    g0123(.A1(new_n322), .A2(KEYINPUT12), .A3(G68), .ZN(new_n324));
  INV_X1    g0124(.A(new_n322), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n310), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n218), .B1(new_n205), .B2(G20), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n323), .A2(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n319), .B2(new_n320), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n308), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n303), .A2(new_n304), .A3(G190), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n330), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n297), .B1(new_n292), .B2(new_n296), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n303), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n325), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT69), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n326), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n205), .A2(G20), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT69), .B1(new_n325), .B2(new_n310), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n343), .B1(new_n348), .B2(new_n342), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G58), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n218), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n201), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n315), .A2(G159), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n251), .A2(new_n206), .A3(new_n252), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n251), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n252), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n355), .B1(new_n360), .B2(G68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n310), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(KEYINPUT75), .A3(new_n359), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT75), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n356), .A2(new_n365), .A3(new_n357), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(G68), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n355), .ZN(new_n368));
  AOI21_X1  g0168(.A(KEYINPUT16), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n350), .B1(new_n363), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n275), .A2(G232), .A3(new_n283), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n294), .B2(new_n295), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT77), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n374), .B(new_n371), .C1(new_n294), .C2(new_n295), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n250), .A2(new_n220), .ZN(new_n376));
  NOR2_X1   g0176(.A1(G223), .A2(G1698), .ZN(new_n377));
  INV_X1    g0177(.A(G226), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(G1698), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n376), .B1(new_n379), .B2(new_n289), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n380), .A2(KEYINPUT76), .B1(new_n268), .B2(new_n269), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(G1698), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G223), .B2(G1698), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n259), .A2(new_n260), .ZN(new_n384));
  OAI22_X1  g0184(.A1(new_n383), .A2(new_n384), .B1(new_n250), .B2(new_n220), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT76), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  AND4_X1   g0188(.A1(G179), .A2(new_n373), .A3(new_n375), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G169), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n372), .A2(KEYINPUT77), .B1(new_n381), .B2(new_n387), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n375), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n370), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT18), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n367), .A2(new_n368), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n310), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n361), .B2(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n349), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n373), .A2(new_n375), .A3(new_n388), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G200), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n391), .A2(G190), .A3(new_n375), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n407), .B(new_n370), .C1(new_n389), .C2(new_n392), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT17), .A4(new_n403), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n394), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  XOR2_X1   g0211(.A(new_n341), .B(KEYINPUT70), .Z(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n315), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT15), .B(G87), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n413), .B1(new_n206), .B2(new_n312), .C1(new_n311), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n310), .ZN(new_n416));
  INV_X1    g0216(.A(new_n326), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n346), .A2(G77), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(G77), .B2(new_n322), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n281), .A2(new_n282), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n284), .A2(G244), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n253), .A2(new_n258), .ZN(new_n425));
  INV_X1    g0225(.A(G107), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n289), .A2(G1698), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n425), .B1(new_n426), .B2(new_n289), .C1(new_n427), .C2(new_n219), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(new_n270), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G179), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n429), .A2(G169), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n421), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n419), .B1(new_n415), .B2(new_n310), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(G190), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n434), .B(new_n435), .C1(new_n336), .C2(new_n429), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n256), .A2(G222), .ZN(new_n438));
  INV_X1    g0238(.A(G223), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n438), .B1(new_n312), .B2(new_n289), .C1(new_n439), .C2(new_n427), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n270), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n284), .A2(G226), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n441), .A2(new_n422), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n345), .A2(G50), .A3(new_n346), .A4(new_n347), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n325), .A2(new_n314), .ZN(new_n445));
  INV_X1    g0245(.A(G150), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n341), .A2(new_n311), .B1(new_n446), .B2(new_n316), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n206), .B1(new_n201), .B2(new_n314), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n310), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n445), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n443), .A2(new_n336), .B1(KEYINPUT9), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n441), .A2(new_n422), .A3(new_n442), .ZN(new_n453));
  INV_X1    g0253(.A(G190), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT9), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n453), .A2(new_n454), .B1(new_n455), .B2(new_n450), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT10), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n456), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n453), .A2(G200), .B1(new_n455), .B2(new_n450), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT10), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n443), .A2(new_n430), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n453), .A2(new_n390), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n450), .A3(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n437), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n340), .A2(new_n411), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n322), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n205), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n322), .A2(new_n470), .A3(new_n214), .A4(new_n309), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n469), .B1(new_n472), .B2(new_n468), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(KEYINPUT78), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n364), .A2(G107), .A3(new_n366), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n426), .A2(KEYINPUT6), .A3(G97), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n468), .A2(new_n426), .ZN(new_n477));
  NOR2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(KEYINPUT6), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(G20), .B1(G77), .B2(new_n315), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n398), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g0283(.A(KEYINPUT5), .B(G41), .Z(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n275), .B(G257), .C1(new_n484), .C2(new_n487), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n275), .A2(G274), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(G244), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n491), .B1(new_n270), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT79), .B1(new_n499), .B2(new_n336), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n270), .ZN(new_n501));
  INV_X1    g0301(.A(new_n491), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT79), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n504), .A3(G200), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n499), .A2(G190), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n483), .A2(new_n500), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT78), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n473), .B(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n475), .A2(new_n481), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n398), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(new_n390), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n499), .A2(new_n430), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n206), .B(G87), .C1(new_n259), .C2(new_n260), .ZN(new_n515));
  XOR2_X1   g0315(.A(KEYINPUT82), .B(KEYINPUT22), .Z(new_n516));
  XNOR2_X1  g0316(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT24), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT23), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(new_n426), .A3(G20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G116), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  OAI221_X1 g0323(.A(new_n520), .B1(G20), .B2(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n517), .A2(new_n518), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n518), .B1(new_n517), .B2(new_n526), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n310), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT25), .B1(new_n325), .B2(new_n426), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n325), .A2(KEYINPUT25), .A3(new_n426), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n531), .A2(new_n532), .B1(G107), .B2(new_n472), .ZN(new_n533));
  OAI211_X1 g0333(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n535));
  INV_X1    g0335(.A(G294), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n535), .C1(new_n250), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n214), .B1(KEYINPUT66), .B2(new_n265), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n274), .A2(new_n538), .B1(new_n489), .B2(new_n486), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n537), .A2(new_n270), .B1(new_n539), .B2(G264), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(G190), .A3(new_n490), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n490), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n529), .A2(new_n533), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n507), .A2(new_n514), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n275), .B(G270), .C1(new_n484), .C2(new_n487), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n546), .A2(new_n490), .ZN(new_n547));
  OAI211_X1 g0347(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n548));
  OAI211_X1 g0348(.A(G257), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n251), .A2(G303), .A3(new_n252), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n270), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(G116), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n325), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n309), .A2(new_n214), .B1(G20), .B2(new_n554), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n496), .B(new_n206), .C1(G33), .C2(new_n468), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n556), .A2(KEYINPUT20), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT20), .B1(new_n556), .B2(new_n557), .ZN(new_n559));
  OAI221_X1 g0359(.A(new_n555), .B1(new_n554), .B2(new_n471), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n553), .A2(G169), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n560), .A2(G179), .A3(new_n552), .A4(new_n547), .ZN(new_n564));
  INV_X1    g0364(.A(new_n560), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n551), .A2(new_n270), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n546), .A2(new_n490), .ZN(new_n567));
  OAI21_X1  g0367(.A(G200), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n565), .B(new_n568), .C1(new_n553), .C2(new_n454), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n553), .A2(KEYINPUT21), .A3(new_n560), .A4(G169), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n563), .A2(new_n564), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n529), .A2(new_n533), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n390), .B1(new_n540), .B2(new_n490), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n540), .A2(G179), .A3(new_n490), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n311), .B2(new_n468), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n289), .A2(new_n206), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n218), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT81), .B(G87), .ZN(new_n583));
  NAND3_X1  g0383(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n583), .A2(new_n478), .B1(new_n206), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n310), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n414), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(new_n322), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n472), .A2(G87), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n486), .B2(new_n221), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n275), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n260), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT80), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n289), .A2(KEYINPUT80), .A3(G244), .A4(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n289), .A2(G238), .A3(new_n258), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n521), .A4(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n595), .B1(new_n601), .B2(new_n270), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n591), .B1(G190), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n336), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(new_n270), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G179), .A3(new_n594), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n390), .B2(new_n602), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n586), .A2(new_n589), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n472), .A2(new_n587), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n603), .A2(new_n605), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n571), .A2(new_n578), .A3(new_n612), .ZN(new_n613));
  NOR3_X1   g0413(.A1(new_n467), .A2(new_n545), .A3(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n465), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n332), .B1(new_n339), .B2(new_n433), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n406), .A3(new_n409), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n394), .A2(new_n408), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n615), .B1(new_n619), .B2(new_n462), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n507), .A2(new_n514), .A3(new_n544), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n570), .A2(new_n564), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n390), .B1(new_n547), .B2(new_n552), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT21), .B1(new_n623), .B2(new_n560), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n578), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n602), .A2(G190), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n627), .A2(new_n604), .A3(new_n591), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n602), .A2(new_n390), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n430), .B(new_n595), .C1(new_n601), .C2(new_n270), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT85), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT85), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n607), .B(new_n632), .C1(new_n390), .C2(new_n602), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n628), .B1(new_n634), .B2(new_n611), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n621), .A2(new_n626), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n611), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n514), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n603), .A2(new_n605), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n608), .A2(new_n611), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n514), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n643), .A2(KEYINPUT86), .B1(KEYINPUT26), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT86), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n641), .A2(new_n648), .A3(new_n642), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n638), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n620), .B1(new_n467), .B2(new_n650), .ZN(G369));
  NAND3_X1  g0451(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n565), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n622), .B2(new_n624), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n563), .A2(new_n569), .A3(new_n564), .A4(new_n570), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(G330), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n578), .A2(new_n657), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n572), .A2(new_n657), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n544), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n666), .B1(new_n578), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n658), .B1(new_n622), .B2(new_n624), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n578), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(G399));
  INV_X1    g0475(.A(new_n209), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G1), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n583), .A2(new_n554), .A3(new_n478), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n679), .A2(new_n680), .B1(new_n212), .B2(new_n678), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT28), .Z(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT26), .B1(new_n639), .B2(new_n612), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n609), .A2(new_n610), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n631), .B2(new_n633), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n685), .A2(new_n514), .A3(new_n628), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n687));
  OAI211_X1 g0487(.A(KEYINPUT29), .B(new_n658), .C1(new_n638), .C2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n641), .A2(new_n642), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n637), .B(new_n636), .C1(new_n691), .C2(new_n683), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(KEYINPUT91), .A3(KEYINPUT29), .A4(new_n658), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT86), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n646), .A2(KEYINPUT26), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n649), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n638), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n657), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n690), .B(new_n693), .C1(KEYINPUT29), .C2(new_n698), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n613), .A2(new_n545), .A3(new_n657), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT90), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n503), .A2(new_n430), .A3(new_n553), .ZN(new_n702));
  INV_X1    g0502(.A(new_n542), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n702), .A2(new_n703), .A3(new_n602), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n552), .A2(G179), .A3(new_n490), .A4(new_n546), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT89), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT89), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n547), .A2(new_n707), .A3(G179), .A4(new_n552), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n503), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT88), .B1(new_n602), .B2(new_n540), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n602), .A2(KEYINPUT88), .A3(new_n540), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n704), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n709), .B(KEYINPUT30), .C1(new_n710), .C2(new_n711), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n658), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n700), .A2(new_n701), .B1(KEYINPUT31), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(KEYINPUT31), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n703), .A2(G179), .B1(new_n573), .B2(KEYINPUT84), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n573), .A2(KEYINPUT84), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n720), .A2(new_n721), .B1(new_n529), .B2(new_n533), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n645), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n621), .A3(new_n571), .A4(new_n658), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT90), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n717), .A2(new_n719), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n699), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n682), .B1(new_n728), .B2(new_n205), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT92), .ZN(G364));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n205), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n677), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n676), .A2(new_n384), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G355), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G116), .B2(new_n209), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n245), .A2(G45), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT93), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n676), .A2(new_n289), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n742), .B1(new_n485), .B2(new_n213), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n738), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n214), .B1(G20), .B2(new_n390), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT94), .Z(new_n750));
  OAI21_X1  g0550(.A(new_n735), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G179), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n468), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n206), .A2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n430), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n206), .A2(new_n454), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n758), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n289), .B1(new_n759), .B2(new_n312), .C1(new_n351), .C2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G190), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n756), .B(new_n762), .C1(G68), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n757), .A2(new_n752), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT32), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n763), .A2(new_n454), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n768), .A2(KEYINPUT32), .B1(new_n770), .B2(G50), .ZN(new_n771));
  INV_X1    g0571(.A(new_n583), .ZN(new_n772));
  OR3_X1    g0572(.A1(new_n336), .A2(KEYINPUT95), .A3(G179), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT95), .B1(new_n336), .B2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n773), .A2(new_n774), .A3(new_n760), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n773), .A2(new_n774), .A3(new_n757), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n772), .A2(new_n776), .B1(new_n778), .B2(G107), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n765), .A2(new_n769), .A3(new_n771), .A4(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n776), .A2(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(KEYINPUT96), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n384), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT97), .Z(new_n786));
  INV_X1    g0586(.A(new_n761), .ZN(new_n787));
  INV_X1    g0587(.A(new_n759), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G322), .A2(new_n787), .B1(new_n788), .B2(G311), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n767), .A2(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n777), .ZN(new_n792));
  INV_X1    g0592(.A(G317), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT33), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT33), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n764), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n770), .ZN(new_n797));
  INV_X1    g0597(.A(G326), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n797), .B2(new_n798), .C1(new_n755), .C2(new_n536), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n792), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n780), .B1(new_n786), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n751), .B1(new_n801), .B2(new_n748), .ZN(new_n802));
  INV_X1    g0602(.A(new_n747), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n662), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT98), .Z(new_n805));
  INV_X1    g0605(.A(new_n735), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n663), .B2(new_n664), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n664), .B2(new_n663), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n421), .A2(new_n657), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n436), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n433), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n433), .A2(new_n657), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n437), .A2(new_n658), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n698), .A2(new_n815), .B1(new_n650), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n735), .B1(new_n817), .B2(new_n727), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n727), .B2(new_n817), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n748), .A2(new_n745), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n806), .B1(new_n312), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n748), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G143), .A2(new_n787), .B1(new_n788), .B2(G159), .ZN(new_n823));
  INV_X1    g0623(.A(new_n764), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n446), .C1(new_n825), .C2(new_n797), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT34), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n783), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(G50), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n777), .A2(new_n218), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n289), .B1(new_n766), .B2(new_n832), .C1(new_n755), .C2(new_n351), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(new_n826), .C2(new_n827), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT99), .B(G283), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n756), .B1(new_n764), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n784), .B2(new_n797), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n777), .A2(new_n220), .ZN(new_n839));
  INV_X1    g0639(.A(G311), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n384), .B1(new_n766), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n761), .A2(new_n536), .B1(new_n759), .B2(new_n554), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n829), .A2(G107), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n830), .A2(new_n834), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n821), .B1(new_n822), .B2(new_n845), .C1(new_n815), .C2(new_n746), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n819), .A2(new_n846), .ZN(G384));
  OAI21_X1  g0647(.A(new_n620), .B1(new_n699), .B2(new_n467), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT102), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n332), .A2(new_n657), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n350), .B1(new_n363), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n655), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n410), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n852), .B1(new_n389), .B2(new_n392), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(new_n404), .A3(new_n854), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n370), .A2(new_n853), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n393), .A2(new_n404), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n856), .A2(new_n863), .A3(KEYINPUT38), .ZN(new_n864));
  XNOR2_X1  g0664(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n865));
  INV_X1    g0665(.A(new_n861), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n393), .A2(new_n404), .A3(new_n861), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n410), .A2(new_n866), .B1(new_n868), .B2(new_n862), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n864), .B(new_n865), .C1(KEYINPUT38), .C2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT39), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n856), .A2(new_n863), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT38), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n872), .B1(new_n875), .B2(new_n864), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n850), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n864), .ZN(new_n878));
  INV_X1    g0678(.A(new_n339), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n330), .A2(new_n658), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n332), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n331), .B(new_n657), .C1(new_n308), .C2(new_n339), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n816), .B1(new_n696), .B2(new_n697), .ZN(new_n885));
  INV_X1    g0685(.A(new_n814), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n878), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n618), .A2(new_n853), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  AND4_X1   g0689(.A1(KEYINPUT101), .A2(new_n877), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n856), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT38), .B1(new_n856), .B2(new_n863), .ZN(new_n892));
  OAI21_X1  g0692(.A(KEYINPUT39), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n870), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n888), .B1(new_n894), .B2(new_n850), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT101), .B1(new_n895), .B2(new_n887), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n849), .B(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n813), .A2(new_n814), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n882), .B2(new_n883), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n712), .A2(new_n713), .ZN(new_n902));
  INV_X1    g0702(.A(new_n704), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n715), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n905));
  INV_X1    g0705(.A(new_n613), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n906), .A2(new_n701), .A3(new_n621), .A4(new_n658), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n725), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT103), .B1(new_n716), .B2(KEYINPUT31), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n904), .A2(new_n657), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT103), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT31), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n901), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n891), .A2(new_n892), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n899), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n410), .A2(new_n866), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n868), .A2(new_n862), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n874), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n899), .B1(new_n921), .B2(new_n864), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n717), .A2(new_n725), .A3(new_n909), .A4(new_n913), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n901), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n467), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n923), .ZN(new_n927));
  OAI21_X1  g0727(.A(G330), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n928), .B1(new_n925), .B2(new_n927), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n898), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n898), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n205), .B2(new_n732), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n930), .B1(new_n932), .B2(KEYINPUT104), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(KEYINPUT104), .B2(new_n932), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(G116), .A3(new_n215), .A4(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n212), .A2(new_n312), .A3(new_n352), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n218), .A2(G50), .ZN(new_n940));
  OAI211_X1 g0740(.A(G1), .B(new_n731), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(G367));
  OAI221_X1 g0742(.A(new_n749), .B1(new_n209), .B2(new_n414), .C1(new_n742), .C2(new_n237), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n759), .A2(new_n314), .B1(new_n766), .B2(new_n825), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n384), .B(new_n944), .C1(G150), .C2(new_n787), .ZN(new_n945));
  INV_X1    g0745(.A(G159), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n755), .A2(new_n218), .B1(new_n946), .B2(new_n824), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G143), .B2(new_n770), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n776), .A2(G58), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n778), .A2(G77), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n945), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n829), .A2(KEYINPUT46), .A3(G116), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT110), .Z(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT46), .B1(new_n776), .B2(G116), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n754), .A2(G107), .B1(G294), .B2(new_n764), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n840), .B2(new_n797), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n777), .A2(new_n468), .ZN(new_n957));
  AOI22_X1  g0757(.A1(G303), .A2(new_n787), .B1(new_n767), .B2(G317), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n289), .B1(new_n788), .B2(new_n836), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR4_X1    g0760(.A1(new_n954), .A2(new_n956), .A3(new_n957), .A4(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n951), .B1(new_n953), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  OAI211_X1 g0763(.A(new_n735), .B(new_n943), .C1(new_n963), .C2(new_n822), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n591), .A2(new_n657), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n637), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n635), .B2(new_n965), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(new_n747), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT109), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n507), .B(new_n514), .C1(new_n483), .C2(new_n658), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n639), .A2(new_n657), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OR3_X1    g0775(.A1(new_n674), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n972), .B1(new_n674), .B2(new_n975), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n674), .A2(new_n975), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n674), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AND3_X1   g0783(.A1(new_n978), .A2(new_n983), .A3(new_n670), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n670), .B1(new_n978), .B2(new_n983), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n669), .B(new_n672), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT107), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n665), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n987), .B(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n728), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n677), .B(new_n993), .Z(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT108), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n977), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n674), .A2(new_n972), .A3(new_n975), .ZN(new_n998));
  INV_X1    g0798(.A(new_n982), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT45), .B1(new_n674), .B2(new_n975), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n997), .A2(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n670), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n978), .A2(new_n983), .A3(new_n670), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n727), .B(new_n699), .C1(new_n1005), .C2(new_n990), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT108), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n1007), .A3(new_n994), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n996), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n733), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n669), .A2(new_n672), .A3(new_n975), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT42), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n514), .B1(new_n973), .B2(new_n578), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1012), .B1(new_n658), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n1015));
  AND2_X1   g0815(.A1(new_n967), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  MUX2_X1   g0817(.A(KEYINPUT43), .B(new_n1015), .S(new_n967), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n975), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n670), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n670), .A2(new_n1020), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1017), .B(new_n1022), .C1(new_n1014), .C2(new_n1018), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n971), .B1(new_n1010), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n734), .B1(new_n996), .B2(new_n1008), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1027), .A2(KEYINPUT109), .A3(new_n1024), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n970), .B1(new_n1026), .B2(new_n1028), .ZN(G387));
  AOI22_X1  g0829(.A1(new_n736), .A2(new_n680), .B1(new_n426), .B2(new_n676), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n412), .A2(new_n314), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n485), .B1(new_n218), .B2(new_n312), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n1032), .A2(new_n680), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n741), .B1(new_n233), .B2(new_n485), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1030), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n750), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n806), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G50), .A2(new_n787), .B1(new_n767), .B2(G150), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n1039), .B(new_n289), .C1(new_n218), .C2(new_n759), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n587), .A2(new_n754), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n824), .B2(new_n341), .C1(new_n946), .C2(new_n797), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n775), .A2(new_n312), .ZN(new_n1043));
  NOR4_X1   g0843(.A1(new_n1040), .A2(new_n1042), .A3(new_n957), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G317), .A2(new_n787), .B1(new_n788), .B2(G303), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n770), .A2(G322), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n840), .C2(new_n824), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT48), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n776), .A2(G294), .B1(new_n754), .B2(new_n836), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n384), .B1(new_n766), .B2(new_n798), .C1(new_n777), .C2(new_n554), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT111), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1044), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1038), .B1(new_n822), .B2(new_n1058), .C1(new_n669), .C2(new_n803), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT112), .Z(new_n1060));
  AND2_X1   g0860(.A1(new_n728), .A2(new_n990), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n677), .B(KEYINPUT113), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n728), .B2(new_n990), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1060), .B1(new_n733), .B2(new_n990), .C1(new_n1061), .C2(new_n1063), .ZN(G393));
  INV_X1    g0864(.A(new_n1062), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n728), .A2(new_n990), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n986), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n984), .A2(KEYINPUT114), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1005), .B2(KEYINPUT114), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1020), .A2(new_n747), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n242), .A2(new_n742), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n749), .B1(new_n468), .B2(new_n209), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n735), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n384), .B1(new_n759), .B2(new_n536), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n755), .A2(new_n554), .B1(new_n784), .B2(new_n824), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1075), .B(new_n1076), .C1(G322), .C2(new_n767), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n426), .B2(new_n777), .C1(new_n775), .C2(new_n835), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n787), .A2(G311), .B1(G317), .B2(new_n770), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n839), .B1(new_n412), .B2(new_n788), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n218), .B2(new_n775), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n824), .A2(new_n314), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n384), .B(new_n1083), .C1(G143), .C2(new_n767), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n787), .A2(G159), .B1(G150), .B2(new_n770), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT51), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(KEYINPUT51), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n754), .A2(G77), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1078), .A2(new_n1080), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1074), .B1(new_n1090), .B2(new_n748), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1069), .A2(new_n734), .B1(new_n1071), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT115), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1070), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1093), .B1(new_n1070), .B2(new_n1092), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(G390));
  OAI211_X1 g0897(.A(new_n658), .B(new_n813), .C1(new_n638), .C2(new_n687), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n1098), .A2(new_n814), .B1(new_n882), .B2(new_n883), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n850), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT38), .B1(new_n918), .B2(new_n919), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n891), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n726), .A2(G330), .A3(new_n815), .A4(new_n884), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n814), .B1(new_n650), .B2(new_n816), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n850), .B1(new_n1106), .B2(new_n884), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1105), .C1(new_n1107), .C2(new_n894), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1100), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n871), .A2(new_n876), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1103), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n923), .A2(G330), .A3(new_n901), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1108), .B(new_n734), .C1(new_n1112), .C2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n820), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n735), .B1(new_n342), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1088), .B1(new_n554), .B2(new_n761), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT116), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n384), .B1(new_n766), .B2(new_n536), .C1(new_n468), .C2(new_n759), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n824), .A2(new_n426), .B1(new_n797), .B2(new_n791), .ZN(new_n1120));
  OR4_X1    g0920(.A1(new_n831), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n783), .A2(new_n220), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n776), .A2(G150), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT53), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n755), .A2(new_n946), .B1(new_n825), .B2(new_n824), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(G128), .B2(new_n770), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n778), .A2(G50), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  AOI21_X1  g0928(.A(new_n384), .B1(new_n788), .B2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(G132), .A2(new_n787), .B1(new_n767), .B2(G125), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1121), .A2(new_n1122), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1116), .B1(new_n1132), .B2(new_n748), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n894), .B2(new_n746), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1114), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1108), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n905), .B1(new_n724), .B2(KEYINPUT90), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n613), .A2(new_n545), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n701), .B1(new_n1138), .B2(new_n658), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n909), .A2(new_n913), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n664), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(G330), .B(new_n815), .C1(new_n908), .C2(new_n718), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n884), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n901), .A2(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1106), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n884), .B1(new_n1142), .B2(new_n815), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n1098), .A2(new_n814), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1105), .A2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1145), .A2(new_n1146), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1142), .A2(new_n926), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n620), .C1(new_n699), .C2(new_n467), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1062), .B1(new_n1136), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1113), .B1(new_n1156), .B2(new_n1104), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1158), .A2(new_n1108), .B1(new_n1153), .B2(new_n1150), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1135), .B1(new_n1155), .B2(new_n1159), .ZN(G378));
  XNOR2_X1  g0960(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT119), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n462), .A2(new_n1163), .A3(new_n465), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n450), .A2(new_n853), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT55), .Z(new_n1167));
  AOI21_X1  g0967(.A(new_n1163), .B1(new_n462), .B2(new_n465), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1167), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n462), .A2(new_n465), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT119), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1170), .B1(new_n1172), .B2(new_n1164), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1162), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1167), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1172), .A2(new_n1170), .A3(new_n1164), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n1161), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  AND4_X1   g0978(.A1(G330), .A2(new_n917), .A3(new_n1178), .A4(new_n924), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n883), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n339), .B(new_n880), .C1(new_n308), .C2(new_n331), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n815), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n664), .B1(new_n1183), .B2(new_n922), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1178), .B1(new_n1184), .B2(new_n917), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n890), .A2(new_n896), .B1(new_n1179), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n877), .A2(new_n887), .A3(new_n889), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT101), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n895), .A2(KEYINPUT101), .A3(new_n887), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(new_n917), .A3(new_n1178), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1178), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT40), .B1(new_n1183), .B2(new_n878), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT40), .B1(new_n891), .B2(new_n1101), .ZN(new_n1194));
  OAI21_X1  g0994(.A(G330), .B1(new_n915), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1192), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1186), .A2(new_n1197), .A3(new_n734), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n735), .B1(G50), .B2(new_n1115), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n289), .A2(G41), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n775), .B2(new_n312), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n1201), .A2(KEYINPUT117), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT117), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n777), .A2(new_n351), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G283), .B2(new_n767), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT118), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n761), .A2(new_n426), .B1(new_n759), .B2(new_n414), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G68), .B2(new_n754), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n764), .A2(G97), .B1(new_n770), .B2(G116), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT58), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1213), .B1(new_n946), .B2(new_n777), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n776), .A2(new_n1128), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G128), .A2(new_n787), .B1(new_n788), .B2(G137), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n764), .A2(G132), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n754), .A2(G150), .B1(G125), .B2(new_n770), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1214), .B1(new_n1219), .B2(KEYINPUT59), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(KEYINPUT59), .B2(new_n1219), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n314), .B1(G33), .B2(G41), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1212), .B(new_n1221), .C1(new_n1200), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1199), .B1(new_n1223), .B2(new_n748), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n1178), .B2(new_n746), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1198), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1186), .A2(new_n1197), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1149), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n923), .A2(G330), .A3(new_n815), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1144), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1113), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1229), .A2(new_n1231), .B1(new_n1233), .B2(new_n1106), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1153), .B1(new_n1136), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1156), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1237), .A2(new_n1157), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1152), .B1(new_n1238), .B2(new_n1150), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1186), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1062), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1227), .B1(new_n1236), .B2(new_n1241), .ZN(G375));
  NAND2_X1  g1042(.A1(new_n1144), .A2(new_n745), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n735), .B1(G68), .B2(new_n1115), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n829), .A2(G97), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1041), .B1(new_n824), .B2(new_n554), .C1(new_n536), .C2(new_n797), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n761), .A2(new_n791), .B1(new_n759), .B2(new_n426), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n289), .B(new_n1248), .C1(G303), .C2(new_n767), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1245), .A2(new_n950), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n829), .A2(G159), .B1(G128), .B2(new_n767), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT122), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1128), .A2(new_n764), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n797), .B2(new_n832), .C1(new_n755), .C2(new_n314), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n289), .B1(new_n759), .B2(new_n446), .C1(new_n825), .C2(new_n761), .ZN(new_n1255));
  OR3_X1    g1055(.A1(new_n1254), .A2(new_n1204), .A3(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1250), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1244), .B1(new_n1257), .B2(new_n748), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1150), .A2(new_n734), .B1(new_n1243), .B2(new_n1258), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n994), .B(KEYINPUT121), .Z(new_n1260));
  NAND2_X1  g1060(.A1(new_n1154), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(G381));
  OR2_X1    g1063(.A1(G393), .A2(G396), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(G390), .A2(G384), .A3(new_n1264), .A4(G381), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1010), .A2(new_n971), .A3(new_n1025), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT109), .B1(new_n1027), .B2(new_n1024), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n969), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G378), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1197), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1065), .B1(new_n1270), .B2(new_n1235), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT57), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1186), .A2(new_n1197), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1239), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1226), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1265), .A2(new_n1268), .A3(new_n1269), .A4(new_n1275), .ZN(G407));
  NAND3_X1  g1076(.A1(new_n1275), .A2(new_n656), .A3(new_n1269), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(G407), .A2(G213), .A3(new_n1277), .ZN(G409));
  INV_X1    g1078(.A(KEYINPUT126), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(G393), .B(new_n809), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT125), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n970), .B(new_n1096), .C1(new_n1026), .C2(new_n1028), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1096), .B1(new_n1288), .B2(new_n970), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1283), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1285), .B1(new_n1268), .B2(new_n1096), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G387), .A2(G390), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1282), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1233), .A2(new_n1106), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1231), .A2(new_n1148), .A3(new_n1105), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1294), .A2(new_n1152), .A3(new_n1295), .A4(KEYINPUT60), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1154), .A2(new_n1296), .A3(new_n1062), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT60), .B1(new_n1234), .B2(new_n1152), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1259), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(G384), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G384), .B(new_n1259), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n656), .A2(G213), .ZN(new_n1303));
  INV_X1    g1103(.A(G2897), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(KEYINPUT123), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1305), .B1(KEYINPUT123), .B2(new_n1304), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1301), .A2(new_n1302), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT124), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT124), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1301), .A2(new_n1309), .A3(new_n1302), .A4(new_n1306), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1308), .A2(new_n1310), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1304), .B(new_n1303), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1228), .A2(new_n1235), .A3(new_n1260), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G378), .B1(new_n1227), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1275), .B2(G378), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1303), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1311), .B(new_n1313), .C1(new_n1316), .C2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1290), .A2(new_n1293), .A3(new_n1318), .A4(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G378), .B(new_n1227), .C1(new_n1236), .C2(new_n1241), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1228), .A2(new_n1235), .A3(new_n1260), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1269), .B1(new_n1322), .B2(new_n1226), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1301), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1302), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1324), .A2(new_n1327), .A3(new_n1303), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1328), .B(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1279), .B1(new_n1320), .B2(new_n1330), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1287), .A2(new_n1289), .A3(new_n1283), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1282), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1328), .B(KEYINPUT63), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1334), .A2(new_n1335), .A3(KEYINPUT126), .A4(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT127), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1318), .A2(new_n1338), .A3(new_n1319), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1338), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1328), .A2(KEYINPUT62), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1324), .A2(new_n1342), .A3(new_n1327), .A4(new_n1303), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1339), .A2(new_n1340), .A3(new_n1344), .ZN(new_n1345));
  OAI211_X1 g1145(.A(new_n1331), .B(new_n1337), .C1(new_n1345), .C2(new_n1334), .ZN(G405));
  NAND2_X1  g1146(.A1(G375), .A2(new_n1269), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(new_n1321), .ZN(new_n1348));
  XOR2_X1   g1148(.A(new_n1348), .B(new_n1327), .Z(new_n1349));
  XNOR2_X1  g1149(.A(new_n1349), .B(new_n1334), .ZN(G402));
endmodule


