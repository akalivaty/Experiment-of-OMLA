//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  NOR3_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(KEYINPUT87), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n206), .B1(KEYINPUT87), .B2(new_n205), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n208), .B(KEYINPUT88), .ZN(new_n209));
  OAI211_X1 g008(.A(KEYINPUT15), .B(new_n203), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n211));
  AOI22_X1  g010(.A1(KEYINPUT89), .A2(new_n211), .B1(new_n209), .B2(KEYINPUT91), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT91), .B2(new_n209), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n205), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n204), .B1(new_n205), .B2(new_n215), .ZN(new_n217));
  OAI221_X1 g016(.A(new_n214), .B1(new_n211), .B2(KEYINPUT89), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n210), .B1(new_n213), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n210), .B(KEYINPUT17), .C1(new_n213), .C2(new_n218), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n221), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT93), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n231), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n219), .B(new_n231), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n236), .B(KEYINPUT13), .Z(new_n241));
  AOI22_X1  g040(.A1(new_n238), .A2(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n236), .A4(new_n237), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT94), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n249), .B1(new_n242), .B2(new_n243), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI211_X1 g052(.A(KEYINPUT94), .B(new_n249), .C1(new_n242), .C2(new_n243), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n202), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n252), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT94), .A3(new_n250), .ZN(new_n257));
  INV_X1    g056(.A(new_n254), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(KEYINPUT95), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT28), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n262));
  INV_X1    g061(.A(G183gat), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT27), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G190gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT27), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT64), .A3(G183gat), .ZN(new_n267));
  AND4_X1   g066(.A1(new_n261), .A2(new_n264), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT27), .B(G183gat), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n261), .B1(new_n269), .B2(new_n265), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT65), .B1(new_n268), .B2(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G169gat), .ZN(new_n276));
  INV_X1    g075(.A(G176gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT66), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(KEYINPUT26), .B2(new_n278), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G120gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G113gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G120gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT67), .A3(G134gat), .ZN(new_n292));
  INV_X1    g091(.A(G134gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G127gat), .ZN(new_n296));
  INV_X1    g095(.A(G127gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n297), .A3(new_n294), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n276), .A2(new_n277), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT23), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n281), .A2(KEYINPUT24), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n263), .A2(new_n265), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(KEYINPUT24), .A3(new_n281), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT25), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n284), .A2(new_n299), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n296), .A2(new_n298), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n282), .B1(new_n273), .B2(new_n274), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n306), .B(KEYINPUT25), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G15gat), .B(G43gat), .Z(new_n317));
  XNOR2_X1  g116(.A(new_n317), .B(KEYINPUT68), .ZN(new_n318));
  XNOR2_X1  g117(.A(G71gat), .B(G99gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT33), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(KEYINPUT32), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT69), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n316), .A2(new_n324), .A3(KEYINPUT32), .A4(new_n321), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT33), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n320), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n316), .B2(KEYINPUT32), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n323), .A2(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n309), .A2(new_n313), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT34), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(new_n314), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT71), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n315), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n338), .B2(KEYINPUT34), .ZN(new_n339));
  AOI211_X1 g138(.A(KEYINPUT71), .B(new_n332), .C1(new_n336), .C2(new_n337), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n330), .B(new_n333), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT70), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT70), .B1(new_n309), .B2(new_n313), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(new_n315), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT71), .B1(new_n345), .B2(new_n332), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n334), .A3(KEYINPUT34), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n330), .B1(new_n348), .B2(new_n333), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n350));
  NOR3_X1   g149(.A1(new_n342), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n333), .B1(new_n339), .B2(new_n340), .ZN(new_n352));
  INV_X1    g151(.A(new_n330), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n354), .A2(new_n341), .B1(KEYINPUT72), .B2(KEYINPUT36), .ZN(new_n355));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356));
  INV_X1    g155(.A(G155gat), .ZN(new_n357));
  INV_X1    g156(.A(G162gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n356), .B1(new_n359), .B2(KEYINPUT2), .ZN(new_n360));
  INV_X1    g159(.A(G141gat), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT76), .B1(new_n361), .B2(G148gat), .ZN(new_n362));
  INV_X1    g161(.A(G148gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(G141gat), .B2(new_n363), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n361), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n360), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G141gat), .B(G148gat), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n356), .B(new_n359), .C1(new_n367), .C2(KEYINPUT2), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n372), .A2(new_n296), .A3(new_n298), .A4(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n369), .B1(new_n296), .B2(new_n298), .ZN(new_n378));
  XOR2_X1   g177(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n375), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n310), .A2(new_n370), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n385), .B2(new_n378), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n378), .B2(new_n380), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n386), .B(KEYINPUT5), .C1(new_n388), .C2(new_n376), .ZN(new_n389));
  XOR2_X1   g188(.A(G1gat), .B(G29gat), .Z(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n383), .A2(new_n389), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n389), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n394), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT6), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n389), .A3(KEYINPUT80), .A4(new_n395), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n394), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT73), .ZN(new_n411));
  XNOR2_X1  g210(.A(G197gat), .B(G204gat), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT22), .ZN(new_n413));
  INV_X1    g212(.A(G211gat), .ZN(new_n414));
  INV_X1    g213(.A(G218gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT73), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n410), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n417), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G226gat), .ZN(new_n424));
  INV_X1    g223(.A(G233gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n284), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT74), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n429), .B1(new_n311), .B2(new_n312), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n311), .A2(new_n312), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n432), .A2(KEYINPUT29), .A3(new_n426), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n423), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT75), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT29), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n428), .A2(new_n430), .A3(new_n436), .A4(new_n427), .ZN(new_n437));
  INV_X1    g236(.A(new_n423), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n426), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n434), .A2(new_n435), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n435), .B1(new_n434), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n409), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n434), .A2(new_n440), .A3(new_n408), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n434), .A2(new_n440), .A3(KEYINPUT30), .A4(new_n408), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n405), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G228gat), .A2(G233gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT3), .B1(new_n423), .B2(new_n436), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n453), .B1(new_n454), .B2(new_n370), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n423), .B1(new_n372), .B2(new_n436), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(KEYINPUT83), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT81), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n418), .A2(new_n422), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n436), .B1(new_n422), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n371), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n457), .B1(new_n466), .B2(new_n369), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT82), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n467), .A2(new_n468), .A3(new_n453), .ZN(new_n469));
  INV_X1    g268(.A(new_n371), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n411), .A2(new_n417), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT29), .B1(new_n471), .B2(KEYINPUT81), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n472), .B2(new_n463), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n458), .B1(new_n473), .B2(new_n370), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT82), .B1(new_n474), .B2(new_n452), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n461), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT84), .B1(new_n476), .B2(G22gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT31), .B(G50gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n476), .A2(G22gat), .ZN(new_n482));
  INV_X1    g281(.A(G22gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n468), .B1(new_n467), .B2(new_n453), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n474), .A2(KEYINPUT82), .A3(new_n452), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n483), .B1(new_n486), .B2(new_n461), .ZN(new_n487));
  OAI22_X1  g286(.A1(new_n477), .A2(new_n481), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n476), .A2(G22gat), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n483), .A3(new_n461), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n489), .A2(KEYINPUT84), .A3(new_n490), .A4(new_n480), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n351), .A2(new_n355), .B1(new_n451), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT36), .ZN(new_n497));
  OAI22_X1  g296(.A1(new_n342), .A2(new_n349), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n350), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n354), .A2(new_n341), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n491), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n484), .A2(new_n485), .B1(new_n460), .B2(new_n459), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n504), .B2(new_n483), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n505), .A2(new_n480), .B1(new_n489), .B2(new_n490), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n443), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n408), .B1(new_n508), .B2(new_n441), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(new_n449), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n405), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n501), .A2(KEYINPUT85), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT40), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n382), .A2(new_n374), .A3(new_n381), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT39), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n384), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n395), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n299), .A2(new_n369), .ZN(new_n519));
  INV_X1    g318(.A(new_n378), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n375), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT39), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n522), .B1(new_n515), .B2(new_n384), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n514), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n524), .A2(new_n400), .ZN(new_n525));
  OR3_X1    g324(.A1(new_n518), .A2(new_n523), .A3(new_n514), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n525), .B(new_n526), .C1(new_n509), .C2(new_n449), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT37), .B1(new_n442), .B2(new_n443), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT37), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n434), .A2(new_n529), .A3(new_n440), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n530), .A2(KEYINPUT38), .A3(new_n409), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n438), .B1(new_n431), .B2(new_n433), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n437), .A2(new_n423), .A3(new_n439), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT37), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n534), .A3(new_n409), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT38), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n528), .A2(new_n531), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n403), .A2(new_n404), .A3(new_n445), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n492), .B(new_n527), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n495), .A2(new_n513), .A3(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n341), .B(new_n354), .C1(new_n502), .C2(new_n506), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT35), .B1(new_n541), .B2(new_n511), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n342), .A2(new_n349), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT35), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n451), .A2(new_n543), .A3(new_n544), .A4(new_n492), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n260), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G57gat), .B(G64gat), .Z(new_n548));
  OR2_X1    g347(.A1(G71gat), .A2(G78gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n548), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n550), .B(new_n549), .C1(new_n555), .C2(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(G127gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n232), .B1(new_n558), .B2(new_n557), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n357), .ZN(new_n566));
  XOR2_X1   g365(.A(G183gat), .B(G211gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n564), .B(new_n568), .Z(new_n569));
  AND2_X1   g368(.A1(G232gat), .A2(G233gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT41), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT96), .ZN(new_n572));
  XOR2_X1   g371(.A(G134gat), .B(G162gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT98), .Z(new_n575));
  NAND2_X1  g374(.A1(G85gat), .A2(G92gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(KEYINPUT97), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n579), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT8), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n578), .A2(new_n580), .A3(new_n582), .A4(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n581), .ZN(new_n587));
  NOR2_X1   g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n586), .B(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n221), .A2(new_n233), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n219), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n570), .ZN(new_n593));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n591), .B2(new_n593), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n575), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n574), .A2(KEYINPUT98), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(new_n601), .A3(new_n596), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n569), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT99), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT100), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n586), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n608), .B2(new_n557), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n587), .A2(new_n588), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n586), .B1(new_n611), .B2(KEYINPUT100), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n607), .A2(new_n613), .A3(new_n578), .A4(new_n580), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n554), .A2(new_n556), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT101), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n590), .A2(new_n557), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n609), .A2(new_n610), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n592), .A2(KEYINPUT10), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT103), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n617), .A3(new_n618), .ZN(new_n625));
  INV_X1    g424(.A(new_n622), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n621), .A2(new_n628), .A3(new_n622), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n626), .B1(new_n621), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(new_n636), .B2(new_n621), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n627), .A3(new_n633), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n605), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n547), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n405), .B(KEYINPUT104), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  INV_X1    g447(.A(new_n510), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT105), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n222), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n644), .A2(new_n649), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n653), .B2(new_n222), .ZN(new_n654));
  MUX2_X1   g453(.A(new_n652), .B(new_n654), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g454(.A(G15gat), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n644), .A2(new_n656), .A3(new_n543), .ZN(new_n657));
  INV_X1    g456(.A(new_n501), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n644), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n657), .B1(new_n659), .B2(new_n656), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT106), .ZN(G1326gat));
  NAND2_X1  g460(.A1(new_n644), .A2(new_n507), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  OR2_X1    g463(.A1(new_n603), .A2(KEYINPUT109), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n603), .A2(KEYINPUT109), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n501), .A2(new_n539), .A3(new_n668), .A4(new_n512), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n546), .A2(new_n669), .ZN(new_n670));
  AOI22_X1  g469(.A1(new_n498), .A2(new_n500), .B1(new_n507), .B2(new_n511), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n671), .B2(new_n539), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n667), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n539), .B1(new_n671), .B2(KEYINPUT85), .ZN(new_n675));
  INV_X1    g474(.A(new_n513), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n546), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n603), .A2(new_n674), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n673), .A2(new_n674), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n569), .A2(new_n640), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n253), .A2(new_n254), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT110), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n492), .A2(new_n527), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n537), .A2(new_n538), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT108), .B1(new_n493), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n546), .A3(new_n669), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n690), .B2(new_n667), .ZN(new_n691));
  INV_X1    g490(.A(new_n678), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n692), .B1(new_n540), .B2(new_n546), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n694));
  INV_X1    g493(.A(new_n684), .ZN(new_n695));
  NOR4_X1   g494(.A1(new_n691), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n685), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n645), .ZN(new_n699));
  INV_X1    g498(.A(new_n603), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n680), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT107), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n547), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(G29gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n646), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(new_n706), .ZN(G1328gat));
  OAI21_X1  g506(.A(G36gat), .B1(new_n698), .B2(new_n510), .ZN(new_n708));
  INV_X1    g507(.A(G36gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n703), .A2(new_n709), .A3(new_n649), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT46), .Z(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n673), .A2(new_n674), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n677), .A2(new_n678), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n684), .ZN(new_n716));
  OAI21_X1  g515(.A(G43gat), .B1(new_n716), .B2(new_n501), .ZN(new_n717));
  INV_X1    g516(.A(G43gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n718), .A3(new_n543), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT47), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n718), .B1(new_n697), .B2(new_n658), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n713), .B(new_n721), .C1(new_n722), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n716), .A2(new_n694), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n679), .A2(KEYINPUT110), .A3(new_n684), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n726), .A2(new_n658), .A3(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n728), .B2(G43gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n723), .B1(new_n717), .B2(new_n719), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT111), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n725), .A2(new_n731), .ZN(G1330gat));
  OAI21_X1  g531(.A(G50gat), .B1(new_n716), .B2(new_n492), .ZN(new_n733));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n703), .A2(new_n734), .A3(new_n507), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(KEYINPUT48), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n735), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n697), .A2(new_n507), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(G50gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n739), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n682), .A2(new_n641), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n690), .A2(new_n605), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n646), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n649), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT49), .B(G64gat), .Z(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n745), .B2(new_n747), .ZN(G1333gat));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n658), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n342), .A2(new_n349), .A3(G71gat), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n749), .A2(G71gat), .B1(new_n742), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n742), .A2(new_n507), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  INV_X1    g553(.A(new_n679), .ZN(new_n755));
  INV_X1    g554(.A(new_n569), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT112), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n755), .A2(new_n645), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n690), .A2(new_n683), .A3(new_n756), .A4(new_n700), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT51), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n646), .A2(new_n583), .A3(new_n640), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n759), .A2(new_n583), .B1(new_n761), .B2(new_n762), .ZN(G1336gat));
  INV_X1    g562(.A(new_n761), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n510), .A2(G92gat), .A3(new_n641), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT52), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n755), .A2(new_n758), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n649), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G92gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n760), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT51), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n768), .A2(G92gat), .B1(new_n773), .B2(new_n765), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(G1337gat));
  NOR3_X1   g575(.A1(new_n755), .A2(new_n501), .A3(new_n758), .ZN(new_n777));
  INV_X1    g576(.A(G99gat), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n543), .A2(new_n778), .A3(new_n640), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n777), .A2(new_n778), .B1(new_n761), .B2(new_n779), .ZN(G1338gat));
  NOR3_X1   g579(.A1(new_n492), .A2(G106gat), .A3(new_n641), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n764), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n507), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n783), .A2(G106gat), .B1(new_n773), .B2(new_n781), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(G1339gat));
  NAND3_X1  g587(.A1(new_n619), .A2(new_n626), .A3(new_n620), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n638), .A2(KEYINPUT54), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT54), .B1(new_n624), .B2(new_n629), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n633), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n628), .B1(new_n621), .B2(new_n622), .ZN(new_n795));
  AOI211_X1 g594(.A(KEYINPUT103), .B(new_n626), .C1(new_n619), .C2(new_n620), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(KEYINPUT114), .A3(new_n634), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n790), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n639), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n801), .B(new_n790), .C1(new_n793), .C2(new_n798), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT115), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n790), .ZN(new_n804));
  INV_X1    g603(.A(new_n798), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT114), .B1(new_n797), .B2(new_n634), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n801), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n804), .B(KEYINPUT55), .C1(new_n805), .C2(new_n806), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n808), .A2(new_n809), .A3(new_n639), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n803), .A2(new_n682), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n240), .A2(new_n241), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT116), .Z(new_n814));
  AOI21_X1  g613(.A(new_n236), .B1(new_n234), .B2(new_n237), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n248), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n250), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n641), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n667), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n667), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n821), .A2(new_n817), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n803), .A3(new_n811), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n756), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n643), .A2(new_n683), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(KEYINPUT117), .A3(new_n826), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n541), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n646), .A2(new_n510), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n835), .A2(new_n287), .A3(new_n260), .ZN(new_n836));
  INV_X1    g635(.A(new_n835), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n682), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n836), .B1(new_n838), .B2(new_n287), .ZN(G1340gat));
  NOR2_X1   g638(.A1(new_n835), .A2(new_n641), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(new_n285), .ZN(G1341gat));
  NAND3_X1  g640(.A1(new_n837), .A2(KEYINPUT118), .A3(new_n569), .ZN(new_n842));
  XOR2_X1   g641(.A(KEYINPUT67), .B(G127gat), .Z(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n845), .B1(new_n835), .B2(new_n756), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n842), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n837), .A2(KEYINPUT118), .A3(new_n569), .A4(new_n843), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1342gat));
  XOR2_X1   g648(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n831), .A2(new_n832), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n833), .A2(new_n603), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n851), .B1(new_n854), .B2(G134gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(G134gat), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n852), .A2(new_n293), .A3(new_n853), .A4(new_n850), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G1343gat));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n829), .A2(new_n859), .A3(new_n507), .A4(new_n830), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n833), .A2(new_n658), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n260), .A2(new_n802), .A3(new_n800), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n603), .B1(new_n863), .B2(new_n818), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n569), .B1(new_n864), .B2(new_n823), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n642), .A2(new_n682), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n507), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n867), .B2(KEYINPUT57), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT122), .B1(new_n869), .B2(new_n260), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871));
  INV_X1    g670(.A(new_n260), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n860), .A2(new_n871), .A3(new_n868), .A4(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n870), .A2(G141gat), .A3(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n829), .A2(new_n507), .A3(new_n830), .A4(new_n861), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n260), .A2(G141gat), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT121), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n875), .A2(KEYINPUT121), .A3(new_n877), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n860), .A2(new_n682), .A3(new_n868), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n884), .A2(new_n885), .A3(G141gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n884), .B2(G141gat), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n875), .A2(new_n877), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n883), .B1(new_n889), .B2(new_n879), .ZN(G1344gat));
  INV_X1    g689(.A(new_n875), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n363), .A3(new_n640), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n507), .A2(new_n859), .ZN(new_n894));
  INV_X1    g693(.A(new_n864), .ZN(new_n895));
  NOR4_X1   g694(.A1(new_n800), .A2(new_n802), .A3(new_n817), .A4(new_n603), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n756), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n643), .A2(new_n260), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n829), .A2(new_n507), .A3(new_n830), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n640), .A3(new_n861), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n893), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n869), .A2(new_n641), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(KEYINPUT59), .A3(new_n363), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n892), .B1(new_n903), .B2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n869), .B2(new_n756), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n357), .A3(new_n569), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n869), .B2(new_n821), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n891), .A2(new_n358), .A3(new_n700), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n646), .A2(new_n510), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n829), .A2(new_n832), .A3(new_n830), .A4(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n276), .A3(new_n682), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n872), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT123), .B1(new_n917), .B2(G169gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n914), .A2(new_n641), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(new_n277), .ZN(G1349gat));
  OAI21_X1  g722(.A(new_n263), .B1(new_n914), .B2(new_n756), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n915), .A2(new_n569), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n269), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n926), .B(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n915), .A2(new_n265), .A3(new_n667), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n914), .B2(new_n603), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT124), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n933), .B(G190gat), .C1(new_n914), .C2(new_n603), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n931), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(G1351gat));
  INV_X1    g736(.A(new_n913), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n492), .A3(new_n658), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n831), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n682), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT125), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n901), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI211_X1 g743(.A(KEYINPUT125), .B(new_n899), .C1(new_n900), .C2(KEYINPUT57), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n938), .A2(new_n658), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(G197gat), .A3(new_n872), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n941), .B1(new_n947), .B2(new_n949), .ZN(G1352gat));
  OAI211_X1 g749(.A(new_n640), .B(new_n948), .C1(new_n943), .C2(new_n945), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G204gat), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n641), .A2(G204gat), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n831), .A2(new_n939), .A3(new_n953), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  NAND2_X1  g754(.A1(new_n952), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n414), .A3(new_n569), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n948), .A2(new_n569), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n414), .B1(new_n901), .B2(new_n959), .ZN(new_n960));
  OR2_X1    g759(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n960), .B2(new_n961), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n957), .B1(new_n962), .B2(new_n964), .ZN(G1354gat));
  AOI21_X1  g764(.A(G218gat), .B1(new_n940), .B2(new_n667), .ZN(new_n966));
  INV_X1    g765(.A(new_n948), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n967), .B1(new_n944), .B2(new_n946), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n603), .A2(new_n415), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT127), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(G1355gat));
endmodule


