//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n456), .A2(G2106), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT69), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n464), .B1(new_n463), .B2(new_n462), .ZN(G319));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n466), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT70), .B(G2105), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT70), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT70), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n471), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n470), .A2(G2104), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n469), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n474), .A2(new_n475), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n468), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n468), .C2(G112), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n482), .B2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n466), .A2(KEYINPUT71), .A3(new_n470), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n486), .B1(G136), .B2(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g070(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n476), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n496), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  MUX2_X1   g076(.A(G102), .B(G114), .S(G2105), .Z(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2104), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n466), .A2(G126), .A3(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n501), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G50), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n515), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT5), .B(G543), .Z(new_n524));
  NAND2_X1  g099(.A1(new_n510), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n517), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n508), .A2(new_n509), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(G90), .B1(new_n534), .B2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  AOI22_X1  g112(.A1(new_n532), .A2(G81), .B1(new_n534), .B2(G43), .ZN(new_n538));
  XOR2_X1   g113(.A(new_n538), .B(KEYINPUT73), .Z(new_n539));
  AOI22_X1  g114(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n517), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G65), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n524), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n555), .B2(new_n513), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n511), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n534), .A2(new_n559), .A3(G53), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n556), .B1(KEYINPUT75), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n558), .A2(new_n563), .A3(new_n560), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND2_X1  g142(.A1(new_n532), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n534), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  INV_X1    g146(.A(G48), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n511), .B1(new_n513), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n517), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(KEYINPUT76), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n574), .A2(new_n576), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n578), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n532), .A2(G85), .B1(new_n534), .B2(G47), .ZN(new_n583));
  XOR2_X1   g158(.A(new_n583), .B(KEYINPUT77), .Z(new_n584));
  AOI22_X1  g159(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n585), .A2(new_n517), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n532), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n524), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n534), .B2(G54), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(new_n588), .ZN(G284));
  AOI21_X1  g172(.A(new_n589), .B1(new_n596), .B2(new_n588), .ZN(G321));
  MUX2_X1   g173(.A(G286), .B(G299), .S(new_n588), .Z(G297));
  MUX2_X1   g174(.A(G286), .B(G299), .S(new_n588), .Z(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n596), .B1(new_n601), .B2(G860), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT78), .ZN(G148));
  NAND3_X1  g178(.A1(new_n596), .A2(KEYINPUT79), .A3(new_n601), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n591), .A2(new_n595), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G559), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g186(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT12), .Z(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT13), .Z(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(G2100), .ZN(new_n617));
  OAI221_X1 g192(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n468), .C2(G111), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n483), .A2(G123), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n618), .B(new_n619), .C1(new_n490), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n616), .A2(new_n617), .A3(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT15), .B(G2435), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2427), .ZN(new_n627));
  INV_X1    g202(.A(G2430), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n624), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(new_n628), .B2(new_n627), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G1341), .B(G1348), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n630), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT17), .Z(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT80), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n645), .ZN(new_n648));
  INV_X1    g223(.A(new_n641), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n648), .B(new_n644), .C1(new_n649), .C2(new_n645), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(new_n643), .A3(new_n645), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT81), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  OR3_X1    g240(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G229));
  MUX2_X1   g248(.A(G6), .B(G305), .S(G16), .Z(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT32), .B(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(G16), .A2(G23), .ZN(new_n677));
  AND3_X1   g252(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT84), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(G288), .A2(KEYINPUT84), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n677), .B1(new_n682), .B2(G16), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT33), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(G16), .A2(G22), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G166), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1971), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n676), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT34), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT82), .B(G29), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G25), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n491), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G119), .ZN(new_n696));
  OAI221_X1 g271(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n468), .C2(G107), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT83), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n701), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  OR2_X1    g280(.A1(G16), .A2(G24), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(G290), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n704), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n705), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n691), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n689), .A2(new_n690), .ZN(new_n713));
  OR4_X1    g288(.A1(KEYINPUT85), .A2(new_n711), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(KEYINPUT85), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n712), .A2(KEYINPUT85), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n715), .B(new_n717), .C1(new_n711), .C2(new_n713), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n693), .A2(G35), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G162), .B2(new_n693), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT93), .Z(new_n724));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G29), .B2(G32), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n483), .A2(G129), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT87), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n491), .A2(G141), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT26), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n732), .A2(new_n733), .B1(G105), .B2(new_n478), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n728), .A2(new_n729), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  MUX2_X1   g312(.A(new_n726), .B(new_n725), .S(new_n737), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT27), .B(G1996), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G19), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n543), .B2(G16), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT86), .B(G1341), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n724), .A2(new_n740), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n707), .A2(G20), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT23), .Z(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G299), .B2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1956), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n722), .B2(new_n721), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT94), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G21), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G168), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT89), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT90), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT25), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n491), .A2(G139), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n466), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n759), .B(new_n760), .C1(new_n468), .C2(new_n761), .ZN(new_n762));
  MUX2_X1   g337(.A(G33), .B(new_n762), .S(G29), .Z(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2072), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n755), .B2(new_n754), .ZN(new_n765));
  NOR2_X1   g340(.A1(G4), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n596), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n692), .A2(G26), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT28), .Z(new_n770));
  OAI221_X1 g345(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n468), .C2(G116), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G128), .ZN(new_n772));
  INV_X1    g347(.A(G140), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n771), .B(new_n772), .C1(new_n490), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n770), .B1(new_n774), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n768), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G11), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT91), .B(G28), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT30), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n779), .B1(new_n781), .B2(G29), .C1(new_n621), .C2(new_n692), .ZN(new_n782));
  INV_X1    g357(.A(G2084), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G34), .Z(new_n784));
  OAI22_X1  g359(.A1(new_n480), .A2(new_n736), .B1(new_n693), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n782), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(G5), .A2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT92), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G301), .B2(new_n707), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n787), .A2(G2084), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n786), .B(new_n792), .C1(new_n788), .C2(new_n791), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n693), .A2(G27), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G164), .B2(new_n693), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2078), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n757), .A2(new_n765), .A3(new_n778), .A4(new_n797), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n745), .A2(new_n751), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n714), .A2(new_n718), .A3(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  INV_X1    g376(.A(G55), .ZN(new_n802));
  INV_X1    g377(.A(G93), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n802), .A2(new_n511), .B1(new_n513), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n517), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G860), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT37), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n542), .B(new_n807), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT38), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n606), .A2(new_n601), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n808), .B1(new_n815), .B2(KEYINPUT39), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n810), .B1(new_n816), .B2(new_n817), .ZN(G145));
  NAND2_X1  g393(.A1(new_n498), .A2(new_n500), .ZN(new_n819));
  INV_X1    g394(.A(new_n495), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(new_n505), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n821), .A2(KEYINPUT95), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n501), .B2(new_n505), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n774), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n735), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n699), .B(new_n613), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n468), .A2(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(KEYINPUT98), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(KEYINPUT98), .B2(new_n831), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n491), .A2(G142), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT97), .B1(new_n483), .B2(G130), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n483), .A2(KEYINPUT97), .A3(G130), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n829), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n828), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n828), .B2(new_n839), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(KEYINPUT96), .B2(new_n762), .ZN(new_n843));
  INV_X1    g418(.A(new_n842), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n840), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(G162), .B(G160), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n621), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G37), .ZN(new_n851));
  INV_X1    g426(.A(new_n849), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n843), .A2(new_n846), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g432(.A1(G305), .A2(G303), .ZN(new_n858));
  OAI21_X1  g433(.A(G166), .B1(new_n578), .B2(new_n581), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n680), .A2(new_n681), .ZN(new_n861));
  NAND2_X1  g436(.A1(G290), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n682), .A2(new_n586), .A3(new_n584), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n858), .A2(new_n862), .A3(new_n863), .A4(new_n859), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n857), .B(KEYINPUT42), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT42), .ZN(new_n871));
  INV_X1    g446(.A(new_n867), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n859), .A2(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT101), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n872), .A2(new_n873), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT102), .B1(new_n877), .B2(new_n871), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n870), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G299), .B(new_n606), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(KEYINPUT100), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n883), .B2(KEYINPUT100), .ZN(new_n884));
  INV_X1    g459(.A(new_n811), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n604), .A2(KEYINPUT99), .A3(new_n607), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT99), .B1(new_n604), .B2(new_n607), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n811), .A3(new_n886), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n882), .A2(new_n884), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n889), .A2(new_n891), .ZN(new_n893));
  INV_X1    g468(.A(new_n880), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n879), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n896), .B1(new_n879), .B2(new_n895), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n879), .A2(new_n895), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n856), .B1(new_n900), .B2(new_n588), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n879), .A2(new_n895), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n879), .A2(new_n895), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n902), .B1(new_n903), .B2(new_n896), .ZN(new_n904));
  OAI211_X1 g479(.A(KEYINPUT104), .B(G868), .C1(new_n904), .C2(new_n897), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n588), .B1(new_n804), .B2(new_n806), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(G295));
  NAND3_X1  g482(.A1(new_n901), .A2(new_n905), .A3(new_n906), .ZN(G331));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n874), .A2(new_n875), .ZN(new_n910));
  AOI21_X1  g485(.A(G168), .B1(G301), .B2(KEYINPUT105), .ZN(new_n911));
  NOR2_X1   g486(.A1(G301), .A2(KEYINPUT105), .ZN(new_n912));
  MUX2_X1   g487(.A(new_n911), .B(G168), .S(new_n912), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n811), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n894), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(KEYINPUT106), .A3(new_n894), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n914), .ZN(new_n920));
  INV_X1    g495(.A(new_n881), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n920), .B1(new_n921), .B2(new_n883), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n910), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n882), .A2(new_n884), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n910), .B(new_n915), .C1(new_n924), .C2(new_n914), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n851), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n915), .B1(new_n924), .B2(new_n914), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(new_n874), .A3(new_n875), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n929), .A2(new_n930), .A3(new_n851), .A4(new_n925), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n909), .B1(new_n927), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n923), .B2(new_n926), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n929), .A2(KEYINPUT43), .A3(new_n851), .A4(new_n925), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n909), .B2(new_n935), .ZN(G397));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n823), .A2(new_n937), .A3(new_n825), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n469), .A2(G40), .A3(new_n479), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n942), .A2(new_n705), .A3(new_n586), .A4(new_n584), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT48), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n774), .B(new_n776), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT107), .ZN(new_n947));
  INV_X1    g522(.A(G1996), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n735), .B(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n700), .A2(new_n703), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n700), .A2(new_n703), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(new_n949), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n942), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n944), .B2(new_n943), .ZN(new_n956));
  INV_X1    g531(.A(new_n735), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n947), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n942), .B(new_n948), .C1(KEYINPUT126), .C2(KEYINPUT46), .ZN(new_n959));
  NAND2_X1  g534(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n960));
  OAI22_X1  g535(.A1(new_n958), .A2(new_n954), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n963));
  XOR2_X1   g538(.A(new_n962), .B(new_n963), .Z(new_n964));
  NAND2_X1  g539(.A1(new_n947), .A2(new_n949), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n965), .A2(new_n951), .B1(G2067), .B2(new_n774), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n956), .B(new_n964), .C1(new_n942), .C2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT62), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n937), .B1(new_n501), .B2(new_n505), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n939), .ZN(new_n970));
  INV_X1    g545(.A(new_n941), .ZN(new_n971));
  OAI211_X1 g546(.A(KEYINPUT45), .B(new_n937), .C1(new_n501), .C2(new_n505), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n755), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n941), .B1(new_n969), .B2(KEYINPUT50), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n821), .A2(new_n822), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n977), .A4(new_n937), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n977), .B(new_n937), .C1(new_n501), .C2(new_n505), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n975), .A2(new_n978), .A3(new_n783), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n974), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(KEYINPUT114), .B(G8), .Z(new_n984));
  NOR2_X1   g559(.A1(G168), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(G8), .ZN(new_n988));
  INV_X1    g563(.A(new_n985), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n984), .ZN(new_n991));
  AOI211_X1 g566(.A(KEYINPUT51), .B(new_n985), .C1(new_n983), .C2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n968), .B(new_n986), .C1(new_n990), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n823), .A2(new_n825), .A3(KEYINPUT45), .A4(new_n937), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n969), .A2(new_n996), .A3(new_n939), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n969), .B2(new_n939), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n971), .B(new_n995), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n994), .B1(new_n999), .B2(G2078), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT121), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1002), .B(new_n994), .C1(new_n999), .C2(G2078), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G2078), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n970), .A2(new_n1005), .A3(new_n971), .A4(new_n972), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT120), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n941), .B1(new_n969), .B2(new_n939), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n1005), .A4(new_n972), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(KEYINPUT53), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n975), .A2(new_n978), .A3(new_n981), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n788), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G301), .B1(new_n1004), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n993), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n995), .A2(new_n971), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n970), .A2(KEYINPUT108), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n969), .A2(new_n996), .A3(new_n939), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1971), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(KEYINPUT110), .B(G2090), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1012), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1018), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT113), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OR3_X1    g609(.A1(new_n1028), .A2(KEYINPUT112), .A3(new_n1029), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT112), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1971), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n999), .A2(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n975), .A2(new_n978), .A3(new_n981), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1024), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1041), .A3(KEYINPUT111), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1027), .A2(G8), .A3(new_n1037), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1037), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n975), .A2(new_n979), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n1025), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n991), .B1(new_n1023), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n969), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n971), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n991), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1052), .B(new_n1054), .C1(new_n1053), .C2(new_n861), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n579), .B(G1981), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1056), .A2(KEYINPUT49), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(KEYINPUT49), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1052), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n861), .A2(new_n1053), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT52), .B1(new_n1051), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1055), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1043), .A2(new_n1048), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT125), .B1(new_n1017), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1043), .A2(new_n1048), .A3(new_n1063), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1016), .A4(new_n993), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n988), .A2(new_n989), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT51), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n983), .A2(new_n991), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(new_n987), .A3(new_n989), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1070), .A2(new_n1072), .B1(new_n985), .B2(new_n983), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1073), .A2(new_n968), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1065), .A2(new_n1068), .A3(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1059), .A2(new_n1053), .A3(new_n678), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n577), .A2(G1981), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1052), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1043), .B2(new_n1062), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT63), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n983), .A2(G168), .A3(new_n991), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1080), .B1(new_n1064), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1027), .A2(G8), .A3(new_n1042), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n1044), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1081), .A2(new_n1080), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1043), .A3(new_n1063), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1079), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1075), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1012), .A2(KEYINPUT122), .A3(new_n788), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT122), .B1(new_n1012), .B2(new_n788), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1005), .A2(KEYINPUT53), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n941), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n469), .A2(KEYINPUT123), .A3(new_n479), .A4(G40), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n940), .A2(new_n995), .A3(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1090), .A2(new_n1091), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1019), .A2(new_n1005), .A3(new_n1022), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1002), .B1(new_n1099), .B2(new_n994), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1003), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1089), .B1(new_n1102), .B2(G171), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n1104));
  AND4_X1   g679(.A1(new_n1104), .A2(new_n1004), .A3(G301), .A4(new_n1015), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1014), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n1106), .B2(G301), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1103), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1102), .A2(G171), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1089), .B1(new_n1109), .B2(new_n1016), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1064), .A2(new_n1073), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n556), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(KEYINPUT57), .A4(new_n564), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n562), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n564), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n556), .B1(new_n558), .B2(new_n560), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1117), .B(new_n1118), .C1(KEYINPUT57), .C2(new_n1119), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT56), .B(G2072), .Z(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1019), .A2(new_n1022), .A3(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT115), .B(G1956), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1045), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1120), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI22_X1  g701(.A1(new_n1040), .A2(G1348), .B1(G2067), .B2(new_n1050), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1127), .A2(new_n596), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1129), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(new_n1126), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT61), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1050), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n999), .A2(G1996), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1138), .A2(new_n1139), .A3(new_n543), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1138), .B2(new_n543), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1131), .B(new_n1144), .C1(new_n1132), .C2(new_n1126), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1134), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1127), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1127), .B(new_n596), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1147), .B1(new_n1148), .B2(KEYINPUT60), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1142), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(KEYINPUT59), .A3(new_n1140), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1130), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1112), .B1(KEYINPUT119), .B2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1153), .A2(KEYINPUT119), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1088), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(G290), .B(new_n705), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n954), .B1(new_n953), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n967), .B1(new_n1156), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g734(.A1(G227), .A2(G229), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n854), .A2(G319), .A3(new_n639), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g736(.A1(new_n1162), .A2(new_n935), .ZN(G308));
  INV_X1    g737(.A(G308), .ZN(G225));
endmodule


