//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT77), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT77), .A2(G107), .ZN(new_n193));
  AOI21_X1  g007(.A(G104), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G107), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(KEYINPUT3), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n192), .A3(new_n193), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G107), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(new_n195), .B2(G107), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT68), .B1(new_n205), .B2(G119), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n207));
  INV_X1    g021(.A(G119), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G116), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n206), .A2(new_n209), .B1(new_n205), .B2(G119), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT2), .B(G113), .Z(new_n211));
  AND2_X1   g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n204), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(KEYINPUT5), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n205), .A2(KEYINPUT5), .A3(G119), .ZN(new_n215));
  INV_X1    g029(.A(G113), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT84), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G104), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT77), .A2(G107), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT77), .A2(G107), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n202), .A2(new_n201), .ZN(new_n228));
  OAI211_X1 g042(.A(G101), .B(new_n222), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n199), .A2(new_n201), .A3(new_n202), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n232), .A2(KEYINPUT79), .A3(G101), .A4(new_n222), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n235));
  INV_X1    g049(.A(new_n228), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n200), .B1(new_n236), .B2(new_n199), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n210), .A2(new_n211), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n235), .A2(new_n237), .B1(new_n212), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n221), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n203), .A2(KEYINPUT4), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n232), .A2(G101), .ZN(new_n242));
  INV_X1    g056(.A(new_n238), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n210), .A2(new_n211), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n231), .A2(new_n233), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(KEYINPUT84), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n220), .B1(new_n240), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n189), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT0), .B(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT0), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT0), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G128), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n261), .A2(new_n266), .A3(KEYINPUT64), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n264), .A2(new_n262), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n258), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n252), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n261), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT1), .B1(new_n256), .B2(G146), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n255), .A2(KEYINPUT67), .A3(KEYINPUT1), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(G128), .A3(new_n277), .ZN(new_n278));
  AOI211_X1 g092(.A(G125), .B(new_n273), .C1(new_n278), .C2(new_n261), .ZN(new_n279));
  OAI211_X1 g093(.A(G224), .B(new_n251), .C1(new_n271), .C2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n273), .B1(new_n278), .B2(new_n261), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n252), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n251), .A2(G224), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n260), .A2(new_n267), .B1(new_n258), .B2(new_n269), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n282), .B(new_n283), .C1(new_n252), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n234), .A2(new_n221), .A3(new_n239), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT84), .B1(new_n245), .B2(new_n246), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n219), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n187), .A2(new_n249), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n189), .B1(new_n290), .B2(new_n188), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n250), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n248), .A2(new_n187), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT7), .B1(new_n251), .B2(G224), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n280), .B2(new_n285), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n271), .B2(new_n279), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT86), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n214), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n210), .A2(KEYINPUT86), .A3(KEYINPUT5), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n217), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n218), .A2(new_n244), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n301), .A2(new_n213), .B1(new_n302), .B2(new_n204), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n187), .B(KEYINPUT8), .Z(new_n304));
  OAI21_X1  g118(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n296), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n294), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n293), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(new_n307), .A3(new_n309), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(KEYINPUT87), .A3(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n312), .A2(KEYINPUT87), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G140), .B1(new_n252), .B2(KEYINPUT71), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n252), .A2(G140), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT72), .A4(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n254), .ZN(new_n330));
  NOR2_X1   g144(.A1(G237), .A2(G953), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G214), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT88), .A3(G143), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT88), .A2(G143), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT88), .A2(G143), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(G214), .A3(new_n331), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT17), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n333), .A2(G131), .A3(new_n336), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n341), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n327), .A2(G146), .A3(new_n328), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n330), .A2(new_n342), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT18), .A2(G131), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n333), .A2(new_n347), .A3(new_n336), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n347), .B1(new_n333), .B2(new_n336), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n254), .B1(new_n319), .B2(new_n322), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(KEYINPUT89), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n254), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n351), .B2(KEYINPUT89), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n349), .A2(new_n350), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n346), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G113), .B(G122), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(new_n195), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n357), .B(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G475), .B1(new_n360), .B2(G902), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT19), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n321), .A2(G125), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n326), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT19), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n367), .A2(new_n254), .B1(new_n339), .B2(new_n341), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n352), .A2(new_n355), .ZN(new_n369));
  INV_X1    g183(.A(new_n350), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n348), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n368), .A2(new_n345), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT90), .B1(new_n372), .B2(new_n359), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n339), .A2(new_n341), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(G146), .B2(new_n366), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n327), .A2(G146), .A3(new_n328), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n356), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT90), .ZN(new_n378));
  INV_X1    g192(.A(new_n359), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n346), .A2(new_n359), .A3(new_n356), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n373), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n383));
  NOR2_X1   g197(.A1(G475), .A2(G902), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n361), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n251), .A2(G952), .ZN(new_n388));
  INV_X1    g202(.A(G234), .ZN(new_n389));
  INV_X1    g203(.A(G237), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G902), .ZN(new_n393));
  AOI211_X1 g207(.A(new_n393), .B(new_n251), .C1(G234), .C2(G237), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT21), .B(G898), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n205), .A2(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT14), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n205), .B2(G122), .ZN(new_n400));
  INV_X1    g214(.A(G122), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT91), .A3(G116), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G107), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n225), .A2(new_n226), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n406), .A3(new_n397), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT93), .B1(new_n262), .B2(G143), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n256), .A3(G128), .ZN(new_n411));
  AOI22_X1  g225(.A1(new_n409), .A2(new_n411), .B1(new_n262), .B2(G143), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(G134), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT13), .B1(new_n262), .B2(G143), .ZN(new_n416));
  INV_X1    g230(.A(G134), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n412), .B(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT92), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n406), .B1(new_n403), .B2(new_n397), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(new_n407), .ZN(new_n423));
  INV_X1    g237(.A(new_n407), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n424), .A2(KEYINPUT92), .A3(new_n421), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n419), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT9), .B(G234), .ZN(new_n427));
  INV_X1    g241(.A(G217), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(G953), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n415), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n429), .B1(new_n415), .B2(new_n426), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n393), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  OAI221_X1 g250(.A(new_n393), .B1(KEYINPUT15), .B2(new_n434), .C1(new_n431), .C2(new_n432), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n387), .A2(new_n396), .A3(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  INV_X1    g254(.A(G227), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n440), .B(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n262), .B1(new_n274), .B2(KEYINPUT80), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n255), .A2(new_n445), .A3(KEYINPUT1), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n258), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n203), .B(new_n197), .C1(new_n447), .C2(new_n273), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n197), .A2(new_n203), .A3(KEYINPUT10), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n278), .A2(new_n261), .ZN(new_n451));
  INV_X1    g265(.A(new_n273), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n246), .A2(new_n284), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n457));
  INV_X1    g271(.A(G137), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G134), .ZN(new_n459));
  NOR2_X1   g273(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(G134), .A3(new_n458), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n458), .A2(G134), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n461), .A2(new_n338), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g281(.A(new_n459), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n464), .B1(new_n468), .B2(new_n462), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(new_n470), .A3(new_n338), .A4(new_n461), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n461), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n467), .A2(new_n471), .B1(G131), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n454), .A2(new_n456), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n454), .B2(new_n456), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n443), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n454), .A2(new_n456), .A3(new_n473), .ZN(new_n479));
  INV_X1    g293(.A(new_n443), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n281), .A2(new_n204), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n281), .A2(new_n204), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n448), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n471), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n472), .A2(G131), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n486), .A2(KEYINPUT81), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT12), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n473), .A2(KEYINPUT12), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n486), .A2(KEYINPUT81), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n481), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(KEYINPUT83), .B(new_n443), .C1(new_n474), .C2(new_n475), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n478), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G469), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n393), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n479), .A3(new_n493), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n443), .ZN(new_n500));
  INV_X1    g314(.A(new_n475), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n481), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(G469), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(G469), .A2(G902), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G221), .B1(new_n427), .B2(G902), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n439), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G472), .A2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT32), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n331), .A2(G210), .ZN(new_n512));
  XOR2_X1   g326(.A(new_n512), .B(KEYINPUT27), .Z(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT26), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n200), .ZN(new_n515));
  OAI21_X1  g329(.A(G131), .B1(new_n468), .B2(new_n464), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n487), .A2(new_n453), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n267), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT64), .B1(new_n261), .B2(new_n266), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n270), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n487), .B2(new_n488), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n212), .A2(new_n238), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n489), .A2(new_n284), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n487), .A2(new_n453), .A3(new_n516), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT28), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n522), .A3(new_n526), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n515), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n517), .B2(new_n521), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n526), .B(KEYINPUT30), .C1(new_n473), .C2(new_n520), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n523), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT69), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT69), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n535), .A2(new_n539), .A3(new_n523), .A4(new_n536), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n515), .A2(new_n529), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n533), .B1(new_n544), .B2(KEYINPUT31), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n542), .B1(new_n538), .B2(new_n540), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT31), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n511), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n523), .B1(new_n517), .B2(new_n521), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n530), .B1(new_n550), .B2(new_n529), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n517), .A2(new_n521), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT28), .B1(new_n552), .B2(new_n522), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n514), .B(G101), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(G902), .B1(new_n555), .B2(KEYINPUT29), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n515), .B1(new_n541), .B2(new_n529), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n528), .A2(new_n515), .A3(new_n531), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n556), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G472), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n544), .A2(KEYINPUT31), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n532), .B1(new_n546), .B2(new_n547), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n509), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n549), .B(new_n562), .C1(KEYINPUT32), .C2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n251), .A2(G221), .A3(G234), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT22), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(G137), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT23), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(new_n208), .B2(G128), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n208), .A2(G128), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G110), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n262), .A2(G119), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n573), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT24), .B(G110), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n575), .A2(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n330), .B2(new_n345), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n572), .A2(new_n574), .A3(new_n576), .A4(new_n573), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n582), .A2(KEYINPUT73), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n579), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(KEYINPUT73), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n586), .A2(new_n345), .A3(new_n354), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n570), .B1(new_n581), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n586), .A2(new_n345), .A3(new_n354), .ZN(new_n589));
  AOI21_X1  g403(.A(G146), .B1(new_n327), .B2(new_n328), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n376), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n589), .B(new_n569), .C1(new_n591), .C2(new_n580), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G217), .B1(new_n389), .B2(G902), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT70), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(G902), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT75), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n598), .A2(KEYINPUT76), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n588), .A2(new_n393), .A3(new_n592), .ZN(new_n600));
  AND2_X1   g414(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n588), .A2(new_n592), .A3(new_n393), .A4(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n602), .A2(new_n605), .A3(new_n595), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n598), .A2(KEYINPUT76), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n599), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n318), .A2(new_n507), .A3(new_n566), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT94), .B(G101), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G3));
  NAND2_X1  g426(.A1(new_n563), .A2(new_n564), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n508), .ZN(new_n614));
  INV_X1    g428(.A(G472), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n563), .B2(new_n564), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n614), .B(new_n609), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n505), .A2(new_n506), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n396), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  OR3_X1    g435(.A1(new_n431), .A2(new_n621), .A3(new_n432), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n621), .B1(new_n431), .B2(new_n432), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n434), .A2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT95), .B(G478), .Z(new_n626));
  NAND2_X1  g440(.A1(new_n433), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n387), .A2(new_n620), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n311), .A2(new_n312), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(KEYINPUT96), .A3(new_n630), .A4(new_n316), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n293), .A2(new_n307), .A3(new_n309), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n309), .B1(new_n293), .B2(new_n307), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n316), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n387), .A2(new_n628), .A3(new_n620), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n619), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  OAI211_X1 g455(.A(new_n438), .B(new_n361), .C1(new_n385), .C2(new_n386), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n635), .A2(new_n396), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n619), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT35), .B(G107), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  OAI21_X1  g460(.A(new_n393), .B1(new_n545), .B2(new_n548), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n565), .B1(new_n647), .B2(G472), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n589), .B1(new_n591), .B2(new_n580), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n570), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n597), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n606), .A2(KEYINPUT97), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT97), .B1(new_n606), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n649), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n606), .A2(new_n653), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n606), .A2(new_n653), .A3(KEYINPUT97), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(KEYINPUT98), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n318), .A2(new_n507), .A3(new_n648), .A4(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  INV_X1    g479(.A(new_n387), .ZN(new_n666));
  INV_X1    g480(.A(new_n394), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT99), .B(G900), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n392), .B1(new_n670), .B2(KEYINPUT100), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(KEYINPUT100), .B2(new_n670), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n666), .A2(new_n438), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n635), .ZN(new_n674));
  INV_X1    g488(.A(new_n618), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n566), .A2(new_n674), .A3(new_n662), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  OAI21_X1  g491(.A(new_n549), .B1(new_n565), .B2(KEYINPUT32), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n524), .A2(new_n527), .ZN(new_n679));
  AOI21_X1  g493(.A(G902), .B1(new_n679), .B2(new_n554), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n524), .B1(new_n538), .B2(new_n540), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n680), .B1(new_n681), .B2(new_n554), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n682), .A2(KEYINPUT101), .A3(G472), .ZN(new_n683));
  AOI21_X1  g497(.A(KEYINPUT101), .B1(new_n682), .B2(G472), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(KEYINPUT102), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n672), .B(KEYINPUT103), .Z(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT39), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n675), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT40), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n315), .B(KEYINPUT38), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n659), .A2(new_n660), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n387), .A2(new_n438), .ZN(new_n698));
  NOR4_X1   g512(.A1(new_n696), .A2(new_n317), .A3(new_n697), .A4(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n690), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n690), .A2(KEYINPUT104), .A3(new_n695), .A4(new_n699), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n256), .ZN(G45));
  NAND3_X1  g519(.A1(new_n387), .A2(new_n628), .A3(new_n672), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n635), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n566), .A2(new_n662), .A3(new_n675), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NAND2_X1  g523(.A1(new_n614), .A2(new_n510), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n613), .A2(new_n511), .B1(new_n561), .B2(G472), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n608), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n496), .A2(new_n393), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n506), .A3(new_n498), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n712), .A2(new_n638), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n566), .A2(new_n643), .A3(new_n609), .A4(new_n716), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n712), .A2(KEYINPUT105), .A3(new_n643), .A4(new_n716), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR2_X1   g539(.A1(new_n715), .A2(new_n635), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n566), .A2(new_n726), .A3(new_n662), .A4(new_n439), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NOR2_X1   g542(.A1(new_n715), .A2(new_n396), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n635), .A2(new_n698), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n648), .A3(new_n609), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND4_X1  g546(.A1(new_n648), .A2(new_n697), .A3(new_n707), .A4(new_n716), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  NAND2_X1  g548(.A1(new_n315), .A2(new_n316), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n618), .ZN(new_n736));
  INV_X1    g550(.A(new_n706), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n712), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT42), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n736), .A2(new_n712), .A3(new_n740), .A4(new_n737), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  INV_X1    g557(.A(new_n673), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n736), .A2(new_n712), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT106), .B(G134), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G36));
  AND2_X1   g561(.A1(new_n500), .A2(new_n502), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n748), .A2(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n750), .B(G469), .C1(KEYINPUT45), .C2(new_n748), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n504), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT46), .B(new_n504), .C1(new_n751), .C2(new_n752), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n498), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n506), .A3(new_n693), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT43), .B1(new_n666), .B2(new_n628), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n387), .A2(KEYINPUT108), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n387), .A2(KEYINPUT108), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n628), .A2(KEYINPUT43), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT109), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n760), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n616), .A2(new_n615), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n697), .B1(new_n770), .B2(new_n565), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(new_n774), .A3(KEYINPUT44), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n735), .B(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n774), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n759), .A2(new_n775), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  NAND2_X1  g595(.A1(new_n757), .A2(new_n506), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n757), .A2(new_n784), .A3(new_n506), .ZN(new_n785));
  INV_X1    g599(.A(new_n566), .ZN(new_n786));
  INV_X1    g600(.A(new_n735), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n706), .A2(new_n609), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n783), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G140), .ZN(G42));
  AND2_X1   g606(.A1(new_n714), .A2(new_n498), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n761), .A2(new_n762), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n609), .A2(new_n316), .A3(new_n506), .A4(new_n628), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n689), .A2(new_n696), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n783), .A2(new_n785), .ZN(new_n801));
  INV_X1    g615(.A(new_n506), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n793), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n768), .A2(new_n391), .A3(new_n617), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n776), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n715), .A2(new_n316), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n805), .A2(new_n696), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT50), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n735), .A2(new_n608), .A3(new_n391), .A4(new_n715), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n689), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n387), .A3(new_n628), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n768), .A2(new_n391), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n735), .A2(new_n715), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n648), .A2(new_n813), .A3(new_n697), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n809), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n387), .A2(new_n628), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n388), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n813), .A2(new_n712), .A3(new_n814), .ZN(new_n820));
  NAND2_X1  g634(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n821));
  OR2_X1    g635(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n820), .B2(new_n821), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n819), .B(new_n824), .C1(new_n726), .C2(new_n805), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n809), .A2(new_n816), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n805), .A2(new_n776), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n803), .B(KEYINPUT115), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n801), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n817), .B(new_n825), .C1(new_n830), .C2(KEYINPUT51), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n676), .A2(new_n708), .A3(new_n733), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n635), .A2(new_n657), .A3(new_n698), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n505), .A2(new_n506), .A3(new_n672), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n834), .B(new_n835), .C1(new_n678), .C2(new_n685), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(KEYINPUT113), .A3(KEYINPUT52), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n676), .A2(new_n708), .A3(new_n836), .A4(new_n733), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n656), .A2(new_n661), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n710), .B2(new_n711), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n618), .A2(new_n673), .A3(new_n635), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n618), .A2(new_n635), .A3(new_n706), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT114), .A3(new_n733), .A4(new_n836), .ZN(new_n850));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n629), .A2(new_n313), .A3(new_n316), .A4(new_n314), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n313), .A2(new_n314), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT112), .A3(new_n316), .A4(new_n629), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n619), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(new_n610), .A3(new_n727), .A4(new_n731), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n666), .A2(new_n620), .A3(new_n438), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n315), .A2(new_n860), .A3(new_n317), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n609), .A3(new_n675), .A4(new_n648), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n717), .A2(new_n862), .A3(new_n663), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n745), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n387), .A2(new_n438), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n566), .A2(new_n866), .A3(new_n662), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n648), .A2(new_n697), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n867), .B1(new_n818), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n787), .A2(new_n835), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n864), .A2(new_n742), .A3(new_n871), .A4(new_n724), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n832), .B1(new_n852), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n844), .A2(new_n850), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n840), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n850), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n717), .A2(new_n862), .A3(new_n663), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n610), .A2(new_n727), .A3(new_n731), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n724), .A3(new_n858), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n869), .A2(new_n870), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n739), .A3(new_n741), .A4(new_n745), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n877), .A2(KEYINPUT53), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n873), .A2(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n852), .A2(new_n872), .A3(new_n832), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT53), .B1(new_n877), .B2(new_n883), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  MUX2_X1   g703(.A(new_n885), .B(new_n888), .S(new_n889), .Z(new_n890));
  NOR2_X1   g704(.A1(new_n831), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n800), .B1(new_n891), .B2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n251), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n896));
  OAI211_X1 g710(.A(G210), .B(G902), .C1(new_n886), .C2(new_n887), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n250), .A2(new_n292), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT117), .Z(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT55), .Z(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n286), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(KEYINPUT56), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(G210), .A2(G902), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n850), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n851), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n832), .B1(new_n906), .B2(new_n872), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n883), .B(KEYINPUT53), .C1(new_n851), .C2(new_n842), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n902), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n895), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g729(.A(KEYINPUT118), .B(new_n904), .C1(new_n907), .C2(new_n908), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n901), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT119), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT119), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n919), .B(new_n901), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n912), .B1(new_n918), .B2(new_n920), .ZN(G51));
  NAND2_X1  g735(.A1(new_n907), .A2(new_n908), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n889), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n504), .B(KEYINPUT57), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n496), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n888), .A2(new_n393), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n751), .A2(new_n752), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n894), .B1(new_n925), .B2(new_n928), .ZN(G54));
  NAND3_X1  g743(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .ZN(new_n930));
  INV_X1    g744(.A(new_n382), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n894), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n926), .A2(KEYINPUT58), .A3(G475), .A4(new_n382), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G60));
  AND2_X1   g748(.A1(new_n622), .A2(new_n623), .ZN(new_n935));
  XNOR2_X1  g749(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n434), .A2(new_n393), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n935), .B1(new_n890), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n935), .A2(new_n939), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n895), .B1(new_n923), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n652), .B(new_n946), .C1(new_n886), .C2(new_n887), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n947), .A2(KEYINPUT61), .A3(new_n895), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n945), .B1(new_n907), .B2(new_n908), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n593), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n950), .A2(KEYINPUT123), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n949), .A2(new_n952), .A3(new_n593), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n948), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n947), .B(new_n895), .C1(new_n593), .C2(new_n949), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(KEYINPUT122), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(KEYINPUT122), .B1(new_n955), .B2(new_n956), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G66));
  NAND2_X1  g773(.A1(G224), .A2(G953), .ZN(new_n960));
  OAI22_X1  g774(.A1(new_n880), .A2(G953), .B1(new_n395), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n899), .B1(G898), .B2(new_n251), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT124), .Z(new_n963));
  XNOR2_X1  g777(.A(new_n961), .B(new_n963), .ZN(G69));
  NAND3_X1  g778(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n535), .A2(new_n536), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n367), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n783), .A2(new_n785), .A3(new_n790), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n702), .A2(new_n703), .A3(new_n833), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(KEYINPUT62), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n702), .A2(new_n703), .A3(new_n971), .A4(new_n833), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n818), .A2(new_n642), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n712), .A2(new_n787), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n975), .A2(new_n694), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT125), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n780), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n251), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n965), .B(new_n967), .C1(new_n973), .C2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n779), .A2(new_n775), .A3(new_n776), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n712), .A2(new_n730), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n758), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT126), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n742), .A2(new_n745), .A3(new_n833), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n984), .A2(new_n985), .A3(new_n791), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n791), .A2(new_n986), .ZN(new_n988));
  OAI21_X1  g802(.A(KEYINPUT126), .B1(new_n988), .B2(new_n983), .ZN(new_n989));
  AOI21_X1  g803(.A(G953), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n441), .A2(G900), .A3(G953), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n967), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n980), .B1(new_n990), .B2(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(new_n681), .A2(new_n554), .ZN(new_n994));
  INV_X1    g808(.A(new_n880), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n987), .A2(new_n989), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT127), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n994), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n681), .A2(new_n554), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n970), .A2(new_n978), .A3(new_n995), .A4(new_n972), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n999), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n544), .B1(new_n515), .B2(new_n681), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n885), .A2(new_n998), .A3(new_n1005), .ZN(new_n1006));
  NOR4_X1   g820(.A1(new_n1000), .A2(new_n1004), .A3(new_n1006), .A4(new_n894), .ZN(G57));
endmodule


