//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n868, new_n869, new_n870,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(G1gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT94), .ZN(new_n204));
  AOI21_X1  g003(.A(G8gat), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n203), .B(new_n207), .C1(new_n204), .C2(G8gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT92), .B(G29gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G36gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT15), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G43gat), .B(G50gat), .Z(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(G50gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G43gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n219), .B1(new_n221), .B2(KEYINPUT93), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n216), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n217), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n223), .A2(new_n218), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT17), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT17), .B1(new_n224), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n211), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n224), .A2(new_n209), .A3(new_n225), .A4(new_n210), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT18), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n228), .A2(KEYINPUT18), .A3(new_n229), .A4(new_n230), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n211), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n230), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n229), .B(KEYINPUT13), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n233), .A2(new_n234), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT90), .B(G197gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT11), .B(G169gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT12), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n240), .A2(KEYINPUT91), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n240), .B2(KEYINPUT91), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT80), .ZN(new_n251));
  INV_X1    g050(.A(G141gat), .ZN(new_n252));
  INV_X1    g051(.A(G148gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n254), .A2(KEYINPUT2), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G155gat), .B(G162gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G155gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(G162gat), .ZN(new_n260));
  INV_X1    g059(.A(G162gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(G155gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(G141gat), .B(G148gat), .ZN(new_n263));
  OAI221_X1 g062(.A(KEYINPUT80), .B1(new_n260), .B2(new_n262), .C1(new_n263), .C2(KEYINPUT2), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(KEYINPUT82), .A2(G155gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(KEYINPUT82), .A2(G155gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT2), .B1(new_n268), .B2(new_n261), .ZN(new_n269));
  INV_X1    g068(.A(new_n263), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n257), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT81), .B1(new_n260), .B2(new_n262), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n269), .A2(new_n270), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n265), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n265), .A2(new_n277), .A3(new_n274), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G127gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281));
  INV_X1    g080(.A(G127gat), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n281), .B1(new_n282), .B2(G134gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(new_n281), .A3(G127gat), .ZN(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G113gat), .ZN(new_n287));
  INV_X1    g086(.A(G113gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G120gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT1), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  XNOR2_X1  g093(.A(G127gat), .B(G134gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n276), .A2(new_n278), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n275), .B2(new_n297), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n272), .A2(new_n273), .A3(new_n270), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n302), .A2(new_n269), .B1(new_n258), .B2(new_n264), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n285), .A2(new_n292), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n304), .A2(new_n284), .B1(new_n294), .B2(new_n295), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT4), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n298), .A2(new_n299), .A3(new_n301), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n299), .ZN(new_n308));
  AND4_X1   g107(.A1(new_n265), .A2(new_n274), .A3(new_n293), .A4(new_n296), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n265), .A2(new_n274), .B1(new_n293), .B2(new_n296), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT5), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n301), .A2(new_n306), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n314), .A2(KEYINPUT5), .A3(new_n299), .A4(new_n298), .ZN(new_n315));
  XOR2_X1   g114(.A(G1gat), .B(G29gat), .Z(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G57gat), .B(G85gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n313), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT89), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n313), .A2(new_n315), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n320), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n327));
  NAND4_X1  g126(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT89), .A4(new_n321), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n322), .A2(new_n327), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n331), .A2(KEYINPUT77), .B1(G211gat), .B2(G218gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(KEYINPUT77), .B2(new_n331), .ZN(new_n333));
  XNOR2_X1  g132(.A(G197gat), .B(G204gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(G211gat), .B(G218gat), .Z(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n333), .B2(new_n334), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(new_n336), .ZN(new_n340));
  INV_X1    g139(.A(G226gat), .ZN(new_n341));
  INV_X1    g140(.A(G233gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(KEYINPUT29), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI22_X1  g152(.A1(new_n349), .A2(new_n350), .B1(KEYINPUT26), .B2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n349), .A2(new_n350), .ZN(new_n355));
  INV_X1    g154(.A(G183gat), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  OAI22_X1  g156(.A1(new_n354), .A2(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n356), .A2(KEYINPUT27), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT27), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G183gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT67), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n361), .B2(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n357), .A2(KEYINPUT28), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT27), .B(G183gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n369), .B1(new_n357), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n360), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n364), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n362), .A2(G183gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n356), .A2(KEYINPUT27), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT67), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n367), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n357), .ZN(new_n379));
  INV_X1    g178(.A(new_n369), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n378), .A2(KEYINPUT68), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n359), .A2(new_n372), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n347), .A2(KEYINPUT23), .ZN(new_n384));
  INV_X1    g183(.A(new_n346), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT23), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n353), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT64), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(G183gat), .B2(G190gat), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n384), .B(new_n387), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT65), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n384), .B1(new_n396), .B2(new_n346), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT25), .B1(new_n347), .B2(KEYINPUT23), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n385), .A2(KEYINPUT65), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n392), .A2(new_n388), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n383), .A2(KEYINPUT79), .A3(new_n403), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n345), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n404), .A2(new_n341), .A3(new_n342), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n340), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n343), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n337), .A2(new_n338), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n339), .A2(new_n336), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n404), .A2(new_n344), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND3_X1  g218(.A1(new_n410), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n329), .A2(new_n330), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n410), .A2(new_n416), .ZN(new_n424));
  INV_X1    g223(.A(new_n419), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n422), .B1(new_n410), .B2(new_n416), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT38), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT38), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n408), .A2(new_n409), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(new_n340), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n340), .A3(new_n415), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT37), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n419), .B1(new_n410), .B2(new_n416), .ZN(new_n434));
  OAI221_X1 g233(.A(new_n429), .B1(new_n431), .B2(new_n433), .C1(new_n434), .C2(new_n423), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n421), .A2(new_n428), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(G22gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT31), .B(G50gat), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(G228gat), .A2(G233gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n442), .B(KEYINPUT85), .Z(new_n443));
  AND3_X1   g242(.A1(new_n333), .A2(new_n338), .A3(new_n334), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n444), .A2(new_n339), .A3(KEYINPUT29), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n275), .B1(new_n445), .B2(KEYINPUT3), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT29), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n340), .B1(new_n278), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n448), .B2(KEYINPUT86), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450));
  AOI211_X1 g249(.A(new_n450), .B(new_n340), .C1(new_n447), .C2(new_n278), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n443), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT87), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n454), .B(new_n443), .C1(new_n449), .C2(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n340), .A2(new_n447), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n303), .B1(new_n457), .B2(new_n277), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n458), .A2(new_n448), .A3(new_n442), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n441), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  AOI211_X1 g260(.A(new_n440), .B(new_n459), .C1(new_n453), .C2(new_n455), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n439), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n303), .B2(new_n277), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n450), .B1(new_n464), .B2(new_n340), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n448), .A2(KEYINPUT86), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n446), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n454), .B1(new_n467), .B2(new_n443), .ZN(new_n468));
  INV_X1    g267(.A(new_n455), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n460), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n440), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n441), .A3(new_n460), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n438), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n463), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n297), .B1(new_n303), .B2(new_n277), .ZN(new_n476));
  INV_X1    g275(.A(new_n278), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n301), .B(new_n306), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n478), .A2(new_n479), .A3(new_n308), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n478), .B2(new_n308), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n277), .B1(new_n265), .B2(new_n274), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n477), .A2(new_n483), .A3(new_n305), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n301), .A2(new_n306), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n308), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT88), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(new_n479), .A3(new_n308), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n309), .A2(new_n310), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n475), .B1(new_n489), .B2(new_n299), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(new_n491), .A3(new_n320), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT40), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT40), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n482), .A2(new_n491), .A3(new_n494), .A4(new_n320), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OR3_X1    g295(.A1(new_n424), .A2(KEYINPUT30), .A3(new_n425), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n424), .A2(new_n425), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n420), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n324), .A2(new_n328), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n496), .A2(new_n497), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n436), .A2(new_n474), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n497), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n326), .A2(new_n322), .A3(new_n327), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n330), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n463), .A2(new_n473), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n378), .A2(KEYINPUT68), .A3(new_n381), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT68), .B1(new_n378), .B2(new_n381), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n509), .A2(new_n510), .A3(new_n358), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n393), .A2(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n305), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n383), .A2(new_n297), .A3(new_n403), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT34), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT34), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n515), .A2(new_n519), .A3(new_n516), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n513), .A2(G227gat), .A3(new_n514), .A4(G233gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT32), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT33), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(G15gat), .B(G43gat), .Z(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G71gat), .B(G99gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n522), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n521), .B(KEYINPUT32), .C1(new_n523), .C2(new_n529), .ZN(new_n532));
  AOI221_X4 g331(.A(KEYINPUT76), .B1(new_n518), .B2(new_n520), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n532), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n520), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n519), .B1(new_n515), .B2(new_n516), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(new_n531), .A3(new_n532), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT75), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n541), .A2(new_n531), .A3(KEYINPUT75), .A4(new_n532), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT36), .B1(new_n538), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n535), .A2(new_n536), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(KEYINPUT36), .A3(new_n542), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT74), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n502), .B(new_n508), .C1(new_n548), .C2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n533), .A2(new_n537), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(new_n546), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT35), .B1(new_n329), .B2(new_n330), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n554), .A2(new_n503), .A3(new_n474), .A4(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n463), .A2(new_n473), .A3(new_n549), .A4(new_n542), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT35), .B1(new_n557), .B2(new_n506), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n250), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT100), .ZN(new_n567));
  AND2_X1   g366(.A1(G99gat), .A2(G106gat), .ZN(new_n568));
  NOR2_X1   g367(.A1(G99gat), .A2(G106gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n572), .A2(KEYINPUT98), .B1(G85gat), .B2(G92gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n574), .A2(KEYINPUT99), .A3(KEYINPUT7), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT99), .B1(new_n574), .B2(KEYINPUT7), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n573), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G85gat), .A2(G92gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n574), .B2(KEYINPUT7), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n572), .B2(KEYINPUT98), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(KEYINPUT99), .A3(KEYINPUT7), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT8), .ZN(new_n585));
  OAI22_X1  g384(.A1(new_n568), .A2(new_n585), .B1(G85gat), .B2(G92gat), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n571), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  AOI211_X1 g387(.A(new_n570), .B(new_n586), .C1(new_n577), .C2(new_n583), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n235), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT17), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n590), .A2(new_n225), .A3(new_n224), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n567), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n590), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n226), .B2(new_n227), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(KEYINPUT100), .A3(new_n595), .A4(new_n596), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n566), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  INV_X1    g404(.A(new_n603), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n605), .B1(new_n604), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n565), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT101), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n564), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n583), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n587), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n570), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n584), .A2(new_n571), .A3(new_n587), .ZN(new_n620));
  NAND2_X1  g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  OR2_X1    g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT9), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G57gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G64gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(G64gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(KEYINPUT95), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n629), .A2(new_n625), .A3(G64gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n624), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G64gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(G57gat), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT9), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n621), .A3(new_n622), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n635), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n588), .B2(new_n589), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n644), .B1(new_n648), .B2(new_n641), .ZN(new_n649));
  AOI211_X1 g448(.A(KEYINPUT102), .B(new_n642), .C1(new_n646), .C2(new_n647), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n643), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n648), .A2(new_n641), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n643), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT21), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n638), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G231gat), .A2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G127gat), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n211), .B1(new_n660), .B2(new_n638), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(G183gat), .B(G211gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT96), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(new_n259), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n668), .B(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n666), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n615), .A2(new_n659), .A3(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n560), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n505), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g479(.A1(new_n560), .A2(new_n676), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n681), .B2(new_n503), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  INV_X1    g482(.A(new_n503), .ZN(new_n684));
  XOR2_X1   g483(.A(KEYINPUT16), .B(G8gat), .Z(new_n685));
  NAND3_X1  g484(.A1(new_n677), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n686), .A2(KEYINPUT103), .A3(new_n683), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT103), .B1(new_n686), .B2(new_n683), .ZN(new_n688));
  OAI221_X1 g487(.A(new_n682), .B1(new_n683), .B2(new_n686), .C1(new_n687), .C2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n677), .A2(new_n690), .A3(new_n554), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n548), .A2(new_n551), .ZN(new_n692));
  OAI21_X1  g491(.A(G15gat), .B1(new_n681), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(G1326gat));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n507), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT43), .B(G22gat), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n697), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n610), .A2(new_n614), .ZN(new_n701));
  INV_X1    g500(.A(new_n675), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(new_n702), .A3(new_n659), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n560), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n505), .A3(new_n215), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n702), .A2(new_n659), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n249), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n552), .A2(new_n559), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n615), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(KEYINPUT107), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n701), .B1(new_n552), .B2(new_n559), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n714), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n709), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n215), .B1(new_n721), .B2(new_n505), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n722), .ZN(G1328gat));
  NOR3_X1   g522(.A1(new_n704), .A2(G36gat), .A3(new_n503), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G36gat), .B1(new_n721), .B2(new_n503), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n726), .A2(KEYINPUT46), .A3(new_n727), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(G1329gat));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n692), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n720), .B2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n704), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n553), .A2(new_n546), .A3(G43gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT47), .B1(new_n739), .B2(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(new_n739), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n736), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n740), .B1(new_n736), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  NAND2_X1  g543(.A1(new_n717), .A2(new_n719), .ZN(new_n745));
  INV_X1    g544(.A(new_n709), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n507), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G50gat), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n737), .A2(new_n220), .A3(new_n507), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n749), .B1(new_n748), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1331gat));
  NAND3_X1  g552(.A1(new_n701), .A2(new_n250), .A3(new_n702), .ZN(new_n754));
  INV_X1    g553(.A(new_n659), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n710), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n505), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(new_n625), .ZN(G1332gat));
  NOR2_X1   g560(.A1(new_n759), .A2(new_n503), .ZN(new_n762));
  NOR2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  AND2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n759), .B2(new_n692), .ZN(new_n767));
  INV_X1    g566(.A(G71gat), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n554), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n759), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g569(.A(new_n770), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g570(.A1(new_n759), .A2(new_n474), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT111), .B(G78gat), .Z(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n702), .A2(new_n249), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT51), .B1(new_n718), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n710), .A2(new_n615), .A3(new_n775), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n781), .B2(new_n777), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n505), .A2(G85gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n659), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n775), .A2(new_n659), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(KEYINPUT112), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n745), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788), .B2(new_n505), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(G1336gat));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n710), .A2(new_n615), .B1(new_n715), .B2(new_n714), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n701), .B(new_n713), .C1(new_n552), .C2(new_n559), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n684), .B(new_n787), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n503), .A2(G92gat), .A3(new_n755), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n791), .B(new_n795), .C1(new_n782), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n779), .A2(new_n780), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n796), .B1(new_n799), .B2(new_n776), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n801), .B2(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  AOI211_X1 g602(.A(new_n803), .B(new_n791), .C1(new_n795), .C2(new_n800), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n798), .B1(new_n802), .B2(new_n804), .ZN(G1337gat));
  NOR3_X1   g604(.A1(new_n553), .A2(new_n546), .A3(G99gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n783), .A2(new_n659), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n788), .B2(new_n692), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1338gat));
  NOR3_X1   g608(.A1(new_n474), .A2(G106gat), .A3(new_n755), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n782), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n745), .A2(new_n507), .A3(new_n787), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n813), .A2(G106gat), .B1(new_n781), .B2(new_n810), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n812), .A2(new_n816), .B1(new_n817), .B2(new_n815), .ZN(G1339gat));
  INV_X1    g617(.A(new_n658), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n657), .A2(KEYINPUT102), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n648), .A2(new_n644), .A3(new_n641), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n648), .B2(new_n641), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n646), .A2(new_n642), .A3(new_n647), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n654), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n819), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n823), .A2(new_n826), .A3(KEYINPUT115), .A4(KEYINPUT55), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n238), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n236), .A2(new_n230), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT116), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n229), .B1(new_n228), .B2(new_n230), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n245), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n233), .A2(new_n234), .A3(new_n239), .A4(new_n246), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n615), .A2(new_n834), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n659), .A2(new_n841), .A3(new_n839), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT54), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n657), .A2(KEYINPUT54), .A3(new_n825), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n655), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n828), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n658), .A3(new_n830), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n846), .B1(new_n250), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n701), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n702), .B1(new_n845), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n754), .A2(new_n659), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n505), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(new_n503), .A3(new_n474), .A4(new_n554), .ZN(new_n858));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n250), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n557), .A2(new_n684), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT118), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n249), .A2(new_n288), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G1340gat));
  OAI21_X1  g663(.A(G120gat), .B1(new_n858), .B2(new_n755), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n659), .A2(new_n286), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n865), .B1(new_n862), .B2(new_n866), .ZN(G1341gat));
  INV_X1    g666(.A(new_n861), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n282), .A3(new_n702), .ZN(new_n869));
  OAI21_X1  g668(.A(G127gat), .B1(new_n858), .B2(new_n675), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(G1342gat));
  NAND3_X1  g670(.A1(new_n868), .A2(new_n279), .A3(new_n615), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n858), .B2(new_n701), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n684), .A2(new_n505), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n692), .A2(new_n877), .ZN(new_n878));
  AND4_X1   g677(.A1(new_n614), .A2(new_n834), .A3(new_n610), .A4(new_n844), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n851), .A2(KEYINPUT120), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n829), .A2(new_n833), .A3(new_n881), .A4(new_n830), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n249), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n846), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n879), .B1(new_n884), .B2(new_n701), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT121), .B1(new_n885), .B2(new_n702), .ZN(new_n886));
  INV_X1    g685(.A(new_n855), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n851), .A2(KEYINPUT120), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(new_n249), .A3(new_n882), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n615), .B1(new_n890), .B2(new_n846), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n888), .B(new_n675), .C1(new_n891), .C2(new_n879), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n887), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n507), .A2(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n897), .B1(new_n856), .B2(new_n474), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n878), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n252), .B1(new_n899), .B2(new_n249), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n735), .A2(new_n474), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n503), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n903), .A2(new_n252), .A3(new_n249), .A4(new_n857), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT122), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT58), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n878), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n675), .B1(new_n891), .B2(new_n879), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n855), .B1(new_n908), .B2(KEYINPUT121), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n894), .B1(new_n909), .B2(new_n892), .ZN(new_n910));
  INV_X1    g709(.A(new_n897), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n854), .A2(new_n855), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n912), .B2(new_n507), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n907), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G141gat), .B1(new_n914), .B2(new_n250), .ZN(new_n915));
  INV_X1    g714(.A(new_n905), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n906), .A2(new_n918), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n908), .A2(new_n887), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT57), .B1(new_n920), .B2(new_n507), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n856), .A2(new_n474), .A3(new_n897), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n659), .A3(new_n907), .ZN(new_n924));
  AND2_X1   g723(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n902), .A2(new_n505), .A3(new_n856), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n253), .A3(new_n659), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n253), .B1(new_n899), .B2(new_n659), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n926), .B(new_n928), .C1(KEYINPUT59), .C2(new_n929), .ZN(G1345gat));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n268), .A3(new_n702), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n675), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n268), .ZN(G1346gat));
  AOI21_X1  g732(.A(G162gat), .B1(new_n927), .B2(new_n615), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n701), .A2(new_n261), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n899), .B2(new_n935), .ZN(G1347gat));
  NOR4_X1   g735(.A1(new_n507), .A2(new_n553), .A3(new_n503), .A4(new_n546), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n912), .A2(new_n505), .A3(new_n937), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n938), .A2(new_n351), .A3(new_n250), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n505), .B1(new_n854), .B2(new_n855), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n557), .A2(new_n503), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT124), .Z(new_n944));
  NAND3_X1  g743(.A1(new_n942), .A2(new_n249), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n939), .B1(new_n945), .B2(new_n351), .ZN(G1348gat));
  OAI21_X1  g745(.A(G176gat), .B1(new_n938), .B2(new_n755), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n942), .A2(new_n944), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n659), .A2(new_n352), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(G1349gat));
  OAI21_X1  g749(.A(G183gat), .B1(new_n938), .B2(new_n675), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n702), .A2(new_n376), .A3(new_n373), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT60), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT60), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n955), .B(new_n951), .C1(new_n948), .C2(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1350gat));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n357), .A3(new_n615), .A4(new_n944), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n912), .A2(new_n505), .A3(new_n615), .A4(new_n937), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(G190gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n959), .B2(G190gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n958), .B(KEYINPUT125), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1351gat));
  NOR3_X1   g766(.A1(new_n735), .A2(new_n678), .A3(new_n503), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n923), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(G197gat), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(new_n250), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n901), .A2(new_n684), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n942), .A2(new_n249), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g773(.A1(new_n974), .A2(new_n970), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n971), .A2(new_n975), .ZN(G1352gat));
  XOR2_X1   g775(.A(KEYINPUT126), .B(G204gat), .Z(new_n977));
  OAI21_X1  g776(.A(new_n977), .B1(new_n969), .B2(new_n755), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n755), .A2(new_n977), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n942), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(G1353gat));
  NOR2_X1   g782(.A1(new_n675), .A2(G211gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n942), .A2(new_n973), .A3(new_n984), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n702), .B(new_n968), .C1(new_n921), .C2(new_n922), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(G1354gat));
  OAI21_X1  g788(.A(G218gat), .B1(new_n969), .B2(new_n701), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n701), .A2(G218gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n942), .A2(new_n973), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1355gat));
endmodule


