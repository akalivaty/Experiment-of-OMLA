//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G221), .A2(G218), .A3(G220), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g041(.A(KEYINPUT67), .B(G125), .C1(new_n462), .C2(new_n463), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n471), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n471), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G101), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g049(.A(G137), .B(new_n471), .C1(new_n462), .C2(new_n463), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n470), .A2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n481));
  INV_X1    g056(.A(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n471), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT69), .Z(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n483), .B2(new_n484), .ZN(new_n488));
  AOI211_X1 g063(.A(new_n480), .B(new_n487), .C1(G136), .C2(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n471), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n462), .B2(new_n463), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n463), .C2(new_n462), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G62), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n503), .A2(KEYINPUT71), .B1(G75), .B2(G543), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n501), .B2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n511), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n502), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n506), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n512), .A2(G51), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT72), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n523), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n522), .A2(new_n520), .A3(new_n524), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n519), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT5), .B(G543), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n515), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n527), .A2(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n512), .A2(G52), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n533), .B(KEYINPUT74), .C1(new_n534), .C2(new_n516), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OR2_X1    g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(G77), .A2(G543), .ZN(new_n540));
  OAI211_X1 g115(.A(KEYINPUT73), .B(G651), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  OAI21_X1  g116(.A(G651), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n535), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n515), .A2(new_n502), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G90), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT74), .B1(new_n547), .B2(new_n533), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n501), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n512), .A2(G43), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n546), .A2(G81), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT75), .Z(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n515), .A2(G91), .A3(new_n502), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT77), .B(G65), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n502), .A2(new_n563), .B1(G78), .B2(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(KEYINPUT76), .ZN(new_n567));
  AND3_X1   g142(.A1(new_n512), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n565), .B1(new_n512), .B2(new_n567), .ZN(new_n569));
  OAI221_X1 g144(.A(new_n562), .B1(new_n501), .B2(new_n564), .C1(new_n568), .C2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  OR2_X1    g146(.A1(new_n527), .A2(new_n531), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND2_X1  g148(.A1(new_n546), .A2(G87), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n512), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n528), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n512), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n546), .A2(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n501), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n512), .A2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n546), .A2(G85), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  XOR2_X1   g165(.A(KEYINPUT79), .B(G66), .Z(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n528), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  XNOR2_X1  g169(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n516), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n516), .B2(new_n594), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT80), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G284));
  XOR2_X1   g175(.A(G284), .B(KEYINPUT81), .Z(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n485), .A2(G123), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n471), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(G135), .B2(new_n488), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT83), .Z(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  XNOR2_X1  g193(.A(KEYINPUT3), .B(G2104), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n472), .B2(new_n473), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT13), .B(G2100), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT85), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT86), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n644), .B2(new_n647), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n652), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2096), .B(G2100), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT20), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n663), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  MUX2_X1   g243(.A(new_n667), .B(new_n668), .S(new_n661), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G23), .ZN(new_n679));
  AND3_X1   g254(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT33), .ZN(new_n682));
  INV_X1    g257(.A(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(G166), .A2(new_n678), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(G22), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(G1971), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(G1971), .ZN(new_n689));
  NOR2_X1   g264(.A1(G6), .A2(G16), .ZN(new_n690));
  INV_X1    g265(.A(G305), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XOR2_X1   g268(.A(new_n692), .B(new_n693), .Z(new_n694));
  NOR4_X1   g269(.A1(new_n684), .A2(new_n688), .A3(new_n689), .A4(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  INV_X1    g273(.A(G290), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(new_n678), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(new_n678), .B2(G24), .ZN(new_n701));
  INV_X1    g276(.A(G1986), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  AOI22_X1  g278(.A1(G119), .A2(new_n485), .B1(new_n488), .B2(G131), .ZN(new_n704));
  OAI21_X1  g279(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n707));
  OAI221_X1 g282(.A(G2104), .B1(G107), .B2(new_n471), .C1(new_n706), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G25), .B(new_n709), .S(G29), .Z(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n701), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(G1986), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n697), .A2(new_n698), .A3(new_n703), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT90), .B(KEYINPUT36), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT31), .B(G11), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT95), .B(G28), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(KEYINPUT30), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n720), .B2(KEYINPUT30), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n488), .A2(G141), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n485), .A2(G129), .ZN(new_n725));
  OAI21_X1  g300(.A(G105), .B1(new_n472), .B2(new_n473), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT26), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n724), .A2(new_n725), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(new_n722), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n722), .B2(G32), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n719), .B1(new_n721), .B2(new_n723), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n722), .A2(G26), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT91), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n488), .A2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n485), .A2(G128), .ZN(new_n740));
  OR2_X1    g315(.A1(G104), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n738), .B1(new_n744), .B2(new_n722), .ZN(new_n745));
  INV_X1    g320(.A(G2067), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n555), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G16), .B2(G19), .ZN(new_n749));
  INV_X1    g324(.A(G1341), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n735), .B(new_n751), .C1(new_n750), .C2(new_n749), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT24), .ZN(new_n753));
  INV_X1    g328(.A(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n753), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G160), .B2(new_n722), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(G2084), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n617), .A2(new_n722), .ZN(new_n759));
  NOR2_X1   g334(.A1(G27), .A2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G164), .B2(G29), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n759), .B1(G2078), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(G2078), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n733), .B2(new_n734), .ZN(new_n764));
  AND4_X1   g339(.A1(new_n752), .A2(new_n758), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G29), .A2(G33), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT92), .Z(new_n767));
  INV_X1    g342(.A(G127), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n483), .B2(new_n484), .ZN(new_n769));
  NAND2_X1  g344(.A1(G115), .A2(G2104), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(G2105), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G103), .A2(G2104), .ZN(new_n773));
  OAI21_X1  g348(.A(KEYINPUT93), .B1(new_n773), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n775), .A2(new_n471), .A3(G103), .A4(G2104), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n488), .A2(G139), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n774), .A2(new_n776), .A3(KEYINPUT25), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n772), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(G127), .B1(new_n462), .B2(new_n463), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(new_n770), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n786), .A2(G2105), .B1(G139), .B2(new_n488), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n774), .A2(KEYINPUT25), .A3(new_n776), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT25), .B1(new_n774), .B2(new_n776), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n790), .A3(KEYINPUT94), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n784), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n767), .B1(new_n792), .B2(new_n722), .ZN(new_n793));
  INV_X1    g368(.A(G2072), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(G2090), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n722), .A2(G35), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G162), .B2(new_n722), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT29), .Z(new_n799));
  OAI211_X1 g374(.A(new_n765), .B(new_n795), .C1(new_n796), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n678), .A2(G5), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G171), .B2(new_n678), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1961), .ZN(new_n803));
  NOR2_X1   g378(.A1(G168), .A2(new_n678), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n678), .B2(G21), .ZN(new_n805));
  INV_X1    g380(.A(G1966), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(new_n806), .B1(new_n757), .B2(G2084), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n806), .B2(new_n805), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n799), .A2(new_n796), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n678), .A2(G4), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n599), .B2(new_n678), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n793), .A2(new_n794), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n678), .A2(G20), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT23), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n603), .B2(new_n678), .ZN(new_n817));
  INV_X1    g392(.A(G1956), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n809), .A2(new_n813), .A3(new_n814), .A4(new_n819), .ZN(new_n820));
  NOR4_X1   g395(.A1(new_n800), .A2(new_n803), .A3(new_n808), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n718), .A2(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  AND3_X1   g398(.A1(new_n510), .A2(KEYINPUT6), .A3(G651), .ZN(new_n824));
  AOI21_X1  g399(.A(KEYINPUT6), .B1(new_n510), .B2(G651), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n502), .B(G93), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(G55), .B(G543), .C1(new_n824), .C2(new_n825), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT96), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n502), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(new_n501), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT97), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n826), .A2(new_n827), .A3(KEYINPUT96), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT96), .B1(new_n826), .B2(new_n827), .ZN(new_n837));
  OAI211_X1 g412(.A(KEYINPUT97), .B(new_n834), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n554), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n554), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n599), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n848));
  AOI21_X1  g423(.A(G860), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n848), .B2(new_n847), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT98), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n841), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n838), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT99), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n857), .ZN(G145));
  XOR2_X1   g433(.A(KEYINPUT105), .B(G37), .Z(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n617), .B(G160), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(G162), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n730), .B1(new_n792), .B2(new_n863), .ZN(new_n864));
  AOI211_X1 g439(.A(KEYINPUT101), .B(new_n731), .C1(new_n784), .C2(new_n791), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n744), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n782), .A2(new_n783), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT94), .B1(new_n787), .B2(new_n790), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n731), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n792), .A2(new_n863), .A3(new_n730), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n743), .A3(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n873));
  INV_X1    g448(.A(new_n499), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n498), .B1(new_n619), .B2(new_n495), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n873), .B1(new_n876), .B2(new_n493), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n497), .A2(new_n499), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n491), .A2(new_n492), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n485), .B2(G126), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT100), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n866), .A2(new_n872), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n883), .B1(new_n866), .B2(new_n872), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n622), .B(new_n709), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n485), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n471), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n488), .A2(G142), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(KEYINPUT102), .ZN(new_n893));
  OAI221_X1 g468(.A(new_n888), .B1(new_n889), .B2(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n887), .B(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n886), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n862), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n864), .A2(new_n865), .A3(new_n744), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n743), .B1(new_n870), .B2(new_n871), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n882), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n866), .A2(new_n872), .A3(new_n883), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT103), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n900), .A2(new_n895), .A3(new_n904), .A4(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n860), .B1(new_n897), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n903), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n903), .B2(new_n905), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n909), .A2(new_n910), .A3(new_n896), .ZN(new_n911));
  INV_X1    g486(.A(new_n862), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n907), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g489(.A(new_n844), .B(new_n608), .Z(new_n915));
  XNOR2_X1  g490(.A(new_n598), .B(G299), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT41), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n916), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(G288), .A2(KEYINPUT106), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(G288), .A2(KEYINPUT106), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n699), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(G290), .A3(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G303), .A2(G305), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  NAND2_X1  g505(.A1(G166), .A2(new_n691), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n928), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT107), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n921), .B(new_n938), .ZN(new_n939));
  MUX2_X1   g514(.A(new_n854), .B(new_n939), .S(G868), .Z(G295));
  MUX2_X1   g515(.A(new_n854), .B(new_n939), .S(G868), .Z(G331));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  OAI21_X1  g517(.A(G286), .B1(new_n545), .B2(new_n548), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n544), .A2(new_n541), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n533), .B1(new_n534), .B2(new_n516), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT74), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n944), .A2(G168), .A3(new_n947), .A4(new_n535), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n840), .A2(new_n843), .A3(new_n943), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n943), .A2(new_n948), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n555), .B1(new_n853), .B2(new_n838), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(new_n842), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n949), .A2(new_n920), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n844), .B2(new_n950), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n954), .B(new_n950), .C1(new_n951), .C2(new_n842), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n949), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n953), .B1(new_n958), .B2(new_n917), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n942), .B1(new_n959), .B2(new_n937), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n951), .A2(new_n950), .A3(new_n842), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(new_n916), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n952), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n952), .A2(KEYINPUT108), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n961), .B1(new_n964), .B2(new_n956), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n937), .B(new_n963), .C1(new_n965), .C2(new_n918), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n959), .A2(new_n968), .A3(new_n937), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n960), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n962), .B1(new_n955), .B2(new_n957), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n949), .A2(new_n952), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n918), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n937), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n860), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n968), .B1(new_n959), .B2(new_n937), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT43), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n971), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n980), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n970), .B2(new_n980), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(G397));
  OR3_X1    g562(.A1(new_n882), .A2(KEYINPUT110), .A3(G1384), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT110), .B1(new_n882), .B2(G1384), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT46), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n743), .B(new_n746), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n730), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT126), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT126), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n996), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(KEYINPUT47), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n993), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1005), .A2(G1986), .A3(G290), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT48), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n730), .B(G1996), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n998), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n704), .A2(new_n711), .A3(new_n708), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n709), .A2(new_n712), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1006), .A2(KEYINPUT48), .B1(new_n993), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1010), .B(KEYINPUT125), .ZN(new_n1015));
  AOI22_X1  g590(.A1(new_n1009), .A2(new_n1015), .B1(new_n746), .B2(new_n744), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1004), .B(new_n1014), .C1(new_n1005), .C2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT47), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n877), .A2(KEYINPUT45), .A3(new_n1020), .A4(new_n881), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n474), .A2(G40), .A3(new_n475), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(G2105), .B2(new_n469), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n876), .B2(new_n493), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n989), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1021), .A2(new_n1023), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n878), .B2(new_n880), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1023), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n818), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n568), .A2(new_n569), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n562), .B1(new_n564), .B2(new_n501), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1035), .B(new_n1036), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1038), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(KEYINPUT57), .C1(new_n569), .C2(new_n568), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1035), .B1(G299), .B2(new_n1036), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1034), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT117), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(KEYINPUT118), .A3(new_n1041), .A4(new_n1039), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1033), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n1023), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n992), .A2(new_n1024), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1051), .A2(new_n812), .B1(new_n1052), .B2(new_n746), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1048), .A2(new_n598), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1027), .A2(new_n1055), .A3(new_n1032), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(KEYINPUT119), .B2(new_n1033), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1054), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n812), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1023), .A2(new_n1028), .A3(new_n746), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT60), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1060), .B1(new_n1063), .B2(new_n598), .ZN(new_n1064));
  INV_X1    g639(.A(new_n598), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT121), .B(new_n1065), .C1(new_n1053), .C2(KEYINPUT60), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1053), .A2(KEYINPUT60), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1033), .A2(KEYINPUT119), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1070), .A2(new_n1056), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1033), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1057), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1033), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1076), .B2(new_n1048), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1064), .A2(new_n1066), .A3(KEYINPUT60), .A4(new_n1053), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1069), .A2(new_n1075), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1023), .B1(new_n1028), .B2(KEYINPUT45), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n994), .A3(new_n1021), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1052), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  AOI22_X1  g662(.A1(new_n1083), .A2(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1080), .B1(new_n1089), .B2(new_n555), .ZN(new_n1090));
  AOI211_X1 g665(.A(KEYINPUT59), .B(new_n554), .C1(new_n1085), .C2(new_n1088), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1059), .B1(new_n1079), .B2(new_n1092), .ZN(new_n1093));
  AOI211_X1 g668(.A(new_n989), .B(G1384), .C1(new_n878), .C2(new_n880), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n806), .B1(new_n1081), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(G2084), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1049), .A2(new_n1050), .A3(new_n1096), .A4(new_n1023), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G8), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G168), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1099), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1102), .A2(KEYINPUT51), .A3(new_n1100), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1102), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT122), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1100), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1105), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1104), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1098), .A2(new_n1108), .A3(G8), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1100), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1102), .A2(new_n1108), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT51), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(KEYINPUT123), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1101), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G303), .A2(G8), .ZN(new_n1120));
  XOR2_X1   g695(.A(new_n1120), .B(KEYINPUT55), .Z(new_n1121));
  AOI21_X1  g696(.A(G1971), .B1(new_n1082), .B2(new_n1021), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT111), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1122), .A2(new_n1123), .B1(G2090), .B2(new_n1051), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1121), .B(G8), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G2078), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1082), .A2(new_n1127), .A3(new_n1021), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n1129));
  INV_X1    g704(.A(G1961), .ZN(new_n1130));
  AOI22_X1  g705(.A1(new_n1128), .A2(new_n1129), .B1(new_n1130), .B2(new_n1051), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G171), .B(new_n1132), .ZN(new_n1133));
  AND4_X1   g708(.A1(KEYINPUT53), .A2(new_n1021), .A3(new_n1127), .A4(new_n1023), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n991), .B2(new_n1134), .ZN(new_n1135));
  OR4_X1    g710(.A1(new_n1129), .A2(new_n1081), .A3(G2078), .A4(new_n1094), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1131), .A2(new_n1135), .B1(new_n1137), .B2(new_n1133), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1052), .A2(new_n1099), .ZN(new_n1139));
  XNOR2_X1  g714(.A(G305), .B(G1981), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT49), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT112), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(KEYINPUT112), .A3(new_n1141), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(G288), .A2(new_n683), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1052), .A2(new_n1099), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT52), .B1(G288), .B2(new_n683), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT52), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1149), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1147), .A2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1120), .B(KEYINPUT55), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT114), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1051), .A2(G2090), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(new_n1122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G8), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1157), .A2(new_n1122), .A3(new_n1156), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1155), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND4_X1   g736(.A1(new_n1126), .A2(new_n1138), .A3(new_n1154), .A4(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1093), .A2(new_n1119), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n680), .A2(new_n683), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1147), .A2(new_n1164), .B1(G1981), .B2(G305), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1139), .B(KEYINPUT113), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1154), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1126), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1102), .A2(G168), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1170), .A2(KEYINPUT115), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(KEYINPUT115), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1173), .A2(new_n1161), .A3(new_n1126), .A4(new_n1154), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT63), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1177));
  OAI21_X1  g752(.A(G8), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1155), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1177), .A2(new_n1126), .A3(new_n1154), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1169), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(G301), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1182));
  AND4_X1   g757(.A1(new_n1126), .A2(new_n1161), .A3(new_n1182), .A4(new_n1154), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1101), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1103), .B1(new_n1117), .B2(KEYINPUT123), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1183), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1188), .B(new_n1101), .C1(new_n1112), .C2(new_n1118), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1163), .B(new_n1181), .C1(new_n1189), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n1193));
  XNOR2_X1  g768(.A(G290), .B(G1986), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n993), .B1(new_n1012), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1192), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1193), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1019), .B1(new_n1196), .B2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n1200));
  NOR3_X1   g774(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1201), .A2(new_n676), .ZN(new_n1202));
  INV_X1    g776(.A(new_n1202), .ZN(new_n1203));
  AND4_X1   g777(.A1(new_n1200), .A2(new_n984), .A3(new_n913), .A4(new_n1203), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n904), .B1(new_n886), .B2(new_n895), .ZN(new_n1205));
  INV_X1    g779(.A(new_n905), .ZN(new_n1206));
  OAI21_X1  g780(.A(KEYINPUT104), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n903), .A2(new_n908), .A3(new_n905), .ZN(new_n1208));
  INV_X1    g782(.A(new_n896), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n1207), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1210), .A2(new_n862), .ZN(new_n1211));
  AOI21_X1  g785(.A(new_n1202), .B1(new_n1211), .B2(new_n907), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1200), .B1(new_n1212), .B2(new_n984), .ZN(new_n1213));
  NOR2_X1   g787(.A1(new_n1204), .A2(new_n1213), .ZN(G308));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n984), .ZN(G225));
endmodule


