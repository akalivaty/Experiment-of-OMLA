//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n455), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n464), .A2(new_n465), .A3(G137), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(G101), .A3(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n468), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n465), .A2(KEYINPUT69), .A3(new_n470), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n479), .A2(new_n464), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n482), .A2(G136), .B1(G124), .B2(new_n483), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n464), .C2(G112), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n476), .B(new_n478), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n488), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(new_n470), .B2(G114), .ZN(new_n494));
  NOR2_X1   g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT70), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT4), .A4(G138), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n493), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT71), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n509), .B(new_n511), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(G543), .B1(new_n517), .B2(new_n518), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n514), .A2(new_n525), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n516), .A2(new_n524), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  OAI21_X1  g103(.A(G89), .B1(new_n517), .B2(new_n518), .ZN(new_n529));
  INV_X1    g104(.A(G63), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n512), .ZN(new_n533));
  INV_X1    g108(.A(new_n521), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(G51), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n519), .A2(new_n541), .B1(new_n521), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n533), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n531), .B2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n519), .A2(new_n548), .B1(new_n521), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT73), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n533), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n531), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND3_X1  g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n534), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(new_n519), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n566), .A2(KEYINPUT75), .A3(G91), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n519), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(KEYINPUT76), .B(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n512), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n567), .A2(new_n570), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n565), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G74), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n531), .B1(new_n512), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(G87), .B2(new_n566), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n534), .A2(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G288));
  OAI211_X1 g155(.A(G48), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n519), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n509), .A2(new_n511), .A3(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n531), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n583), .A2(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n566), .A2(G85), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n534), .A2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n533), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n531), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT77), .B(G66), .Z(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n512), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n534), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT10), .B1(new_n519), .B2(new_n597), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n592), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  OR3_X1    g179(.A1(G168), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT78), .B1(G168), .B2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(G299), .A2(new_n604), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G297));
  NAND3_X1  g183(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n601), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n554), .A2(new_n604), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n600), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n604), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n483), .A2(G123), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT79), .Z(new_n617));
  NAND2_X1  g192(.A1(new_n482), .A2(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n464), .C2(G111), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2096), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT80), .ZN(new_n639));
  OAI21_X1  g214(.A(G14), .B1(new_n636), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2067), .B(G2678), .Z(new_n642));
  XNOR2_X1  g217(.A(G2084), .B(G2090), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(KEYINPUT17), .B2(new_n646), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(new_n643), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n650), .C1(KEYINPUT17), .C2(new_n646), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n645), .B(KEYINPUT81), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n648), .B(new_n651), .C1(new_n650), .C2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2096), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(G227));
  XOR2_X1   g230(.A(G1956), .B(G2474), .Z(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  NOR2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n672), .B(new_n673), .Z(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G1981), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G229));
  NAND2_X1  g252(.A1(G115), .A2(G2104), .ZN(new_n678));
  INV_X1    g253(.A(G127), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n479), .B2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n464), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT93), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n482), .A2(G139), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT25), .Z(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G29), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G29), .B2(G33), .ZN(new_n690));
  INV_X1    g265(.A(G2072), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(G29), .A2(G32), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT26), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n482), .B2(G141), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n483), .A2(G129), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n470), .A2(G105), .A3(G2104), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT96), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n693), .B1(new_n701), .B2(G29), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT27), .B(G1996), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  INV_X1    g279(.A(KEYINPUT98), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G5), .B2(G16), .ZN(new_n706));
  OR3_X1    g281(.A1(new_n705), .A2(G5), .A3(G16), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n706), .B(new_n707), .C1(G301), .C2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT99), .B(G1961), .Z(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(G160), .A2(G29), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  NOR2_X1   g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT94), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(KEYINPUT94), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n713), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT95), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2084), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT91), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G4), .B2(G16), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n723), .A2(G4), .A3(G16), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n724), .B(new_n725), .C1(new_n600), .C2(new_n708), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT92), .B(G1348), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(G299), .A2(G16), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n708), .A2(KEYINPUT23), .A3(G20), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT23), .ZN(new_n731));
  INV_X1    g306(.A(G20), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G16), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n729), .A2(new_n730), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1956), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n712), .A2(new_n722), .A3(new_n728), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n714), .A2(G35), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n714), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT29), .B(G2090), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n714), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n714), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT100), .B(G2078), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n555), .A2(new_n708), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n708), .B2(G19), .ZN(new_n748));
  INV_X1    g323(.A(G1341), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n748), .A2(new_n749), .B1(new_n690), .B2(new_n691), .ZN(new_n750));
  NAND2_X1  g325(.A1(G168), .A2(G16), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G16), .B2(G21), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT31), .B(G11), .Z(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n752), .B2(new_n753), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n620), .A2(G29), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n760), .B(new_n714), .C1(new_n758), .C2(G28), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n754), .A2(new_n756), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  NOR4_X1   g337(.A1(new_n737), .A2(new_n746), .A3(new_n750), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n708), .A2(G23), .ZN(new_n764));
  INV_X1    g339(.A(G288), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n708), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT33), .B(G1976), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT89), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(G6), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G305), .B2(new_n708), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT32), .B(G1981), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n771), .A2(new_n772), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n775), .ZN(new_n778));
  INV_X1    g353(.A(new_n776), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n773), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n769), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G22), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G166), .B2(G16), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT90), .B(G1971), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OR3_X1    g360(.A1(new_n781), .A2(new_n785), .A3(KEYINPUT34), .ZN(new_n786));
  OAI21_X1  g361(.A(KEYINPUT34), .B1(new_n781), .B2(new_n785), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n708), .A2(G24), .ZN(new_n788));
  XNOR2_X1  g363(.A(G290), .B(KEYINPUT85), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n708), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT86), .B(G1986), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n714), .A2(G25), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n482), .A2(G131), .B1(G119), .B2(new_n483), .ZN(new_n794));
  OAI221_X1 g369(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n793), .B1(new_n797), .B2(new_n714), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT35), .B(G1991), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT84), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n786), .A2(new_n787), .A3(new_n792), .A4(new_n801), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(KEYINPUT36), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n692), .B(new_n763), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n714), .A2(G26), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n482), .A2(G140), .B1(G128), .B2(new_n483), .ZN(new_n807));
  OAI221_X1 g382(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n464), .C2(G116), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n806), .B1(new_n810), .B2(new_n714), .ZN(new_n811));
  MUX2_X1   g386(.A(new_n806), .B(new_n811), .S(KEYINPUT28), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G2067), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n748), .A2(new_n749), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n805), .A2(new_n813), .A3(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  INV_X1    g393(.A(G67), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n512), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G651), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT101), .Z(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI22_X1  g399(.A1(new_n519), .A2(new_n823), .B1(new_n521), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT37), .Z(new_n828));
  NOR2_X1   g403(.A1(new_n600), .A2(new_n610), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT39), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n826), .A2(new_n555), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n822), .A2(new_n825), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n554), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n832), .B(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n828), .B1(new_n837), .B2(G860), .ZN(G145));
  XNOR2_X1  g413(.A(new_n809), .B(new_n505), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n688), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n700), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n482), .A2(G142), .B1(G130), .B2(new_n483), .ZN(new_n842));
  OAI221_X1 g417(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n623), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n796), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT104), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT104), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n841), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(G160), .B(KEYINPUT103), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G162), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(new_n620), .Z(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n849), .B(new_n853), .C1(new_n841), .C2(new_n847), .ZN(new_n854));
  INV_X1    g429(.A(G37), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n840), .B(new_n701), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(KEYINPUT105), .A3(new_n846), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n846), .A2(KEYINPUT105), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n841), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n852), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n855), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g437(.A(G299), .B(new_n601), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n836), .A2(KEYINPUT106), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n836), .A2(KEYINPUT106), .ZN(new_n866));
  INV_X1    g441(.A(new_n613), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n836), .A2(KEYINPUT106), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n613), .B1(new_n869), .B2(new_n864), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n863), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n863), .A2(new_n873), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n869), .A2(new_n613), .A3(new_n864), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(KEYINPUT108), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G305), .B(KEYINPUT107), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G303), .ZN(new_n884));
  XNOR2_X1  g459(.A(G288), .B(G290), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(KEYINPUT108), .B2(new_n880), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n871), .B(new_n878), .C1(KEYINPUT108), .C2(new_n880), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n882), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n882), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(G868), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n826), .A2(new_n604), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(G295));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n893), .ZN(G331));
  XNOR2_X1  g470(.A(G301), .B(G286), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n836), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n833), .A2(new_n835), .A3(new_n896), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n863), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n876), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n886), .B(new_n900), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n855), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT111), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n874), .A2(KEYINPUT109), .A3(new_n875), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n901), .B(new_n908), .C1(KEYINPUT109), .C2(new_n874), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n886), .B1(new_n909), .B2(new_n900), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT111), .B1(new_n905), .B2(new_n910), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(KEYINPUT43), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n905), .B1(new_n915), .B2(new_n887), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(KEYINPUT110), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n887), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n906), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n914), .A2(new_n918), .A3(new_n922), .A4(KEYINPUT44), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n906), .A2(new_n917), .A3(new_n911), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(new_n916), .B2(new_n917), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(G397));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n505), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g505(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G125), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n467), .B1(new_n479), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n681), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n936), .A2(G40), .A3(new_n471), .A4(new_n469), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G2067), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n809), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n700), .A2(G1996), .ZN(new_n941));
  INV_X1    g516(.A(G1996), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n796), .A2(new_n799), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n796), .A2(new_n799), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(G290), .A2(G1986), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(G290), .A2(G1986), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n938), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT53), .ZN(new_n952));
  INV_X1    g527(.A(G40), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n468), .A2(new_n472), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n933), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n956), .B2(G2078), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n937), .B1(new_n930), .B2(KEYINPUT50), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT50), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n505), .A2(new_n959), .A3(new_n929), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(G1961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n957), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n505), .A2(new_n929), .A3(new_n931), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n954), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n505), .B2(new_n929), .ZN(new_n967));
  OR4_X1    g542(.A1(new_n952), .A2(new_n966), .A3(G2078), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(G171), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n753), .B1(new_n966), .B2(new_n967), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT120), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n930), .A2(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G2084), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n954), .A4(new_n960), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G8), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n973), .B1(new_n972), .B2(new_n976), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT51), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(G168), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n972), .A2(new_n976), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(G8), .A3(G168), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n985), .A2(KEYINPUT51), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT62), .ZN(new_n987));
  INV_X1    g562(.A(new_n982), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT51), .B(new_n988), .C1(new_n978), .C2(new_n979), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n983), .A2(new_n986), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2090), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n958), .A2(new_n991), .A3(new_n960), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n931), .B1(new_n505), .B2(new_n929), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n993), .A2(new_n994), .A3(new_n937), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n992), .B1(new_n995), .B2(G1971), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G8), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n999), .A3(G8), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1971), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n956), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n981), .B1(new_n1004), .B2(new_n992), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(KEYINPUT113), .A3(new_n999), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT123), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n578), .A2(G1976), .A3(new_n579), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(G160), .A2(new_n505), .A3(G40), .A4(new_n929), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n578), .A2(KEYINPUT114), .A3(G1976), .A4(new_n579), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1011), .A2(new_n1012), .A3(G8), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1015));
  OR3_X1    g590(.A1(new_n583), .A2(new_n586), .A3(G1981), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1981), .B1(new_n583), .B2(new_n586), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1017), .A3(KEYINPUT49), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(G8), .A3(new_n1012), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n765), .B2(G1976), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1015), .B(new_n1022), .C1(new_n1014), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n960), .A2(KEYINPUT116), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n505), .A2(new_n1027), .A3(new_n959), .A4(new_n929), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n958), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1029), .A2(G2090), .B1(new_n995), .B2(G1971), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(G8), .ZN(new_n1031));
  INV_X1    g606(.A(new_n999), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1025), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1007), .A2(new_n1008), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1008), .B1(new_n1007), .B2(new_n1033), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n971), .B(new_n990), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n983), .A2(new_n986), .A3(new_n989), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1039), .A2(new_n1040), .A3(KEYINPUT62), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1039), .B2(KEYINPUT62), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT113), .B1(new_n1005), .B2(new_n999), .ZN(new_n1044));
  AND4_X1   g619(.A1(KEYINPUT113), .A2(new_n996), .A3(G8), .A4(new_n999), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1033), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT123), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1007), .A2(new_n1008), .A3(new_n1033), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(KEYINPUT124), .A3(new_n971), .A4(new_n990), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1038), .A2(new_n1043), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1022), .A2(new_n1052), .A3(new_n765), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1016), .ZN(new_n1054));
  XOR2_X1   g629(.A(new_n1054), .B(KEYINPUT115), .Z(new_n1055));
  NAND2_X1  g630(.A1(new_n1012), .A2(G8), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT63), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1005), .A2(new_n999), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1058), .A2(new_n1025), .A3(new_n985), .ZN(new_n1059));
  OAI22_X1  g634(.A1(new_n1055), .A2(new_n1056), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n999), .B1(new_n1030), .B2(G8), .ZN(new_n1061));
  OR3_X1    g636(.A1(new_n1061), .A2(KEYINPUT63), .A3(new_n985), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1025), .B1(new_n1062), .B2(new_n1007), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(KEYINPUT121), .A2(G2078), .ZN(new_n1065));
  NAND2_X1  g640(.A1(KEYINPUT121), .A2(G2078), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n952), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n995), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1068), .B(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(new_n964), .A3(G301), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT54), .B1(new_n1071), .B2(new_n970), .ZN(new_n1072));
  XOR2_X1   g647(.A(G299), .B(KEYINPUT57), .Z(new_n1073));
  NAND2_X1  g648(.A1(new_n1029), .A2(new_n735), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT56), .B(G2072), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n995), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1073), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1012), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1012), .A2(new_n1079), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n939), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1348), .B1(new_n958), .B2(new_n960), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(KEYINPUT61), .B(new_n1078), .C1(new_n1085), .C2(new_n600), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1077), .B1(new_n1086), .B2(KEYINPUT119), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1078), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1072), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1083), .A2(new_n601), .A3(new_n1084), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1084), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n600), .B1(new_n1092), .B2(new_n1082), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT60), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1085), .A2(new_n1095), .A3(new_n601), .ZN(new_n1096));
  OR3_X1    g671(.A1(new_n956), .A2(KEYINPUT118), .A3(G1996), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1098));
  XOR2_X1   g673(.A(KEYINPUT58), .B(G1341), .Z(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n956), .B2(G1996), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n555), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1102), .B2(new_n555), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1094), .B(new_n1096), .C1(new_n1104), .C2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1077), .B1(new_n1078), .B2(new_n1093), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1090), .A2(new_n1108), .A3(new_n1049), .ZN(new_n1109));
  INV_X1    g684(.A(new_n969), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G301), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1070), .A2(new_n964), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1111), .B(KEYINPUT54), .C1(G301), .C2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n1039), .C1(KEYINPUT61), .C2(new_n1078), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1064), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n951), .B1(new_n1051), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n938), .A2(new_n942), .ZN(new_n1117));
  XOR2_X1   g692(.A(new_n1117), .B(KEYINPUT46), .Z(new_n1118));
  INV_X1    g693(.A(new_n938), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n940), .B2(new_n701), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(new_n1121), .B(KEYINPUT47), .Z(new_n1122));
  INV_X1    g697(.A(new_n946), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n944), .A2(new_n1123), .B1(G2067), .B2(new_n809), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n938), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT126), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n938), .A2(new_n950), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT48), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n947), .B2(new_n1119), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1122), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1116), .A2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g706(.A1(new_n462), .A2(G227), .ZN(new_n1133));
  INV_X1    g707(.A(KEYINPUT127), .ZN(new_n1134));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AND3_X1   g709(.A1(new_n861), .A2(new_n676), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1137));
  NOR2_X1   g711(.A1(new_n1137), .A2(G401), .ZN(new_n1138));
  AND3_X1   g712(.A1(new_n1136), .A2(new_n925), .A3(new_n1138), .ZN(G308));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n925), .A3(new_n1138), .ZN(G225));
endmodule


