//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT69), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT68), .Z(new_n213));
  OAI21_X1  g0013(.A(new_n206), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT70), .Z(new_n215));
  INV_X1    g0015(.A(KEYINPUT1), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n216), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT64), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n206), .B2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G13), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n221), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g0029(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  INV_X1    g0032(.A(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n226), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AND3_X1   g0037(.A1(new_n217), .A2(new_n218), .A3(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  INV_X1    g0047(.A(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT71), .B(G50), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT72), .ZN(new_n253));
  XOR2_X1   g0053(.A(G107), .B(G116), .Z(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT73), .B1(new_n259), .B2(new_n227), .ZN(new_n260));
  INV_X1    g0060(.A(new_n227), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT73), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(new_n258), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n257), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n260), .B2(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n268), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT74), .ZN(new_n273));
  OR2_X1    g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT75), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n279), .B1(new_n276), .B2(new_n278), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G223), .A3(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n284), .B(new_n285), .C1(new_n286), .C2(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n231), .A2(new_n258), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n272), .A2(new_n273), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n274), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n203), .A2(G20), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G150), .ZN(new_n296));
  XNOR2_X1  g0096(.A(KEYINPUT8), .B(G58), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n233), .A2(G33), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n294), .B(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n229), .A2(new_n230), .A3(new_n300), .ZN(new_n301));
  NOR3_X1   g0101(.A1(new_n221), .A2(new_n233), .A3(G1), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n299), .A2(new_n301), .B1(new_n202), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n302), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n233), .A2(G1), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT76), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n306), .A3(G50), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT78), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(KEYINPUT78), .B1(new_n303), .B2(new_n307), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n293), .A2(G190), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  AOI22_X1  g0116(.A1(G200), .A2(new_n292), .B1(new_n312), .B2(KEYINPUT9), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n316), .B1(new_n315), .B2(new_n317), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n293), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n292), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n308), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n297), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n295), .B1(G20), .B2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT15), .B(G87), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n298), .B2(new_n328), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n301), .B1(new_n286), .B2(new_n302), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n304), .A2(new_n306), .A3(G77), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n276), .A2(new_n278), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT75), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT3), .B(G33), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n279), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G107), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n288), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  MUX2_X1   g0140(.A(G232), .B(G238), .S(G1698), .Z(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(G244), .A2(new_n269), .B1(new_n264), .B2(new_n267), .ZN(new_n343));
  AOI21_X1  g0143(.A(G169), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OR3_X1    g0144(.A1(new_n332), .A2(new_n333), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n333), .B1(new_n332), .B2(new_n344), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n342), .A2(new_n343), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n321), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(G190), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n332), .C1(new_n351), .C2(new_n347), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n320), .A2(new_n325), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n306), .A2(new_n326), .ZN(new_n355));
  INV_X1    g0155(.A(new_n304), .ZN(new_n356));
  INV_X1    g0156(.A(new_n302), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n355), .A2(new_n356), .B1(new_n357), .B2(new_n326), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G68), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n248), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G20), .B1(new_n361), .B2(new_n201), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n295), .A2(G159), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n277), .A2(G33), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT7), .B(new_n233), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n233), .B1(new_n280), .B2(new_n281), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n365), .B1(new_n372), .B2(new_n360), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n301), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n368), .A2(KEYINPUT81), .ZN(new_n377));
  AOI21_X1  g0177(.A(G20), .B1(new_n276), .B2(new_n278), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT80), .B1(new_n378), .B2(KEYINPUT7), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT80), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n371), .C1(new_n336), .C2(G20), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT81), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT7), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n377), .A2(new_n379), .A3(new_n381), .A4(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G68), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n364), .A2(new_n374), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n376), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT82), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n375), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(new_n375), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n359), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(KEYINPUT83), .B(new_n359), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n271), .A2(G1698), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(G223), .B2(G1698), .ZN(new_n396));
  INV_X1    g0196(.A(G87), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n396), .A2(new_n334), .B1(new_n275), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n289), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G232), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n268), .C1(new_n270), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G169), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n321), .B2(new_n401), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n393), .A2(new_n394), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT18), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n393), .A2(new_n406), .A3(new_n394), .A4(new_n403), .ZN(new_n407));
  INV_X1    g0207(.A(G190), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(G200), .B2(new_n401), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n359), .B(new_n410), .C1(new_n389), .C2(new_n390), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n385), .A2(new_n386), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n301), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT7), .B1(new_n338), .B2(new_n233), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n416), .B2(new_n369), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT16), .B1(new_n417), .B2(new_n365), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT82), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n375), .A2(new_n387), .A3(new_n388), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n421), .A2(KEYINPUT17), .A3(new_n359), .A4(new_n410), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n405), .A2(new_n407), .A3(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(G238), .A2(new_n269), .B1(new_n264), .B2(new_n267), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT13), .ZN(new_n427));
  NOR2_X1   g0227(.A1(G226), .A2(G1698), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n400), .B2(G1698), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n335), .A2(new_n337), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G97), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n426), .B(new_n427), .C1(new_n432), .C2(new_n288), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n269), .A2(G238), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n268), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n288), .B1(new_n430), .B2(new_n431), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT13), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(G169), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n433), .A2(new_n437), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n439), .A2(KEYINPUT14), .B1(new_n440), .B2(G179), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT79), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n323), .B1(new_n433), .B2(new_n437), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND4_X1   g0245(.A1(new_n442), .A2(new_n438), .A3(new_n444), .A4(G169), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n441), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n233), .A2(G33), .A3(G77), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n295), .A2(G50), .B1(G20), .B2(new_n360), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n376), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n450), .A2(KEYINPUT11), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(KEYINPUT11), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n302), .A2(new_n360), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n453), .B(KEYINPUT12), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n304), .A2(new_n306), .A3(G68), .ZN(new_n455));
  AND4_X1   g0255(.A1(new_n451), .A2(new_n452), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n447), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n440), .A2(new_n351), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n456), .B1(new_n438), .B2(new_n408), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n354), .A2(new_n425), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n335), .A2(new_n337), .A3(G250), .A4(G1698), .ZN(new_n466));
  AND2_X1   g0266(.A1(KEYINPUT4), .A2(G244), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n335), .A2(new_n337), .A3(new_n283), .A4(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n276), .A2(new_n278), .A3(G244), .A4(new_n283), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  AOI22_X1  g0270(.A1(new_n469), .A2(new_n470), .B1(G33), .B2(G283), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT84), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT84), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n466), .A2(new_n468), .A3(new_n474), .A4(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n289), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n265), .A2(G45), .ZN(new_n477));
  OR2_X1    g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n260), .B2(new_n263), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n481), .A2(G257), .B1(new_n264), .B2(new_n480), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT85), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n476), .A2(KEYINPUT85), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(G200), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n339), .A2(KEYINPUT6), .A3(G97), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(new_n339), .ZN(new_n490));
  NOR2_X1   g0290(.A1(G97), .A2(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n488), .B1(new_n492), .B2(KEYINPUT6), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n493), .A2(G20), .B1(G77), .B2(new_n295), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n372), .B2(new_n339), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n301), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n357), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n265), .A2(G33), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n304), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n482), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n475), .A2(new_n289), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(new_n473), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n501), .B1(G190), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n476), .A2(new_n321), .A3(new_n482), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n483), .A2(new_n323), .B1(new_n496), .B2(new_n500), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n487), .A2(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n336), .A2(G244), .A3(G1698), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n336), .A2(G238), .A3(new_n283), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n477), .A2(G274), .ZN(new_n513));
  INV_X1    g0313(.A(G250), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n513), .B1(new_n514), .B2(new_n477), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n260), .A2(new_n263), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n512), .A2(new_n289), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G190), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n351), .B2(new_n517), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n233), .B1(new_n431), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n491), .A2(new_n397), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n276), .A2(new_n278), .A3(new_n233), .A4(G68), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n520), .B1(new_n298), .B2(new_n489), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT86), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n376), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT86), .A4(new_n525), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n328), .A2(new_n302), .ZN(new_n531));
  INV_X1    g0331(.A(new_n499), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n397), .C2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n519), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n328), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n499), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n530), .A2(new_n536), .A3(new_n531), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT87), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n530), .A2(new_n536), .A3(KEYINPUT87), .A4(new_n531), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n517), .A2(G169), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n321), .B2(new_n517), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n534), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n508), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n264), .A2(new_n480), .ZN(new_n546));
  INV_X1    g0346(.A(new_n480), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n516), .A2(new_n547), .A3(G270), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT88), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G264), .A2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n334), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n336), .A2(KEYINPUT88), .A3(G264), .A4(G1698), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n336), .A2(G257), .A3(new_n283), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G303), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n335), .B2(new_n337), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n289), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n323), .B1(new_n550), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n304), .A2(G116), .A3(new_n498), .ZN(new_n561));
  INV_X1    g0361(.A(G116), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n302), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(G20), .B1(G33), .B2(G283), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n275), .A2(G97), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n564), .A2(new_n565), .B1(G20), .B2(new_n562), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n566), .A2(new_n301), .A3(KEYINPUT20), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT20), .B1(new_n566), .B2(new_n301), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n561), .B(new_n563), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n550), .A2(G190), .A3(new_n559), .ZN(new_n573));
  INV_X1    g0373(.A(new_n569), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n556), .A2(new_n558), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n549), .B1(new_n575), .B2(new_n289), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n573), .B(new_n574), .C1(new_n576), .C2(new_n351), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(G179), .A3(new_n569), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n560), .A2(KEYINPUT21), .A3(new_n569), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n572), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n233), .A2(G107), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT23), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(KEYINPUT23), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n583), .A2(new_n584), .B1(G20), .B2(new_n511), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n397), .A2(KEYINPUT22), .A3(G20), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n335), .A2(new_n337), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT89), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n282), .A2(KEYINPUT89), .A3(new_n587), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n336), .A2(new_n233), .A3(G87), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n594));
  OAI211_X1 g0394(.A(KEYINPUT24), .B(new_n586), .C1(new_n592), .C2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT24), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n590), .A2(new_n591), .B1(KEYINPUT22), .B2(new_n593), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(new_n585), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n598), .A3(new_n301), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n221), .A2(G1), .ZN(new_n600));
  OR2_X1    g0400(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n601));
  NAND2_X1  g0401(.A1(KEYINPUT90), .A2(KEYINPUT25), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n581), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n600), .A2(new_n581), .ZN(new_n604));
  OAI221_X1 g0404(.A(new_n603), .B1(new_n602), .B2(new_n604), .C1(new_n532), .C2(new_n339), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n336), .A2(G257), .A3(G1698), .ZN(new_n608));
  NAND2_X1  g0408(.A1(G33), .A2(G294), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n336), .A2(new_n283), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n514), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n289), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n481), .A2(G264), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n546), .A3(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n614), .A2(G179), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n323), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n607), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT91), .B1(new_n614), .B2(G190), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n614), .A2(new_n351), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT91), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n599), .A3(new_n606), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n580), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n465), .A2(new_n545), .A3(new_n625), .ZN(G372));
  INV_X1    g0426(.A(KEYINPUT92), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n579), .A2(new_n578), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT21), .B1(new_n560), .B2(new_n569), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n572), .A2(KEYINPUT92), .A3(new_n578), .A4(new_n579), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n617), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n508), .A3(new_n544), .A4(new_n623), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n541), .A2(new_n543), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(new_n534), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n506), .B(new_n501), .C1(new_n504), .C2(G169), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n544), .A2(KEYINPUT26), .A3(new_n506), .A4(new_n507), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n636), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n464), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n325), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n458), .B1(new_n461), .B2(new_n349), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n424), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n391), .A2(new_n403), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT18), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n391), .A2(new_n406), .A3(new_n403), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n646), .B1(new_n652), .B2(new_n320), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n645), .A2(new_n653), .ZN(G369));
  OR2_X1    g0454(.A1(new_n580), .A2(KEYINPUT93), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n580), .A2(KEYINPUT93), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n600), .A2(new_n233), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n655), .B(new_n656), .C1(new_n574), .C2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n632), .A2(new_n569), .A3(new_n662), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G330), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n607), .A2(KEYINPUT94), .A3(new_n662), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n617), .A2(new_n667), .A3(new_n623), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT94), .B1(new_n607), .B2(new_n662), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n617), .A2(new_n663), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT95), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n617), .A2(new_n662), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n628), .A2(new_n629), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n662), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(new_n675), .A3(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n223), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  NOR4_X1   g0481(.A1(new_n681), .A2(new_n265), .A3(G116), .A4(new_n522), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n682), .B1(new_n236), .B2(new_n681), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  AOI21_X1  g0484(.A(new_n662), .B1(new_n634), .B2(new_n643), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(KEYINPUT29), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n599), .A2(new_n606), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n615), .A2(new_n616), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n676), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n508), .A2(new_n690), .A3(new_n544), .A4(new_n623), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n643), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n663), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n624), .A2(new_n508), .A3(new_n544), .A4(new_n663), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n517), .A2(new_n613), .A3(new_n612), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n576), .A2(new_n698), .A3(G179), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n697), .B1(new_n699), .B2(new_n483), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n550), .A2(new_n559), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(new_n321), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n504), .A2(new_n702), .A3(KEYINPUT30), .A4(new_n698), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n517), .A2(G179), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n483), .A2(new_n614), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n700), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n662), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n710));
  OAI211_X1 g0510(.A(new_n696), .B(new_n709), .C1(new_n707), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n695), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n684), .B1(new_n714), .B2(G1), .ZN(G364));
  NOR2_X1   g0515(.A1(new_n221), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n265), .B1(new_n716), .B2(G45), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n681), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n232), .B1(G20), .B2(new_n323), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n282), .A2(new_n223), .ZN(new_n726));
  INV_X1    g0526(.A(G355), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n726), .A2(new_n727), .B1(G116), .B2(new_n223), .ZN(new_n728));
  INV_X1    g0528(.A(G45), .ZN(new_n729));
  OR2_X1    g0529(.A1(new_n251), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n223), .A2(new_n334), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n729), .B2(new_n236), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n233), .A2(new_n321), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n735), .A2(new_n408), .A3(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n408), .A2(new_n351), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n736), .A2(G322), .B1(new_n739), .B2(G326), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n408), .A2(G179), .A3(G200), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n233), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G294), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n338), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n233), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(new_n408), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G190), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n734), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n748), .A2(G283), .B1(new_n751), .B2(G311), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n737), .A2(new_n746), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n735), .A2(new_n351), .A3(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT33), .B(G317), .Z(new_n756));
  OAI221_X1 g0556(.A(new_n752), .B1(new_n557), .B2(new_n753), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n746), .A2(new_n749), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n745), .B(new_n757), .C1(G329), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n747), .A2(new_n339), .ZN(new_n764));
  INV_X1    g0564(.A(new_n753), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n764), .B(new_n338), .C1(G87), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT99), .Z(new_n767));
  NAND2_X1  g0567(.A1(new_n751), .A2(KEYINPUT97), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n751), .A2(KEYINPUT97), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n286), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n742), .A2(new_n489), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n736), .A2(G58), .B1(new_n739), .B2(G50), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(new_n360), .B2(new_n755), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n767), .A2(new_n772), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n761), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n763), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n720), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n719), .B1(new_n725), .B2(new_n733), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n664), .A2(new_n665), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n723), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT100), .ZN(new_n785));
  INV_X1    g0585(.A(G330), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n719), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(new_n666), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT101), .ZN(G396));
  INV_X1    g0591(.A(KEYINPUT103), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n349), .A2(new_n792), .A3(new_n352), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n332), .A2(new_n663), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(KEYINPUT103), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(new_n794), .B1(new_n349), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n685), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n712), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n798), .B(KEYINPUT104), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n719), .B1(new_n797), .B2(new_n712), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n720), .A2(new_n721), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n788), .B1(new_n802), .B2(new_n286), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n754), .A2(G150), .B1(new_n739), .B2(G137), .ZN(new_n804));
  INV_X1    g0604(.A(G143), .ZN(new_n805));
  INV_X1    g0605(.A(new_n736), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n805), .B2(new_n806), .C1(new_n771), .C2(new_n777), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT34), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n334), .B1(new_n748), .B2(G68), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n809), .B1(new_n202), .B2(new_n753), .C1(new_n248), .C2(new_n742), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G132), .B2(new_n762), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n762), .A2(G311), .B1(G87), .B2(new_n748), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT102), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n736), .A2(G294), .B1(new_n739), .B2(G303), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n339), .B2(new_n753), .C1(new_n815), .C2(new_n755), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n771), .A2(new_n562), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n816), .A2(new_n817), .A3(new_n282), .A4(new_n773), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n808), .A2(new_n811), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n803), .B1(new_n781), .B2(new_n819), .C1(new_n796), .C2(new_n722), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n801), .A2(new_n820), .ZN(G384));
  NOR2_X1   g0621(.A1(new_n716), .A2(new_n265), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT110), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n707), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n706), .A2(KEYINPUT110), .A3(new_n662), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n824), .A2(new_n710), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n696), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n456), .A2(new_n663), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n443), .A2(new_n444), .B1(new_n438), .B2(new_n321), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n438), .A2(new_n444), .A3(G169), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(KEYINPUT79), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n443), .A2(new_n442), .A3(new_n444), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n462), .B(new_n830), .C1(new_n835), .C2(new_n456), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n829), .B1(new_n447), .B2(new_n461), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT106), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT106), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n458), .A2(new_n839), .A3(new_n462), .A4(new_n830), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n838), .A2(new_n796), .A3(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT38), .ZN(new_n843));
  INV_X1    g0643(.A(new_n660), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n393), .A2(new_n394), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g0645(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n846));
  AND2_X1   g0646(.A1(new_n411), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n404), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n385), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n374), .B1(new_n849), .B2(new_n364), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n358), .B1(new_n850), .B2(new_n387), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(KEYINPUT107), .A3(new_n844), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT107), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n851), .B2(new_n660), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n403), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n411), .B1(new_n857), .B2(new_n851), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT37), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AOI221_X4 g0659(.A(new_n843), .B1(new_n848), .B2(new_n859), .C1(new_n425), .C2(new_n856), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n425), .A2(new_n856), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n848), .A2(new_n859), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n828), .B(new_n842), .C1(new_n860), .C2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT40), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n393), .A2(new_n394), .A3(new_n844), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n650), .A2(new_n651), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n866), .B1(new_n867), .B2(new_n423), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n404), .A2(new_n845), .A3(new_n847), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n649), .A2(new_n411), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n846), .B1(new_n870), .B2(new_n845), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n868), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n843), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n824), .A2(new_n710), .A3(new_n825), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n617), .A2(new_n580), .A3(new_n623), .A4(new_n663), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n827), .B1(new_n545), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n879), .A2(new_n841), .A3(new_n865), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n864), .A2(new_n865), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n465), .A2(new_n879), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n786), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT111), .Z(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n458), .A2(new_n662), .ZN(new_n887));
  XNOR2_X1  g0687(.A(KEYINPUT109), .B(KEYINPUT39), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n873), .A2(new_n874), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  INV_X1    g0690(.A(new_n856), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n423), .B1(KEYINPUT18), .B2(new_n404), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n892), .B2(new_n407), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n848), .A2(new_n859), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n843), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n895), .B2(new_n874), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n887), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n874), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n838), .A2(new_n840), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n685), .A2(new_n796), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n349), .A2(new_n662), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n898), .A2(new_n903), .B1(new_n867), .B2(new_n660), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n464), .B1(new_n687), .B2(new_n694), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n653), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n905), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n822), .B1(new_n886), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n886), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n493), .A2(KEYINPUT35), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n234), .B(G116), .C1(new_n493), .C2(KEYINPUT35), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT105), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n913), .B2(new_n912), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT36), .Z(new_n916));
  OAI211_X1 g0716(.A(new_n236), .B(G77), .C1(new_n248), .C2(new_n360), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(G50), .B2(new_n360), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(G1), .A3(new_n221), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n910), .A2(new_n916), .A3(new_n919), .ZN(G367));
  NAND2_X1  g0720(.A1(new_n501), .A2(new_n662), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n508), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n507), .A2(new_n506), .A3(new_n662), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(new_n670), .A3(new_n677), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n487), .A2(new_n505), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n640), .B1(new_n927), .B2(new_n617), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n925), .A2(KEYINPUT42), .B1(new_n663), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n533), .A2(new_n662), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n544), .A2(KEYINPUT112), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n635), .B2(new_n930), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT112), .B1(new_n544), .B2(new_n930), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n926), .A2(new_n929), .B1(KEYINPUT43), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n935), .A2(KEYINPUT43), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n936), .B(new_n937), .Z(new_n938));
  INV_X1    g0738(.A(new_n924), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n674), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n938), .B(new_n940), .Z(new_n941));
  XNOR2_X1  g0741(.A(KEYINPUT113), .B(KEYINPUT41), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n681), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n678), .A2(new_n675), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n939), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT44), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n944), .A2(new_n939), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(new_n674), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n672), .B1(new_n676), .B2(new_n662), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n678), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n666), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n713), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n943), .B1(new_n955), .B2(new_n714), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n941), .B1(new_n956), .B2(new_n718), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n724), .B1(new_n223), .B2(new_n328), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n245), .A2(new_n731), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n719), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n334), .B1(new_n747), .B2(new_n489), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n754), .A2(G294), .B1(new_n739), .B2(G311), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n557), .B2(new_n806), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n961), .B(new_n963), .C1(G107), .C2(new_n743), .ZN(new_n964));
  INV_X1    g0764(.A(G317), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n964), .B1(new_n815), .B2(new_n771), .C1(new_n965), .C2(new_n761), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT114), .B1(new_n753), .B2(new_n562), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT46), .ZN(new_n968));
  INV_X1    g0768(.A(G150), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n806), .A2(new_n969), .B1(new_n753), .B2(new_n248), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n771), .A2(new_n202), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n970), .B(new_n971), .C1(G143), .C2(new_n739), .ZN(new_n972));
  INV_X1    g0772(.A(G137), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n761), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n754), .A2(G159), .B1(G77), .B2(new_n748), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n975), .B(new_n282), .C1(new_n360), .C2(new_n742), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n966), .A2(new_n968), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n960), .B1(new_n978), .B2(new_n720), .ZN(new_n979));
  INV_X1    g0779(.A(new_n723), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n935), .B2(new_n980), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT115), .Z(new_n982));
  NAND2_X1  g0782(.A1(new_n957), .A2(new_n982), .ZN(G387));
  INV_X1    g0783(.A(new_n681), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n954), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n953), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n985), .B1(new_n714), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n672), .A2(new_n723), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n242), .A2(new_n729), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n522), .A2(G116), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n989), .A2(new_n731), .B1(new_n990), .B2(new_n726), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n297), .A2(KEYINPUT50), .A3(G50), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT50), .B1(new_n297), .B2(G50), .ZN(new_n993));
  AOI21_X1  g0793(.A(G45), .B1(G68), .B2(G77), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n992), .A2(new_n990), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n991), .A2(new_n995), .B1(new_n339), .B2(new_n680), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n719), .B1(new_n996), .B2(new_n725), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n754), .A2(G311), .B1(new_n739), .B2(G322), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n965), .B2(new_n806), .C1(new_n771), .C2(new_n557), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT48), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n743), .A2(G283), .B1(new_n765), .B2(G294), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n762), .A2(G326), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n336), .B1(new_n748), .B2(G116), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n755), .A2(new_n297), .B1(new_n753), .B2(new_n286), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n334), .B(new_n1011), .C1(G97), .C2(new_n748), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n743), .A2(new_n535), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n762), .A2(G150), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n806), .A2(new_n202), .B1(new_n750), .B2(new_n360), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G159), .B2(new_n739), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n997), .B1(new_n1018), .B2(new_n720), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n986), .A2(new_n718), .B1(new_n988), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n987), .A2(new_n1020), .ZN(G393));
  AOI21_X1  g0821(.A(new_n984), .B1(new_n950), .B2(new_n954), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n954), .B2(new_n950), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n255), .A2(new_n731), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n724), .B1(new_n489), .B2(new_n223), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n755), .A2(new_n557), .B1(new_n753), .B2(new_n815), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n764), .B(new_n1026), .C1(G294), .C2(new_n751), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n338), .C1(new_n562), .C2(new_n742), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G322), .B2(new_n762), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n736), .A2(G311), .B1(new_n739), .B2(G317), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT52), .Z(new_n1031));
  OAI22_X1  g0831(.A1(new_n771), .A2(new_n297), .B1(new_n202), .B2(new_n755), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT116), .Z(new_n1033));
  OAI22_X1  g0833(.A1(new_n806), .A2(new_n777), .B1(new_n738), .B2(new_n969), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT51), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1034), .A2(new_n1035), .B1(new_n762), .B2(G143), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n1035), .B2(new_n1034), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n742), .A2(new_n286), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n336), .B1(new_n753), .B2(new_n360), .C1(new_n397), .C2(new_n747), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1029), .A2(new_n1031), .B1(new_n1033), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n719), .B1(new_n1024), .B2(new_n1025), .C1(new_n1041), .C2(new_n781), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n939), .B2(new_n723), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n950), .B2(new_n718), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1023), .A2(new_n1044), .ZN(G390));
  INV_X1    g0845(.A(new_n796), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n899), .B1(new_n712), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n879), .A2(new_n786), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n842), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n901), .B1(new_n685), .B2(new_n796), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1048), .A2(new_n796), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n899), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n902), .B1(new_n693), .B2(new_n1046), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n842), .A2(G330), .A3(new_n711), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1053), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n464), .A2(new_n1048), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n906), .A2(new_n653), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(KEYINPUT39), .B1(new_n860), .B2(new_n863), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n873), .A2(new_n874), .A3(new_n888), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n887), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1051), .B2(new_n899), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n838), .A2(new_n840), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1056), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n875), .A2(new_n1071), .A3(new_n1067), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1069), .A2(new_n1058), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1049), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1064), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1062), .B1(new_n1053), .B2(new_n1059), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1069), .A2(new_n1058), .A3(new_n1072), .ZN(new_n1077));
  AND3_X1   g0877(.A1(new_n875), .A2(new_n1071), .A3(new_n1067), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n889), .A2(new_n896), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n1068), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1076), .B(new_n1077), .C1(new_n1080), .C2(new_n1049), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1075), .A2(new_n1081), .A3(new_n681), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n718), .B(new_n1077), .C1(new_n1080), .C2(new_n1049), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT118), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n889), .A2(new_n896), .A3(new_n722), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n788), .B1(new_n802), .B2(new_n297), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G107), .A2(new_n754), .B1(new_n736), .B2(G116), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n815), .B2(new_n738), .C1(new_n771), .C2(new_n489), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G294), .B2(new_n762), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n360), .A2(new_n747), .B1(new_n753), .B2(new_n397), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n1090), .A2(new_n282), .A3(new_n1038), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n282), .B1(new_n202), .B2(new_n747), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n762), .B2(G125), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT117), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n736), .A2(G132), .B1(new_n739), .B2(G128), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT54), .B(G143), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1095), .B1(new_n973), .B2(new_n755), .C1(new_n771), .C2(new_n1096), .ZN(new_n1097));
  OR3_X1    g0897(.A1(new_n753), .A2(KEYINPUT53), .A3(new_n969), .ZN(new_n1098));
  OAI21_X1  g0898(.A(KEYINPUT53), .B1(new_n753), .B2(new_n969), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n777), .C2(new_n742), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1089), .A2(new_n1091), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1086), .B1(new_n1102), .B2(new_n781), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1085), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1083), .A2(new_n1084), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1084), .B1(new_n1083), .B2(new_n1105), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT119), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1073), .A2(new_n1074), .A3(new_n717), .ZN(new_n1110));
  OAI21_X1  g0910(.A(KEYINPUT118), .B1(new_n1110), .B2(new_n1104), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1083), .A2(new_n1105), .A3(new_n1084), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT119), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1082), .B1(new_n1109), .B2(new_n1113), .ZN(G378));
  NOR2_X1   g0914(.A1(new_n312), .A2(new_n660), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n320), .A2(new_n325), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n320), .B2(new_n325), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n881), .A2(G330), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n846), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n649), .A2(new_n411), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n866), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n848), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT38), .B1(new_n1127), .B2(new_n868), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n880), .B1(new_n860), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1070), .A2(new_n796), .A3(new_n828), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n895), .B2(new_n874), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1129), .B(G330), .C1(new_n1131), .C2(KEYINPUT40), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1123), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1122), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT123), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(new_n905), .B2(KEYINPUT122), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT122), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1137), .B(KEYINPUT123), .C1(new_n897), .C2(new_n904), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1132), .B(new_n1121), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1067), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n898), .A2(new_n903), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n867), .A2(new_n660), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT122), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT123), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n905), .A2(KEYINPUT122), .A3(new_n1135), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1140), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1139), .A2(new_n1148), .A3(new_n718), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n736), .A2(G107), .B1(new_n739), .B2(G116), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n336), .A2(G41), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n815), .C2(new_n761), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n742), .A2(new_n360), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n755), .A2(new_n489), .B1(new_n328), .B2(new_n750), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n248), .A2(new_n747), .B1(new_n753), .B2(new_n286), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT58), .Z(new_n1157));
  NAND2_X1  g0957(.A1(new_n754), .A2(G132), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n753), .B2(new_n1096), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n736), .A2(G128), .B1(new_n739), .B2(G125), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n973), .B2(new_n750), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1159), .B(new_n1161), .C1(G150), .C2(new_n743), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n762), .A2(G124), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n748), .C2(G159), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT59), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1166), .C1(new_n1162), .C2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1157), .B1(new_n1164), .B2(new_n1168), .C1(new_n1151), .C2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT120), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n720), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT121), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n788), .B1(new_n802), .B2(new_n202), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n1121), .C2(new_n722), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1149), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1081), .A2(new_n1063), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1177), .A2(new_n1139), .A3(new_n1148), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1140), .A2(new_n897), .A3(new_n904), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1134), .A2(new_n905), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1179), .B1(new_n1081), .B2(new_n1063), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n984), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1176), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n899), .A2(new_n721), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n720), .A2(G68), .A3(new_n721), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n562), .A2(new_n755), .B1(new_n806), .B2(new_n815), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G294), .B2(new_n739), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n339), .B2(new_n771), .C1(new_n557), .C2(new_n761), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G77), .A2(new_n748), .B1(new_n765), .B2(G97), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n338), .A3(new_n1013), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G132), .A2(new_n739), .B1(new_n751), .B2(G150), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n334), .B1(new_n748), .B2(G58), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n202), .C2(new_n742), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n736), .A2(G137), .B1(G159), .B2(new_n765), .ZN(new_n1198));
  INV_X1    g0998(.A(G128), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1198), .B1(new_n755), .B2(new_n1096), .C1(new_n1199), .C2(new_n761), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n1192), .A2(new_n1194), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n788), .B(new_n1189), .C1(new_n1201), .C2(new_n720), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1060), .A2(new_n718), .B1(new_n1188), .B2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n943), .B(KEYINPUT124), .ZN(new_n1204));
  OR2_X1    g1004(.A1(new_n1076), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1059), .A2(new_n1053), .A3(new_n1062), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1203), .B1(new_n1205), .B2(new_n1207), .ZN(G381));
  NOR3_X1   g1008(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1111), .A2(new_n1082), .A3(new_n1112), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT125), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1186), .A3(new_n1210), .A4(new_n1212), .ZN(G407));
  NAND2_X1  g1013(.A1(new_n661), .A2(G213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1186), .A2(new_n1210), .A3(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G407), .A2(G213), .A3(new_n1216), .ZN(G409));
  AOI21_X1  g1017(.A(G387), .B1(new_n1023), .B2(new_n1044), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(G393), .B(G396), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G390), .B1(new_n957), .B2(new_n982), .ZN(new_n1220));
  OR3_X1    g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1186), .A2(G378), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1183), .A2(new_n718), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n1175), .C1(new_n1178), .C2(new_n1204), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1210), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1215), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1064), .A2(KEYINPUT60), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1206), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1053), .A2(new_n1059), .A3(new_n1062), .A4(KEYINPUT60), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n681), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G384), .B1(new_n1235), .B2(new_n1203), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1207), .B1(KEYINPUT60), .B2(new_n1064), .ZN(new_n1237));
  OAI211_X1 g1037(.A(G384), .B(new_n1203), .C1(new_n1237), .C2(new_n1233), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1236), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1229), .A2(KEYINPUT63), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1242), .A2(new_n1214), .A3(new_n1240), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1214), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1233), .B1(new_n1230), .B2(new_n1206), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1203), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT126), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1250), .A2(new_n1238), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1215), .A2(G2897), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT126), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(KEYINPUT126), .B(new_n1254), .C1(new_n1236), .C2(new_n1239), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT61), .B1(new_n1246), .B2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1224), .A2(new_n1241), .A3(new_n1245), .A4(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1229), .B2(new_n1259), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT62), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1243), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1229), .A2(KEYINPUT62), .A3(new_n1240), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1264), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT127), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1223), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT62), .B1(new_n1229), .B2(new_n1240), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1261), .B(new_n1269), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1262), .B1(new_n1270), .B2(new_n1274), .ZN(G405));
  INV_X1    g1075(.A(new_n1210), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1225), .B1(new_n1186), .B2(new_n1276), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1277), .B(new_n1240), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(new_n1223), .ZN(G402));
endmodule


