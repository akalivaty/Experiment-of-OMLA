//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936;
  XOR2_X1   g000(.A(KEYINPUT94), .B(G36gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT95), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT14), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT93), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n207), .A2(KEYINPUT93), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n215), .B(KEYINPUT96), .Z(new_n216));
  NOR2_X1   g015(.A1(new_n213), .A2(new_n207), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n205), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT17), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n222), .B1(new_n225), .B2(KEYINPUT97), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n214), .A2(KEYINPUT17), .A3(new_n218), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n221), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n230), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n219), .B(new_n230), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n234), .B(KEYINPUT13), .Z(new_n239));
  AOI22_X1  g038(.A1(new_n236), .A2(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n233), .A2(new_n235), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n234), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G141gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(G197gat), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT11), .B(G169gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(new_n246), .B(KEYINPUT12), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n240), .A2(new_n242), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT98), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT98), .A4(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n248), .B1(new_n240), .B2(new_n242), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G15gat), .B(G43gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(G71gat), .B(G99gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  INV_X1    g060(.A(G176gat), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT23), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n263), .B1(G169gat), .B2(G176gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n266), .B(new_n269), .C1(G183gat), .C2(G190gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND4_X1   g074(.A1(new_n264), .A2(new_n270), .A3(new_n272), .A4(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n273), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT66), .B(G183gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n265), .B(new_n269), .C1(new_n279), .C2(G190gat), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n277), .A2(KEYINPUT67), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT67), .B1(new_n277), .B2(new_n280), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n276), .A2(KEYINPUT25), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .A4(KEYINPUT27), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  AOI21_X1  g091(.A(G190gat), .B1(new_n292), .B2(G183gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n290), .B1(new_n278), .B2(KEYINPUT27), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n285), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n287), .A2(new_n289), .A3(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT68), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n299), .A2(KEYINPUT69), .A3(new_n293), .A4(new_n291), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT27), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n293), .A2(KEYINPUT28), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  OR3_X1    g104(.A1(new_n305), .A2(new_n271), .A3(KEYINPUT70), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT70), .B1(new_n305), .B2(new_n271), .ZN(new_n307));
  INV_X1    g106(.A(new_n271), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n306), .B(new_n307), .C1(KEYINPUT26), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n267), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n284), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  AOI211_X1 g111(.A(KEYINPUT71), .B(new_n310), .C1(new_n301), .C2(new_n303), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n283), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(G113gat), .B(G120gat), .Z(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT72), .B1(new_n320), .B2(new_n321), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n314), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G227gat), .ZN(new_n329));
  INV_X1    g128(.A(G233gat), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n326), .B(new_n283), .C1(new_n312), .C2(new_n313), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n260), .B1(new_n333), .B2(KEYINPUT32), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT33), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n335), .B1(new_n333), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT74), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n337), .A4(new_n334), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n260), .A2(new_n336), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n333), .A2(KEYINPUT32), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n332), .ZN(new_n349));
  INV_X1    g148(.A(new_n331), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT34), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n348), .A2(KEYINPUT75), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n346), .B1(new_n340), .B2(new_n343), .ZN(new_n355));
  INV_X1    g154(.A(new_n352), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT36), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n355), .B2(new_n356), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n353), .A2(new_n357), .A3(new_n359), .A4(KEYINPUT76), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n352), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT77), .B1(new_n355), .B2(new_n356), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n348), .A2(KEYINPUT77), .A3(new_n352), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(new_n358), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n367), .A2(KEYINPUT78), .A3(new_n358), .A4(new_n368), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n364), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(KEYINPUT79), .B(KEYINPUT29), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G141gat), .B(G148gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(KEYINPUT2), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G155gat), .ZN(new_n379));
  INV_X1    g178(.A(G162gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n377), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n377), .B(new_n381), .C1(new_n376), .C2(KEYINPUT2), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n383), .A2(new_n384), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n375), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G197gat), .B(G204gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT22), .ZN(new_n393));
  INV_X1    g192(.A(G211gat), .ZN(new_n394));
  INV_X1    g193(.A(G218gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n391), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n398), .A2(new_n392), .A3(new_n396), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n403), .B(new_n374), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n385), .B1(new_n405), .B2(new_n387), .ZN(new_n406));
  INV_X1    g205(.A(G228gat), .ZN(new_n407));
  OAI22_X1  g206(.A1(new_n401), .A2(new_n406), .B1(new_n407), .B2(new_n330), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n387), .B1(new_n399), .B2(KEYINPUT29), .ZN(new_n409));
  AOI211_X1 g208(.A(new_n407), .B(new_n330), .C1(new_n409), .C2(new_n389), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n391), .B2(new_n400), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G22gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(G22gat), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n408), .B2(new_n411), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n416), .B1(new_n418), .B2(KEYINPUT85), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n413), .A2(new_n419), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n322), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n385), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n385), .B1(new_n324), .B2(new_n325), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n388), .A2(new_n390), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n424), .B1(KEYINPUT3), .B2(new_n389), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n423), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT39), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(G1gat), .B(G29gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT0), .ZN(new_n437));
  XNOR2_X1  g236(.A(G57gat), .B(G85gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n424), .B(new_n389), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n441), .A2(new_n423), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n433), .A2(new_n434), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT40), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n439), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n430), .A2(new_n431), .B1(G225gat), .B2(G233gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT5), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n423), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n428), .A2(KEYINPUT4), .ZN(new_n452));
  INV_X1    g251(.A(new_n425), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n452), .A2(KEYINPUT82), .B1(new_n426), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n428), .A2(new_n455), .A3(KEYINPUT4), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n451), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT5), .B1(new_n441), .B2(new_n423), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n450), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n446), .A2(KEYINPUT87), .B1(new_n447), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT88), .B1(new_n444), .B2(new_n445), .ZN(new_n461));
  OR4_X1    g260(.A1(KEYINPUT88), .A2(new_n440), .A3(new_n443), .A4(new_n445), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n460), .B(new_n463), .C1(KEYINPUT87), .C2(new_n446), .ZN(new_n464));
  NAND2_X1  g263(.A1(G226gat), .A2(G233gat), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n314), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n304), .A2(new_n311), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n283), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT29), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n400), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n468), .A2(new_n465), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n374), .A2(new_n465), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n314), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n399), .ZN(new_n476));
  XNOR2_X1  g275(.A(G8gat), .B(G36gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT80), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT30), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT80), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n472), .A2(new_n483), .A3(new_n476), .A4(new_n479), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT86), .ZN(new_n486));
  INV_X1    g285(.A(new_n479), .ZN(new_n487));
  INV_X1    g286(.A(new_n476), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n399), .B1(new_n466), .B2(new_n470), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n472), .A2(KEYINPUT30), .A3(new_n476), .A4(new_n479), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n486), .B1(new_n485), .B2(new_n492), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n464), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n472), .A2(new_n476), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n487), .B1(new_n497), .B2(KEYINPUT37), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT38), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n471), .A2(new_n399), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT37), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n501), .B1(new_n475), .B2(new_n400), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n499), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT6), .B1(new_n459), .B2(new_n447), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n439), .B(new_n450), .C1(new_n457), .C2(new_n458), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT89), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n452), .A2(KEYINPUT82), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n453), .A2(new_n426), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n456), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n458), .B1(new_n512), .B2(new_n448), .ZN(new_n513));
  INV_X1    g312(.A(new_n450), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n447), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516));
  AND4_X1   g315(.A1(KEYINPUT89), .A2(new_n515), .A3(new_n516), .A4(new_n508), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n447), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT91), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n501), .B1(new_n472), .B2(new_n476), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT38), .B1(new_n498), .B2(new_n522), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n481), .A2(new_n484), .ZN(new_n524));
  AND4_X1   g323(.A1(new_n506), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n422), .B1(new_n496), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n508), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT83), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n507), .A2(KEYINPUT83), .A3(new_n508), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n529), .A2(new_n530), .A3(new_n519), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n413), .B(new_n419), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n485), .A4(new_n492), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n373), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n422), .B1(new_n518), .B2(new_n520), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n485), .A2(new_n492), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT86), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n537), .B1(new_n539), .B2(new_n493), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n355), .A2(new_n356), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n346), .B(new_n352), .C1(new_n340), .C2(new_n343), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT77), .ZN(new_n543));
  INV_X1    g342(.A(new_n368), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n533), .B1(new_n355), .B2(new_n356), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n353), .A2(new_n548), .A3(new_n357), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT92), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n353), .A2(new_n548), .A3(new_n357), .A4(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n531), .A2(new_n538), .A3(new_n546), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n257), .B1(new_n536), .B2(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G57gat), .B(G64gat), .Z(new_n557));
  INV_X1    g356(.A(KEYINPUT99), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  INV_X1    g358(.A(G71gat), .ZN(new_n560));
  INV_X1    g359(.A(G78gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n557), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n558), .B2(new_n562), .ZN(new_n564));
  XNOR2_X1  g363(.A(G71gat), .B(G78gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G127gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n566), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n230), .B1(new_n572), .B2(KEYINPUT21), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n571), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT101), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(G155gat), .ZN(new_n577));
  XOR2_X1   g376(.A(G183gat), .B(G211gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n579), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(KEYINPUT102), .B(G85gat), .Z(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT7), .ZN(new_n587));
  INV_X1    g386(.A(G99gat), .ZN(new_n588));
  INV_X1    g387(.A(G106gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT8), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT103), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g394(.A1(new_n591), .A2(KEYINPUT103), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(KEYINPUT103), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n221), .A2(new_n600), .A3(new_n232), .ZN(new_n601));
  AND2_X1   g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n599), .A2(new_n219), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n572), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n595), .A2(new_n566), .A3(new_n598), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT104), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n616), .A2(new_n622), .A3(new_n617), .A4(new_n618), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n572), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n615), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n616), .A2(new_n618), .ZN(new_n627));
  INV_X1    g426(.A(new_n615), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n626), .A2(new_n629), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n582), .A2(new_n614), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n556), .A2(new_n531), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g439(.A1(new_n494), .A2(new_n495), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n556), .A2(new_n641), .A3(new_n638), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n642), .A2(G8gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G8gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT42), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(KEYINPUT42), .B2(new_n645), .ZN(G1325gat));
  NAND2_X1  g446(.A1(new_n556), .A2(new_n638), .ZN(new_n648));
  OAI21_X1  g447(.A(G15gat), .B1(new_n648), .B2(new_n373), .ZN(new_n649));
  INV_X1    g448(.A(G15gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n367), .A2(new_n368), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n556), .A2(new_n650), .A3(new_n651), .A4(new_n638), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(G1326gat));
  OR3_X1    g452(.A1(new_n648), .A2(KEYINPUT105), .A3(new_n422), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT105), .B1(new_n648), .B2(new_n422), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT43), .B(G22gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  INV_X1    g457(.A(new_n582), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(new_n613), .A3(new_n637), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n556), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n661), .A2(G29gat), .A3(new_n532), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT45), .Z(new_n663));
  AOI21_X1  g462(.A(new_n613), .B1(new_n536), .B2(new_n555), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT108), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n637), .B(KEYINPUT107), .Z(new_n671));
  AOI21_X1  g470(.A(KEYINPUT106), .B1(new_n253), .B2(new_n255), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673));
  AOI211_X1 g472(.A(new_n673), .B(new_n254), .C1(new_n251), .C2(new_n252), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n671), .A2(new_n582), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n670), .A2(new_n531), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(G29gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n678), .ZN(G1328gat));
  INV_X1    g478(.A(new_n641), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n661), .A2(new_n680), .A3(new_n202), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT46), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n670), .A2(new_n641), .A3(new_n676), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n202), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(new_n651), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n661), .A2(G43gat), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n373), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n670), .A2(new_n688), .A3(new_n676), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(G43gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n690), .B(new_n692), .ZN(G1330gat));
  NAND3_X1  g492(.A1(new_n670), .A2(new_n533), .A3(new_n676), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G50gat), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n661), .A2(G50gat), .A3(new_n422), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT48), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(KEYINPUT110), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n695), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n695), .B2(new_n698), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(G1331gat));
  NAND2_X1  g501(.A1(new_n536), .A2(new_n555), .ZN(new_n703));
  NOR4_X1   g502(.A1(new_n671), .A2(new_n675), .A3(new_n582), .A4(new_n614), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n531), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g506(.A1(new_n641), .A2(KEYINPUT111), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n641), .A2(KEYINPUT111), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n711), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n712));
  XOR2_X1   g511(.A(KEYINPUT49), .B(G64gat), .Z(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n711), .B2(new_n713), .ZN(G1333gat));
  AOI21_X1  g513(.A(new_n560), .B1(new_n705), .B2(new_n688), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n686), .A2(G71gat), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n705), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g517(.A1(new_n705), .A2(new_n533), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g519(.A1(new_n659), .A2(new_n675), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n664), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n531), .A2(new_n583), .A3(new_n637), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT112), .Z(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n721), .A2(new_n637), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n670), .A2(new_n531), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n583), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT113), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n727), .B(new_n733), .C1(new_n583), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1336gat));
  INV_X1    g534(.A(new_n710), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(G92gat), .A3(new_n671), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT52), .B1(new_n724), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n669), .B1(new_n703), .B2(new_n614), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n613), .B(new_n666), .C1(new_n536), .C2(new_n555), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n710), .B(new_n729), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G92gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n742), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n738), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n641), .B(new_n729), .C1(new_n739), .C2(new_n740), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G92gat), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n723), .A2(KEYINPUT114), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n664), .A2(new_n721), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n664), .B2(new_n721), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n737), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT115), .B1(new_n754), .B2(KEYINPUT52), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  AOI211_X1 g556(.A(new_n756), .B(new_n757), .C1(new_n748), .C2(new_n753), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n746), .B1(new_n755), .B2(new_n758), .ZN(G1337gat));
  INV_X1    g558(.A(new_n724), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n651), .A2(new_n588), .A3(new_n637), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n670), .A2(new_n688), .A3(new_n729), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n588), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n670), .A2(new_n533), .A3(new_n729), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n751), .A2(new_n752), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n671), .A2(G106gat), .A3(new_n422), .ZN(new_n766));
  AOI22_X1  g565(.A1(G106gat), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n724), .A2(new_n766), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n768), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n764), .A2(G106gat), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n767), .A2(new_n768), .B1(new_n770), .B2(new_n771), .ZN(G1339gat));
  AND2_X1   g571(.A1(new_n623), .A2(new_n624), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n628), .B1(new_n773), .B2(new_n620), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n633), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n628), .A3(new_n620), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n626), .A2(new_n777), .A3(KEYINPUT54), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(KEYINPUT55), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n776), .A2(new_n778), .A3(KEYINPUT117), .A4(KEYINPUT55), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n636), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n781), .A2(KEYINPUT118), .A3(new_n636), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n776), .A2(new_n778), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n785), .A2(new_n675), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n241), .A2(new_n234), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n238), .A2(new_n239), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n246), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n637), .A2(new_n253), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n614), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n614), .A2(new_n253), .A3(new_n793), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n785), .A2(new_n786), .A3(new_n789), .A4(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n582), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n675), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n638), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n533), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n736), .A2(new_n531), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n686), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(G113gat), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n257), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n532), .B1(new_n799), .B2(new_n801), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n550), .A2(new_n552), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n808), .A2(new_n809), .A3(new_n736), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n675), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n807), .B1(new_n811), .B2(new_n806), .ZN(G1340gat));
  INV_X1    g611(.A(G120gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n805), .A2(new_n813), .A3(new_n671), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n637), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n813), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n810), .A2(new_n817), .A3(new_n659), .ZN(new_n818));
  OAI21_X1  g617(.A(G127gat), .B1(new_n805), .B2(new_n582), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n641), .A2(new_n613), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n808), .A2(new_n821), .A3(new_n809), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(KEYINPUT56), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n802), .A2(new_n804), .A3(new_n614), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(G134gat), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT119), .B1(new_n823), .B2(KEYINPUT56), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n823), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT120), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n826), .B(new_n831), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1343gat));
  AOI21_X1  g632(.A(new_n422), .B1(new_n799), .B2(new_n801), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n803), .A2(new_n688), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n256), .A2(new_n789), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n794), .B1(new_n783), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n613), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n659), .B1(new_n840), .B2(new_n797), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n841), .B1(new_n638), .B2(new_n800), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT57), .B1(new_n842), .B2(new_n422), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n836), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G141gat), .B1(new_n844), .B2(new_n257), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n688), .A2(new_n422), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n808), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n710), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n257), .A2(G141gat), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n845), .B(new_n846), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n844), .A2(KEYINPUT121), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n836), .A2(new_n855), .A3(new_n837), .A4(new_n843), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n675), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n853), .B1(new_n857), .B2(G141gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n852), .B1(new_n858), .B2(new_n846), .ZN(G1344gat));
  INV_X1    g658(.A(G148gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n849), .A2(new_n860), .A3(new_n637), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n854), .A2(new_n637), .A3(new_n856), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n860), .A2(KEYINPUT59), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g663(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n840), .A2(new_n797), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n866), .A2(new_n582), .B1(new_n257), .B2(new_n638), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n422), .A2(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n834), .A2(new_n835), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n837), .A2(new_n637), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(KEYINPUT123), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n860), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT123), .B1(new_n870), .B2(new_n871), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n865), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n861), .B1(new_n864), .B2(new_n875), .ZN(G1345gat));
  NAND3_X1  g675(.A1(new_n849), .A2(new_n379), .A3(new_n659), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n854), .A2(new_n659), .A3(new_n856), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n379), .ZN(G1346gat));
  AND3_X1   g678(.A1(new_n854), .A2(new_n614), .A3(new_n856), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n822), .A2(new_n380), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n880), .A2(new_n380), .B1(new_n848), .B2(new_n881), .ZN(G1347gat));
  NOR3_X1   g681(.A1(new_n686), .A2(new_n680), .A3(new_n531), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n802), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n884), .A2(new_n261), .A3(new_n257), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n531), .B1(new_n799), .B2(new_n801), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT124), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n809), .A2(new_n710), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n675), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n885), .B1(new_n889), .B2(new_n261), .ZN(G1348gat));
  OAI21_X1  g689(.A(G176gat), .B1(new_n884), .B2(new_n671), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n637), .A2(new_n262), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(G1349gat));
  OAI21_X1  g693(.A(new_n279), .B1(new_n884), .B2(new_n582), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n292), .A2(G183gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n659), .A2(new_n896), .A3(new_n302), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g698(.A1(new_n613), .A2(G190gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n887), .A2(new_n888), .A3(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT125), .Z(new_n902));
  OAI21_X1  g701(.A(G190gat), .B1(new_n884), .B2(new_n613), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1351gat));
  NAND3_X1  g704(.A1(new_n373), .A2(new_n641), .A3(new_n532), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI221_X1 g706(.A(new_n907), .B1(new_n867), .B2(new_n869), .C1(new_n834), .C2(new_n835), .ZN(new_n908));
  INV_X1    g707(.A(G197gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n257), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n688), .A2(new_n422), .A3(new_n736), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n887), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n675), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n909), .ZN(G1352gat));
  AOI21_X1  g713(.A(G204gat), .B1(new_n635), .B2(new_n636), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n887), .A2(new_n911), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT62), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n887), .A2(new_n918), .A3(new_n911), .A4(new_n915), .ZN(new_n919));
  OAI21_X1  g718(.A(G204gat), .B1(new_n908), .B2(new_n671), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n917), .A2(new_n920), .A3(KEYINPUT126), .A4(new_n919), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n912), .A2(new_n394), .A3(new_n659), .ZN(new_n926));
  OAI21_X1  g725(.A(G211gat), .B1(new_n908), .B2(new_n582), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(G1354gat));
  NAND2_X1  g730(.A1(new_n908), .A2(KEYINPUT127), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(new_n614), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n908), .A2(KEYINPUT127), .ZN(new_n934));
  OAI21_X1  g733(.A(G218gat), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n912), .A2(new_n395), .A3(new_n614), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1355gat));
endmodule


