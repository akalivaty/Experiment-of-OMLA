//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n208), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n213), .A2(KEYINPUT27), .B1(new_n214), .B2(G183gat), .ZN(new_n215));
  AND4_X1   g014(.A1(KEYINPUT68), .A2(new_n214), .A3(KEYINPUT27), .A4(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR3_X1    g016(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT26), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n209), .B(new_n217), .C1(new_n219), .C2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n213), .A2(new_n207), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(KEYINPUT67), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n236));
  AND4_X1   g035(.A1(new_n230), .A2(new_n232), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  INV_X1    g037(.A(G169gat), .ZN(new_n239));
  INV_X1    g038(.A(G176gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(new_n225), .A3(KEYINPUT25), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n228), .B1(new_n237), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n225), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n232), .A2(new_n230), .A3(new_n235), .A4(new_n236), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT69), .A4(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n233), .A2(KEYINPUT64), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT64), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n252), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n229), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n246), .B1(new_n257), .B2(KEYINPUT65), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n259), .A3(new_n256), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT25), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n227), .B1(new_n250), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G113gat), .ZN(new_n264));
  INV_X1    g063(.A(G113gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G120gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT1), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(KEYINPUT72), .A2(G134gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270));
  NOR3_X1   g069(.A1(new_n270), .A2(KEYINPUT1), .A3(G134gat), .ZN(new_n271));
  OAI21_X1  g070(.A(G127gat), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(KEYINPUT72), .B(G134gat), .C1(new_n270), .C2(KEYINPUT1), .ZN(new_n273));
  INV_X1    g072(.A(G134gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n267), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G127gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G227gat), .A2(G233gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n276), .B1(new_n273), .B2(new_n275), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n284), .B(new_n227), .C1(new_n250), .C2(new_n261), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n281), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT33), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n205), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n288), .A2(new_n289), .B1(KEYINPUT32), .B2(new_n286), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n205), .A2(new_n287), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n292), .B1(new_n288), .B2(KEYINPUT73), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n285), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n254), .A2(new_n259), .A3(new_n256), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n259), .B1(new_n254), .B2(new_n256), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n296), .A2(new_n297), .A3(new_n246), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n245), .B(new_n249), .C1(new_n298), .C2(KEYINPUT25), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n284), .B1(new_n299), .B2(new_n227), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n280), .B1(new_n295), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT75), .B1(new_n301), .B2(KEYINPUT34), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(KEYINPUT34), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n285), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .A4(new_n280), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n294), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n308), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n311), .A2(KEYINPUT36), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n303), .A2(new_n307), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n281), .B1(new_n279), .B2(new_n285), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n305), .B1(new_n315), .B2(new_n306), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n288), .A2(new_n289), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n286), .A2(KEYINPUT32), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n288), .A2(KEYINPUT73), .ZN(new_n321));
  INV_X1    g120(.A(new_n292), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n313), .B(new_n308), .C1(new_n290), .C2(new_n293), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT36), .ZN(new_n326));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327));
  XOR2_X1   g126(.A(G155gat), .B(G162gat), .Z(new_n328));
  OR2_X1    g127(.A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(new_n329));
  NAND2_X1  g128(.A1(KEYINPUT80), .A2(KEYINPUT2), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G141gat), .B(G148gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT81), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT81), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n328), .B(new_n335), .C1(new_n332), .C2(new_n331), .ZN(new_n336));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337));
  INV_X1    g136(.A(G155gat), .ZN(new_n338));
  INV_X1    g137(.A(G162gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n340), .B2(KEYINPUT2), .ZN(new_n341));
  INV_X1    g140(.A(G141gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(G148gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT82), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n342), .B2(G148gat), .ZN(new_n346));
  INV_X1    g145(.A(G148gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n344), .B(new_n346), .C1(G141gat), .C2(new_n347), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n334), .A2(new_n336), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT29), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT76), .B(G211gat), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT22), .B1(new_n354), .B2(G218gat), .ZN(new_n355));
  XOR2_X1   g154(.A(G197gat), .B(G204gat), .Z(new_n356));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  OR3_X1    g157(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n355), .B2(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT90), .B1(new_n351), .B2(new_n361), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n341), .ZN(new_n366));
  INV_X1    g165(.A(new_n336), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n347), .A2(G141gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n329), .B(new_n330), .C1(new_n368), .C2(new_n343), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n335), .B1(new_n369), .B2(new_n328), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n367), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT29), .B1(new_n359), .B2(new_n360), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT89), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT89), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n375), .B(new_n371), .C1(new_n372), .C2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n327), .B1(new_n365), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n361), .B(KEYINPUT77), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT91), .B1(new_n379), .B2(new_n351), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n361), .B(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n352), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n373), .A2(G228gat), .A3(G233gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n380), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G78gat), .B(G106gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G22gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT31), .B(G50gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n378), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n378), .B2(new_n386), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT86), .B(KEYINPUT0), .Z(new_n395));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n395), .B(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G57gat), .B(G85gat), .ZN(new_n398));
  XOR2_X1   g197(.A(new_n397), .B(new_n398), .Z(new_n399));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n349), .A2(new_n278), .A3(KEYINPUT84), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT84), .B1(new_n349), .B2(new_n278), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n349), .A2(new_n278), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n407), .B2(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n349), .A2(new_n350), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n272), .A2(KEYINPUT83), .A3(new_n277), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT83), .B1(new_n272), .B2(new_n277), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n403), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n371), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n401), .B2(new_n402), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n405), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n401), .A2(new_n402), .A3(new_n400), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n400), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n418), .A2(new_n405), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n421), .A2(new_n413), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n399), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n425), .A2(KEYINPUT88), .A3(KEYINPUT6), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT88), .B1(new_n425), .B2(KEYINPUT6), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n424), .A3(new_n399), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n419), .A2(new_n424), .ZN(new_n433));
  INV_X1    g232(.A(new_n399), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT87), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n425), .A2(KEYINPUT87), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n432), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440));
  AOI22_X1  g239(.A1(new_n262), .A2(new_n440), .B1(G226gat), .B2(G233gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n299), .B2(new_n227), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(KEYINPUT78), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT78), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n379), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n441), .A2(new_n443), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n361), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT30), .ZN(new_n453));
  XOR2_X1   g252(.A(G64gat), .B(G92gat), .Z(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT79), .ZN(new_n455));
  XNOR2_X1  g254(.A(G8gat), .B(G36gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n452), .A2(new_n453), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n448), .B2(new_n451), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n444), .A2(KEYINPUT78), .ZN(new_n461));
  INV_X1    g260(.A(new_n441), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n447), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n382), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n450), .A3(new_n458), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n460), .A2(new_n465), .A3(KEYINPUT30), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n428), .A2(new_n439), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n312), .B(new_n326), .C1(new_n394), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n413), .A2(new_n422), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n469), .A2(new_n420), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n470), .A2(new_n404), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n434), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT39), .B1(new_n416), .B2(new_n405), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n473), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT40), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n473), .B(KEYINPUT40), .C1(new_n471), .C2(new_n474), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n435), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n466), .A2(new_n459), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n394), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT37), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n452), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n482), .A3(new_n450), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n457), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT38), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT92), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(KEYINPUT38), .C1(new_n483), .C2(new_n485), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n484), .A2(new_n491), .A3(new_n457), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n463), .A2(new_n382), .B1(new_n361), .B2(new_n449), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(KEYINPUT37), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n433), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n425), .A2(KEYINPUT88), .A3(KEYINPUT6), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n497), .B(new_n498), .C1(new_n425), .C2(new_n431), .ZN(new_n499));
  INV_X1    g298(.A(new_n465), .ZN(new_n500));
  NOR3_X1   g299(.A1(new_n494), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n481), .B1(new_n490), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n468), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT94), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT93), .ZN(new_n505));
  AOI211_X1 g304(.A(new_n505), .B(new_n393), .C1(new_n324), .C2(new_n325), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n425), .A2(KEYINPUT87), .ZN(new_n507));
  AOI211_X1 g306(.A(new_n436), .B(new_n399), .C1(new_n419), .C2(new_n424), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n507), .A2(new_n508), .A3(new_n431), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n497), .A2(new_n498), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n480), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n324), .A2(new_n325), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT93), .B1(new_n512), .B2(new_n394), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n506), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n504), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(new_n394), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n505), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n512), .A2(KEYINPUT93), .A3(new_n394), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n467), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n311), .A2(new_n393), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n523), .A2(new_n515), .A3(new_n480), .A4(new_n499), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n503), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G43gat), .B(G50gat), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(KEYINPUT15), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT95), .B(G29gat), .ZN(new_n530));
  INV_X1    g329(.A(G36gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(G29gat), .A2(G36gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(KEYINPUT14), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n534), .A2(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n527), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT97), .B(KEYINPUT17), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n538), .A2(KEYINPUT17), .A3(new_n539), .A4(new_n541), .ZN(new_n545));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT8), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G85gat), .B2(G92gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT103), .ZN(new_n549));
  NAND2_X1  g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n550), .B(new_n551), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XOR2_X1   g352(.A(G99gat), .B(G106gat), .Z(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n554), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n549), .A2(new_n556), .A3(new_n552), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n544), .A2(new_n545), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n542), .A2(new_n560), .B1(KEYINPUT41), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n563), .A2(new_n566), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT101), .ZN(new_n570));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n567), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n567), .B2(new_n568), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n578));
  XOR2_X1   g377(.A(G15gat), .B(G22gat), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT16), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT98), .B1(new_n581), .B2(G1gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n581), .A2(KEYINPUT98), .A3(G1gat), .ZN(new_n584));
  OAI221_X1 g383(.A(new_n578), .B1(G1gat), .B2(new_n580), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(G8gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G71gat), .B(G78gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n587), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n587), .B2(new_n596), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n212), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G211gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n598), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603));
  XOR2_X1   g402(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n577), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n544), .A2(new_n587), .A3(new_n545), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n587), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n612), .A2(new_n613), .B1(new_n615), .B2(new_n542), .ZN(new_n616));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT18), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n587), .B(new_n542), .Z(new_n621));
  XOR2_X1   g420(.A(new_n617), .B(KEYINPUT13), .Z(new_n622));
  AOI22_X1  g421(.A1(new_n618), .A2(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G197gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT11), .B(G169gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT12), .Z(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n620), .A2(new_n623), .A3(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT106), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n592), .B1(new_n557), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n558), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G176gat), .B(G204gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT108), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n558), .A2(new_n645), .A3(new_n592), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT107), .B(KEYINPUT10), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n637), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n638), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n639), .B(new_n644), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT109), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n648), .A2(new_n649), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n639), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n643), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n634), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n525), .A2(new_n611), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n428), .A2(new_n439), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT110), .B(G1gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  INV_X1    g463(.A(new_n480), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n666), .B2(new_n586), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  MUX2_X1   g468(.A(KEYINPUT42), .B(new_n667), .S(new_n669), .Z(G1325gat));
  INV_X1    g469(.A(new_n311), .ZN(new_n671));
  AOI21_X1  g470(.A(G15gat), .B1(new_n659), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n312), .A2(new_n326), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n673), .A2(G15gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n672), .B1(new_n659), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n393), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  NOR2_X1   g477(.A1(new_n525), .A2(new_n658), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n609), .A3(new_n577), .ZN(new_n680));
  INV_X1    g479(.A(new_n530), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n680), .A2(new_n660), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT111), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT45), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n682), .B(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n608), .B(KEYINPUT112), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n658), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n520), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT94), .B1(new_n520), .B2(KEYINPUT35), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n524), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT114), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT114), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n522), .A2(new_n696), .A3(new_n524), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n503), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(KEYINPUT44), .A3(new_n576), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n468), .A2(new_n502), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n576), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT113), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT113), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n704), .B(KEYINPUT44), .C1(new_n525), .C2(new_n576), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n691), .B1(new_n699), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n681), .B1(new_n707), .B2(new_n660), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n684), .A2(new_n688), .A3(new_n708), .ZN(G1328gat));
  NOR3_X1   g508(.A1(new_n680), .A2(G36gat), .A3(new_n480), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT46), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n707), .B2(new_n480), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1329gat));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  INV_X1    g513(.A(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(new_n691), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n703), .A2(new_n705), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n695), .A2(new_n697), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n576), .B1(new_n718), .B2(new_n700), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n702), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n716), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n715), .B1(new_n721), .B2(new_n673), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n671), .A2(new_n715), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n680), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n714), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n673), .ZN(new_n726));
  OAI21_X1  g525(.A(G43gat), .B1(new_n707), .B2(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n727), .B(KEYINPUT47), .C1(new_n680), .C2(new_n723), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n725), .A2(new_n728), .ZN(G1330gat));
  NAND3_X1  g528(.A1(new_n721), .A2(G50gat), .A3(new_n393), .ZN(new_n730));
  INV_X1    g529(.A(G50gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n680), .B2(new_n394), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n730), .A2(KEYINPUT48), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(KEYINPUT48), .B1(new_n730), .B2(new_n732), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(G1331gat));
  NAND3_X1  g534(.A1(new_n634), .A2(new_n610), .A3(new_n656), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n698), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n661), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  INV_X1    g538(.A(new_n737), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n740), .A2(new_n480), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT49), .B(G64gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n737), .A2(new_n665), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT115), .Z(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n740), .B2(new_n311), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n726), .A2(new_n746), .ZN(new_n748));
  AND3_X1   g547(.A1(new_n737), .A2(KEYINPUT116), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT116), .B1(new_n737), .B2(new_n748), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n393), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g553(.A1(new_n633), .A2(new_n608), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT51), .B1(new_n719), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  INV_X1    g556(.A(new_n755), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n698), .A2(new_n757), .A3(new_n576), .A4(new_n758), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n661), .A3(new_n656), .ZN(new_n761));
  INV_X1    g560(.A(G85gat), .ZN(new_n762));
  INV_X1    g561(.A(new_n656), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n717), .B2(new_n720), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n660), .A2(new_n762), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n761), .A2(new_n762), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n665), .B(new_n764), .C1(new_n699), .C2(new_n706), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G92gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n480), .A2(G92gat), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n656), .B(new_n774), .C1(new_n756), .C2(new_n759), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n769), .A2(new_n770), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  AND4_X1   g576(.A1(new_n771), .A2(new_n773), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n772), .B2(G92gat), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n771), .B1(new_n779), .B2(new_n775), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(new_n780), .ZN(G1337gat));
  NOR2_X1   g580(.A1(new_n311), .A2(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n760), .A2(new_n656), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n784), .A3(new_n673), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(G99gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n766), .B2(new_n673), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(G1338gat));
  NOR3_X1   g587(.A1(new_n763), .A2(G106gat), .A3(new_n394), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n760), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n393), .B(new_n764), .C1(new_n699), .C2(new_n706), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(G106gat), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n789), .B(KEYINPUT119), .Z(new_n795));
  AOI22_X1  g594(.A1(new_n760), .A2(new_n795), .B1(new_n793), .B2(G106gat), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n792), .A2(new_n794), .B1(new_n796), .B2(new_n791), .ZN(G1339gat));
  NAND2_X1  g596(.A1(new_n648), .A2(new_n649), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n798), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n648), .A2(KEYINPUT54), .A3(new_n649), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n799), .A2(KEYINPUT55), .A3(new_n643), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n652), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n800), .A2(new_n643), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n803), .B2(new_n799), .ZN(new_n804));
  OR3_X1    g603(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT120), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT120), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n634), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n617), .B1(new_n614), .B2(new_n616), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n621), .A2(new_n622), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n810), .A2(KEYINPUT121), .A3(new_n628), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT121), .B1(new_n810), .B2(new_n628), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n811), .A2(new_n632), .A3(new_n656), .A4(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n576), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n805), .A2(new_n806), .ZN(new_n816));
  AND4_X1   g615(.A1(new_n577), .A2(new_n811), .A3(new_n632), .A4(new_n812), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n689), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n611), .A2(new_n633), .A3(new_n656), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  AOI211_X1 g621(.A(new_n513), .B(new_n506), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n660), .A2(new_n665), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n265), .A3(new_n633), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n820), .A2(new_n822), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n523), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n824), .ZN(new_n830));
  OAI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n634), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n827), .A2(new_n831), .ZN(G1340gat));
  NAND3_X1  g631(.A1(new_n826), .A2(new_n263), .A3(new_n656), .ZN(new_n833));
  OAI21_X1  g632(.A(G120gat), .B1(new_n830), .B2(new_n763), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1341gat));
  XOR2_X1   g634(.A(KEYINPUT72), .B(G127gat), .Z(new_n836));
  NOR3_X1   g635(.A1(new_n830), .A2(new_n689), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n826), .A2(new_n608), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n836), .ZN(G1342gat));
  NAND3_X1  g638(.A1(new_n826), .A2(new_n274), .A3(new_n577), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n830), .B2(new_n576), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n394), .B1(new_n820), .B2(new_n822), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n726), .A2(new_n824), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n633), .A2(new_n342), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n828), .A2(new_n393), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n802), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n799), .A2(new_n643), .A3(new_n800), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(KEYINPUT122), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT55), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n855), .B2(KEYINPUT122), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n854), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n813), .B1(new_n859), .B2(new_n634), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n576), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n608), .B1(new_n861), .B2(new_n818), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n393), .C1(new_n862), .C2(new_n821), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n634), .B(new_n847), .C1(new_n853), .C2(new_n863), .ZN(new_n864));
  OAI221_X1 g663(.A(new_n845), .B1(new_n849), .B2(new_n850), .C1(new_n864), .C2(new_n342), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n847), .B1(new_n853), .B2(new_n863), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n342), .B1(new_n866), .B2(new_n633), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n849), .A2(new_n850), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT58), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n865), .A2(new_n869), .ZN(G1344gat));
  INV_X1    g669(.A(new_n849), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n347), .A3(new_n656), .ZN(new_n872));
  AOI211_X1 g671(.A(KEYINPUT59), .B(new_n347), .C1(new_n866), .C2(new_n656), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n690), .B1(new_n815), .B2(new_n818), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT57), .B(new_n393), .C1(new_n875), .C2(new_n821), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n876), .A2(KEYINPUT123), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n817), .B(new_n854), .C1(KEYINPUT55), .C2(new_n855), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n608), .B1(new_n861), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n393), .B1(new_n879), .B2(new_n821), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n876), .A2(KEYINPUT123), .B1(new_n852), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n656), .A3(new_n848), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n874), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n872), .B1(new_n873), .B2(new_n884), .ZN(G1345gat));
  AOI21_X1  g684(.A(G155gat), .B1(new_n871), .B2(new_n608), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n689), .A2(new_n338), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n866), .B2(new_n887), .ZN(G1346gat));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n339), .A3(new_n577), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n866), .A2(new_n577), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n339), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n661), .A2(new_n480), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n823), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n239), .A3(new_n633), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n829), .A2(new_n892), .ZN(new_n896));
  OAI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n634), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n894), .B2(new_n656), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n896), .A2(new_n240), .A3(new_n763), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(G1349gat));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n902), .A2(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(KEYINPUT60), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n213), .A2(new_n231), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n896), .B2(new_n689), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n823), .A2(new_n608), .A3(new_n206), .A4(new_n892), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n903), .B(new_n904), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  AND4_X1   g707(.A1(new_n902), .A2(new_n906), .A3(KEYINPUT60), .A4(new_n907), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(G1350gat));
  OAI21_X1  g709(.A(G190gat), .B1(new_n896), .B2(new_n576), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT61), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n207), .A3(new_n577), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1351gat));
  INV_X1    g713(.A(G197gat), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n726), .A2(new_n892), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n877), .B2(new_n881), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n917), .B2(new_n633), .ZN(new_n918));
  INV_X1    g717(.A(new_n916), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n846), .A2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(G197gat), .A3(new_n634), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n918), .A2(new_n921), .ZN(G1352gat));
  NOR2_X1   g721(.A1(new_n763), .A2(G204gat), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT125), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT125), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n846), .A2(new_n927), .A3(new_n919), .A4(new_n923), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n882), .A2(new_n656), .A3(new_n919), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G204gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n925), .A2(new_n928), .ZN(new_n932));
  AOI21_X1  g731(.A(KEYINPUT126), .B1(new_n932), .B2(KEYINPUT62), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n934), .B(new_n926), .C1(new_n925), .C2(new_n928), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n929), .B(new_n931), .C1(new_n933), .C2(new_n935), .ZN(G1353gat));
  OR3_X1    g735(.A1(new_n920), .A2(new_n609), .A3(new_n354), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n882), .A2(new_n608), .A3(new_n919), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  OAI21_X1  g740(.A(new_n577), .B1(new_n917), .B2(KEYINPUT127), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n882), .A2(KEYINPUT127), .A3(new_n919), .ZN(new_n943));
  OAI21_X1  g742(.A(G218gat), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OR3_X1    g743(.A1(new_n920), .A2(G218gat), .A3(new_n576), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1355gat));
endmodule


