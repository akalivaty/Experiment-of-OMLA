//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT2), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G155gat), .B(G162gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n202), .A2(new_n207), .A3(new_n205), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT74), .A3(new_n210), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT3), .ZN(new_n216));
  XOR2_X1   g015(.A(G113gat), .B(G120gat), .Z(new_n217));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(KEYINPUT75), .A3(new_n223), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n228), .A3(new_n210), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n216), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n209), .A2(new_n222), .A3(new_n210), .A4(new_n223), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT5), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n232), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n215), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT5), .B1(new_n244), .B2(new_n238), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n228), .B1(new_n213), .B2(new_n214), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n227), .A3(new_n229), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(KEYINPUT4), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n239), .B1(new_n232), .B2(new_n235), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n241), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G1gat), .B(G29gat), .Z(new_n254));
  XNOR2_X1  g053(.A(G57gat), .B(G85gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(KEYINPUT6), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT6), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT5), .ZN(new_n261));
  INV_X1    g060(.A(new_n214), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT74), .B1(new_n209), .B2(new_n210), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n227), .B(new_n226), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n232), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n265), .B2(new_n239), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n231), .A2(new_n249), .A3(new_n250), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n248), .A2(new_n236), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n240), .ZN(new_n269));
  INV_X1    g068(.A(new_n258), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n260), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n253), .A2(new_n258), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n259), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT37), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  OR3_X1    g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT26), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n280), .B1(new_n278), .B2(new_n279), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT66), .B(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT27), .B1(new_n289), .B2(KEYINPUT67), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT27), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G183gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n288), .B(new_n290), .C1(KEYINPUT67), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT27), .B(G183gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n288), .A2(new_n296), .A3(KEYINPUT28), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n287), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n300));
  NAND2_X1  g099(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n305), .A2(KEYINPUT65), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n286), .A2(KEYINPUT24), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n289), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n305), .A2(KEYINPUT65), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n300), .B1(new_n306), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n288), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n310), .B1(new_n315), .B2(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n305), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT25), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n299), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT29), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n320), .A2(new_n321), .B1(G226gat), .B2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n314), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n323), .A2(new_n318), .B1(new_n298), .B2(new_n287), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328));
  INV_X1    g127(.A(G211gat), .ZN(new_n329));
  INV_X1    g128(.A(G218gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G211gat), .B(G218gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n327), .A3(new_n331), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n322), .A2(new_n326), .A3(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n325), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n320), .A2(G226gat), .A3(G233gat), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n337), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n277), .B1(new_n339), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n338), .B1(new_n322), .B2(new_n326), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n337), .A3(new_n341), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT72), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n276), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(new_n345), .A3(new_n276), .ZN(new_n348));
  XOR2_X1   g147(.A(G8gat), .B(G36gat), .Z(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT73), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT38), .B1(new_n347), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n259), .A2(KEYINPUT83), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n344), .A2(new_n345), .A3(new_n352), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n354), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n345), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT38), .B1(new_n360), .B2(KEYINPUT37), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n275), .A2(new_n355), .A3(new_n356), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n228), .B1(new_n338), .B2(KEYINPUT29), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n364), .B1(new_n215), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n229), .A2(new_n321), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n338), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n332), .A2(KEYINPUT78), .A3(new_n334), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n321), .B(new_n373), .C1(new_n337), .C2(KEYINPUT78), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n374), .A2(new_n228), .B1(new_n209), .B2(new_n210), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n337), .B1(new_n229), .B2(new_n321), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n364), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G22gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n372), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n372), .B2(new_n377), .ZN(new_n381));
  OAI21_X1  g180(.A(G78gat), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n372), .A2(new_n377), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G22gat), .ZN(new_n384));
  INV_X1    g183(.A(G78gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n379), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT31), .B(G50gat), .ZN(new_n387));
  INV_X1    g186(.A(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n382), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n382), .B2(new_n386), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n363), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT39), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n244), .B2(new_n238), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n395), .B1(new_n238), .B2(new_n268), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n394), .B(new_n239), .C1(new_n248), .C2(new_n236), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n397), .A2(KEYINPUT80), .A3(new_n270), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT80), .B1(new_n397), .B2(new_n270), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT40), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(KEYINPUT81), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT81), .B1(new_n400), .B2(new_n401), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n253), .A2(new_n258), .ZN(new_n406));
  OAI211_X1 g205(.A(KEYINPUT40), .B(new_n396), .C1(new_n398), .C2(new_n399), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT30), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n357), .B(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n352), .B1(new_n343), .B2(new_n346), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n406), .B(new_n407), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n405), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(new_n402), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(new_n406), .ZN(new_n416));
  INV_X1    g215(.A(new_n410), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n357), .B(KEYINPUT30), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n393), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n392), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n409), .A2(new_n410), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n273), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n319), .A2(new_n314), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n298), .A2(new_n286), .A3(new_n285), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n224), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G227gat), .ZN(new_n429));
  INV_X1    g228(.A(G233gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n224), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n299), .B(new_n433), .C1(new_n314), .C2(new_n319), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT71), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT34), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(new_n434), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n431), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT32), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(G15gat), .B(G43gat), .Z(new_n443));
  XNOR2_X1  g242(.A(new_n443), .B(KEYINPUT69), .ZN(new_n444));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT70), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n448), .B2(new_n446), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n439), .A2(KEYINPUT32), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n437), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n432), .B1(new_n428), .B2(new_n434), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT32), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n446), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n453), .A2(KEYINPUT33), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n451), .B(new_n437), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n436), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT34), .ZN(new_n461));
  INV_X1    g260(.A(new_n436), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n457), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(KEYINPUT36), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT36), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n461), .A2(new_n462), .A3(new_n457), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n462), .B1(new_n461), .B2(new_n457), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n425), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n392), .B1(new_n466), .B2(new_n467), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT35), .B1(new_n471), .B2(new_n424), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n417), .A2(new_n418), .ZN(new_n473));
  NOR4_X1   g272(.A1(new_n473), .A2(KEYINPUT35), .A3(new_n390), .A4(new_n391), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n275), .A2(new_n356), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT84), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n466), .A2(new_n467), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT84), .B1(new_n459), .B2(new_n463), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n474), .B(new_n475), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n421), .A2(new_n470), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n482));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n484));
  INV_X1    g283(.A(G29gat), .ZN(new_n485));
  INV_X1    g284(.A(G36gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G29gat), .A2(G36gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT85), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT85), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(G29gat), .A3(G36gat), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n483), .A2(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(G43gat), .A2(G50gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(G43gat), .A2(G50gat), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT15), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G43gat), .ZN(new_n497));
  INV_X1    g296(.A(G50gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n493), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n496), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n483), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n489), .A2(new_n491), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n496), .A2(new_n503), .A3(new_n504), .A4(new_n501), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT86), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n496), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n482), .B(new_n502), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n503), .A2(new_n504), .ZN(new_n511));
  INV_X1    g310(.A(new_n496), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(new_n506), .A3(new_n505), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n514), .A2(new_n515), .A3(new_n482), .A4(new_n502), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(G1gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT16), .ZN(new_n519));
  INV_X1    g318(.A(G15gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G22gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n378), .A2(G15gat), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(G1gat), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g323(.A(G8gat), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n526));
  INV_X1    g325(.A(G8gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n526), .B(new_n527), .C1(G1gat), .C2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n525), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n502), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT89), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT18), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n514), .A2(new_n502), .A3(new_n530), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT90), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n514), .A2(new_n530), .A3(new_n539), .A4(new_n502), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n533), .A2(KEYINPUT91), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n540), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n531), .A2(new_n525), .A3(new_n529), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n535), .B(KEYINPUT13), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT91), .B1(new_n533), .B2(new_n541), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n481), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n533), .A2(new_n543), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(new_n535), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n541), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n557), .A2(KEYINPUT92), .A3(new_n547), .A4(new_n542), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n550), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G197gat), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT11), .B(G169gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n563), .B(KEYINPUT12), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT93), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n559), .A2(KEYINPUT93), .A3(new_n564), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n548), .A2(new_n549), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n564), .B1(new_n552), .B2(new_n553), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n567), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n480), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(G71gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n385), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G57gat), .B(G64gat), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT95), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n576), .A2(new_n574), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(KEYINPUT94), .ZN(new_n583));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n577), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n582), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT97), .ZN(new_n596));
  XOR2_X1   g395(.A(G99gat), .B(G106gat), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT97), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n595), .B(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n597), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n588), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n597), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n596), .A2(new_n598), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n581), .A2(new_n587), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n603), .A2(KEYINPUT99), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n604), .A2(new_n605), .A3(new_n606), .A4(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(KEYINPUT10), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT10), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n573), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n608), .A2(new_n610), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(G230gat), .A3(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n573), .B(KEYINPUT100), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n611), .B2(new_n613), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(new_n616), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n620), .B1(new_n624), .B2(new_n619), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT101), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n627), .B(new_n620), .C1(new_n624), .C2(new_n619), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(new_n203), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n588), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(G127gat), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n530), .B1(new_n606), .B2(KEYINPUT21), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n634), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n644), .A3(new_n633), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n604), .A2(new_n605), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n517), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(KEYINPUT41), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n653), .B(new_n655), .C1(new_n531), .C2(new_n652), .ZN(new_n656));
  XNOR2_X1  g455(.A(G134gat), .B(G162gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G190gat), .B(G218gat), .Z(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT98), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n654), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n629), .A2(new_n650), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n572), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n273), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT102), .B(G1gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1324gat));
  INV_X1    g472(.A(new_n670), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n473), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT105), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  OR4_X1    g477(.A1(KEYINPUT105), .A2(new_n670), .A3(new_n423), .A4(new_n677), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OR3_X1    g479(.A1(new_n670), .A2(KEYINPUT103), .A3(new_n423), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT103), .B1(new_n670), .B2(new_n423), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(G8gat), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n676), .B(KEYINPUT104), .Z(new_n684));
  AOI21_X1  g483(.A(new_n684), .B1(new_n681), .B2(new_n682), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n680), .B(new_n683), .C1(KEYINPUT42), .C2(new_n685), .ZN(G1325gat));
  NOR2_X1   g485(.A1(new_n477), .A2(new_n478), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n520), .B1(new_n670), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n468), .A2(new_n464), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n690), .A2(KEYINPUT106), .A3(new_n520), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT106), .B1(new_n690), .B2(new_n520), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n670), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT107), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n572), .A2(new_n422), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n668), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT43), .B(G22gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n629), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n700), .A2(new_n650), .A3(new_n667), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n572), .A2(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(G29gat), .A3(new_n273), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT45), .Z(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT35), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n475), .A2(new_n706), .A3(new_n423), .A4(new_n392), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n472), .B1(new_n687), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n363), .A2(new_n392), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n412), .B1(new_n405), .B2(new_n411), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n415), .A2(KEYINPUT82), .A3(new_n419), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n712), .B2(new_n469), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n705), .B1(new_n713), .B2(new_n666), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n666), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n705), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n421), .A2(new_n470), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n708), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n570), .A2(new_n569), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n559), .A2(KEYINPUT93), .A3(new_n564), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT93), .B1(new_n559), .B2(new_n564), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT108), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n700), .A2(new_n650), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n720), .A2(new_n273), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n704), .B1(new_n485), .B2(new_n731), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n702), .A2(G36gat), .A3(new_n423), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n720), .A2(new_n423), .A3(new_n730), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n486), .B2(new_n735), .ZN(G1329gat));
  NOR3_X1   g535(.A1(new_n702), .A2(G43gat), .A3(new_n687), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n480), .B2(new_n667), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n713), .A2(new_n705), .A3(new_n716), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n740), .A2(new_n689), .A3(new_n728), .A4(new_n729), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n737), .B1(new_n741), .B2(G43gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g542(.A(new_n696), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n498), .A3(new_n701), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n720), .A2(new_n392), .A3(new_n730), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(new_n498), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1331gat));
  NAND2_X1  g548(.A1(new_n726), .A2(new_n727), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n750), .A2(new_n650), .A3(new_n667), .A4(new_n700), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n480), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n273), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n756));
  INV_X1    g555(.A(G64gat), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n752), .B(new_n473), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT110), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1333gat));
  NOR4_X1   g560(.A1(new_n480), .A2(new_n751), .A3(new_n575), .A4(new_n690), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT111), .ZN(new_n763));
  INV_X1    g562(.A(new_n687), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n752), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n575), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n422), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT112), .B(G78gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1335gat));
  NAND3_X1  g570(.A1(new_n700), .A2(new_n592), .A3(new_n753), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT114), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n713), .A2(new_n666), .ZN(new_n775));
  INV_X1    g574(.A(new_n650), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n750), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n667), .B1(new_n718), .B2(new_n708), .ZN(new_n779));
  INV_X1    g578(.A(new_n777), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(KEYINPUT51), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n773), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n777), .A2(new_n629), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n740), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n273), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1336gat));
  OAI21_X1  g588(.A(G92gat), .B1(new_n787), .B2(new_n423), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n629), .A2(new_n423), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n782), .A2(new_n593), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(KEYINPUT115), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n790), .A2(KEYINPUT115), .A3(new_n795), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1337gat));
  NAND2_X1  g596(.A1(new_n764), .A2(new_n700), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(G99gat), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n783), .B2(new_n784), .ZN(new_n800));
  OAI21_X1  g599(.A(G99gat), .B1(new_n787), .B2(new_n690), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1338gat));
  INV_X1    g601(.A(new_n786), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n738), .B2(new_n739), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n388), .B1(new_n804), .B2(new_n422), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT53), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n422), .B(new_n786), .C1(new_n714), .C2(new_n719), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n700), .A2(new_n388), .A3(new_n422), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT116), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT51), .B1(new_n779), .B2(new_n780), .ZN(new_n812));
  NOR4_X1   g611(.A1(new_n480), .A2(new_n774), .A3(new_n667), .A4(new_n777), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n809), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n809), .B2(new_n814), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n807), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n811), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n778), .B2(new_n781), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT118), .B1(new_n805), .B2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n809), .B2(KEYINPUT117), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n809), .A2(new_n814), .A3(new_n815), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n818), .A2(new_n825), .ZN(G1339gat));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n827), .B(new_n622), .C1(new_n611), .C2(new_n613), .ZN(new_n828));
  INV_X1    g627(.A(new_n619), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n613), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n621), .B(new_n831), .C1(new_n615), .C2(KEYINPUT10), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n614), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT55), .B1(new_n830), .B2(new_n833), .ZN(new_n835));
  INV_X1    g634(.A(new_n620), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n726), .A2(new_n727), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT119), .B1(new_n551), .B2(new_n535), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(new_n545), .B2(new_n546), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n551), .A2(KEYINPUT119), .A3(new_n535), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n563), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(new_n721), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n626), .A2(new_n628), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n716), .B1(new_n838), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n716), .A2(new_n837), .A3(new_n843), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n776), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n728), .A2(new_n668), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n422), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n473), .A2(new_n273), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n764), .ZN(new_n853));
  INV_X1    g652(.A(G113gat), .ZN(new_n854));
  NOR3_X1   g653(.A1(new_n853), .A2(new_n854), .A3(new_n571), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n273), .B1(new_n847), .B2(new_n849), .ZN(new_n856));
  INV_X1    g655(.A(new_n471), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n423), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n728), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n855), .A2(new_n861), .ZN(G1340gat));
  AOI21_X1  g661(.A(G120gat), .B1(new_n860), .B2(new_n700), .ZN(new_n863));
  INV_X1    g662(.A(G120gat), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n798), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n852), .B2(new_n865), .ZN(G1341gat));
  AOI21_X1  g665(.A(KEYINPUT121), .B1(new_n860), .B2(new_n650), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n856), .A2(KEYINPUT121), .A3(new_n650), .A4(new_n859), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n639), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n776), .A2(new_n639), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n850), .A2(new_n764), .A3(new_n851), .A4(new_n871), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT120), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n870), .A2(new_n873), .ZN(G1342gat));
  OAI21_X1  g673(.A(G134gat), .B1(new_n853), .B2(new_n667), .ZN(new_n875));
  INV_X1    g674(.A(G134gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n876), .A3(new_n666), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n860), .A2(new_n879), .A3(new_n876), .A4(new_n666), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n878), .A3(new_n880), .ZN(G1343gat));
  AOI21_X1  g680(.A(new_n392), .B1(new_n847), .B2(new_n849), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n690), .A2(new_n851), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n830), .A2(new_n833), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT55), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n833), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n620), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n844), .B1(new_n890), .B2(new_n571), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n667), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n716), .A2(new_n837), .A3(new_n843), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n650), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n422), .B1(new_n894), .B2(new_n848), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n885), .B1(new_n895), .B2(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G141gat), .B1(new_n897), .B2(new_n571), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n690), .A2(new_n422), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n473), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n856), .A2(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n571), .A2(G141gat), .ZN(new_n903));
  AOI21_X1  g702(.A(KEYINPUT58), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n896), .A3(new_n728), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n907), .A2(G141gat), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n906), .B2(new_n908), .ZN(G1344gat));
  NOR2_X1   g708(.A1(new_n629), .A2(G148gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n902), .A2(KEYINPUT122), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912));
  INV_X1    g711(.A(new_n910), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n901), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n847), .A2(new_n849), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n422), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT57), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n837), .A2(KEYINPUT123), .A3(new_n666), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n890), .B2(new_n667), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n920), .A3(new_n843), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n650), .B1(new_n921), .B2(new_n892), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n669), .A2(new_n571), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n883), .B(new_n422), .C1(new_n922), .C2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n885), .A2(new_n629), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n917), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n911), .A2(new_n914), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(G148gat), .B1(new_n897), .B2(new_n629), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n932), .ZN(G1345gat));
  OAI21_X1  g732(.A(G155gat), .B1(new_n897), .B2(new_n776), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n902), .A2(new_n203), .A3(new_n650), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1346gat));
  AOI21_X1  g735(.A(G162gat), .B1(new_n902), .B2(new_n666), .ZN(new_n937));
  INV_X1    g736(.A(new_n897), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n716), .A2(G162gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n423), .A2(new_n753), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n687), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n850), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(G169gat), .B1(new_n944), .B2(new_n571), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n915), .A2(new_n273), .A3(new_n857), .ZN(new_n947));
  NOR4_X1   g746(.A1(new_n947), .A2(G169gat), .A3(new_n423), .A4(new_n750), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT124), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n947), .A2(new_n423), .ZN(new_n950));
  INV_X1    g749(.A(G169gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(new_n728), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n953), .A3(new_n945), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n949), .A2(new_n954), .ZN(G1348gat));
  OAI21_X1  g754(.A(G176gat), .B1(new_n944), .B2(new_n629), .ZN(new_n956));
  INV_X1    g755(.A(G176gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n791), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n947), .B2(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n944), .B2(new_n776), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n650), .A2(new_n296), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n947), .A2(new_n423), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT60), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(new_n963), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT60), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n966), .A3(new_n960), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n964), .A2(new_n967), .ZN(G1350gat));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n288), .A3(new_n716), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n850), .A2(new_n666), .A3(new_n943), .ZN(new_n970));
  NOR2_X1   g769(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n311), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n971), .B1(new_n970), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(G1351gat));
  NOR2_X1   g774(.A1(new_n899), .A2(new_n423), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n915), .A2(new_n273), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n977), .A2(new_n750), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n689), .A2(new_n942), .ZN(new_n979));
  OAI211_X1 g778(.A(new_n925), .B(new_n979), .C1(new_n882), .C2(new_n883), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n724), .A2(G197gat), .ZN(new_n981));
  OAI22_X1  g780(.A1(new_n978), .A2(G197gat), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(G1352gat));
  NOR3_X1   g782(.A1(new_n977), .A2(G204gat), .A3(new_n629), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  OAI21_X1  g786(.A(G204gat), .B1(new_n980), .B2(new_n629), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(G1353gat));
  INV_X1    g788(.A(new_n977), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n990), .A2(new_n329), .A3(new_n650), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT63), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n917), .A2(new_n650), .A3(new_n925), .A4(new_n979), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n329), .B1(KEYINPUT126), .B2(new_n992), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g795(.A(new_n995), .B(new_n993), .C1(new_n980), .C2(new_n776), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n991), .B1(new_n996), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n980), .B2(new_n667), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n990), .A2(new_n330), .A3(new_n716), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(G1355gat));
endmodule


