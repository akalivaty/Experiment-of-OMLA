

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n1049, n517, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U551 ( .A1(n795), .A2(n794), .ZN(n541) );
  AND2_X2 U552 ( .A1(n536), .A2(n537), .ZN(n535) );
  NAND2_X2 U553 ( .A1(n755), .A2(G8), .ZN(n756) );
  NOR2_X2 U554 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U555 ( .A1(n1028), .A2(n1024), .ZN(n712) );
  OR2_X1 U556 ( .A1(n555), .A2(n554), .ZN(n556) );
  AND2_X1 U557 ( .A1(n788), .A2(n791), .ZN(n543) );
  XNOR2_X1 U558 ( .A(n527), .B(KEYINPUT28), .ZN(n526) );
  NOR2_X1 U559 ( .A1(n706), .A2(n707), .ZN(n723) );
  AND2_X1 U560 ( .A1(n525), .A2(n712), .ZN(n713) );
  BUF_X1 U561 ( .A(n1049), .Z(G164) );
  XNOR2_X1 U562 ( .A(n556), .B(KEYINPUT85), .ZN(n1049) );
  XNOR2_X1 U563 ( .A(n756), .B(KEYINPUT32), .ZN(n517) );
  XNOR2_X1 U564 ( .A(n548), .B(KEYINPUT66), .ZN(n519) );
  XNOR2_X1 U565 ( .A(n548), .B(KEYINPUT66), .ZN(n520) );
  XNOR2_X1 U566 ( .A(n756), .B(KEYINPUT32), .ZN(n784) );
  XNOR2_X1 U567 ( .A(n548), .B(KEYINPUT66), .ZN(n632) );
  AND2_X1 U568 ( .A1(n547), .A2(G2105), .ZN(n548) );
  NAND2_X1 U569 ( .A1(n736), .A2(G1341), .ZN(n525) );
  AND2_X2 U570 ( .A1(n587), .A2(n532), .ZN(G160) );
  NOR2_X2 U571 ( .A1(n1049), .A2(G1384), .ZN(n805) );
  INV_X1 U572 ( .A(KEYINPUT64), .ZN(n524) );
  INV_X1 U573 ( .A(n806), .ZN(n703) );
  INV_X1 U574 ( .A(KEYINPUT100), .ZN(n540) );
  NAND2_X1 U575 ( .A1(G160), .A2(G40), .ZN(n806) );
  NOR2_X1 U576 ( .A1(n543), .A2(n793), .ZN(n794) );
  INV_X1 U577 ( .A(KEYINPUT89), .ZN(n734) );
  NAND2_X1 U578 ( .A1(n736), .A2(G8), .ZN(n747) );
  AND2_X1 U579 ( .A1(n826), .A2(n540), .ZN(n539) );
  NOR2_X1 U580 ( .A1(n538), .A2(n523), .ZN(n537) );
  NOR2_X1 U581 ( .A1(n826), .A2(n540), .ZN(n538) );
  NOR2_X1 U582 ( .A1(n588), .A2(n521), .ZN(n532) );
  INV_X1 U583 ( .A(KEYINPUT23), .ZN(n585) );
  AND2_X1 U584 ( .A1(G125), .A2(n519), .ZN(n521) );
  XOR2_X1 U585 ( .A(n781), .B(n780), .Z(n522) );
  AND2_X1 U586 ( .A1(n1034), .A2(n839), .ZN(n523) );
  XNOR2_X2 U587 ( .A(n704), .B(n524), .ZN(n708) );
  NAND2_X1 U588 ( .A1(n714), .A2(n525), .ZN(n710) );
  NAND2_X1 U589 ( .A1(n528), .A2(n526), .ZN(n725) );
  OR2_X1 U590 ( .A1(n723), .A2(n722), .ZN(n527) );
  NAND2_X1 U591 ( .A1(n529), .A2(n721), .ZN(n528) );
  NAND2_X1 U592 ( .A1(n531), .A2(n530), .ZN(n529) );
  OR2_X1 U593 ( .A1(n711), .A2(n912), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n720), .B(n719), .ZN(n531) );
  NAND2_X1 U595 ( .A1(n535), .A2(n533), .ZN(n842) );
  NAND2_X1 U596 ( .A1(n534), .A2(KEYINPUT100), .ZN(n533) );
  INV_X1 U597 ( .A(n541), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n541), .A2(n539), .ZN(n536) );
  NAND2_X1 U599 ( .A1(n542), .A2(G101), .ZN(n586) );
  XNOR2_X2 U600 ( .A(n546), .B(n545), .ZN(n542) );
  NAND2_X1 U601 ( .A1(n542), .A2(G102), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n542), .A2(G103), .ZN(n897) );
  NAND2_X1 U603 ( .A1(n542), .A2(G105), .ZN(n810) );
  NAND2_X1 U604 ( .A1(n542), .A2(G95), .ZN(n820) );
  NAND2_X1 U605 ( .A1(n542), .A2(G99), .ZN(n629) );
  NAND2_X1 U606 ( .A1(n542), .A2(G100), .ZN(n876) );
  NAND2_X1 U607 ( .A1(n542), .A2(G104), .ZN(n796) );
  NAND2_X1 U608 ( .A1(n542), .A2(G106), .ZN(n884) );
  BUF_X1 U609 ( .A(n736), .Z(n749) );
  NOR2_X2 U610 ( .A1(n547), .A2(G2105), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT14), .B(n596), .Z(n544) );
  INV_X1 U612 ( .A(KEYINPUT91), .ZN(n719) );
  OR2_X2 U613 ( .A1(n759), .A2(n738), .ZN(n739) );
  INV_X1 U614 ( .A(KEYINPUT29), .ZN(n724) );
  XNOR2_X1 U615 ( .A(n735), .B(n734), .ZN(n759) );
  INV_X1 U616 ( .A(KEYINPUT98), .ZN(n780) );
  BUF_X1 U617 ( .A(n747), .Z(n791) );
  INV_X1 U618 ( .A(n832), .ZN(n824) );
  NOR2_X1 U619 ( .A1(n825), .A2(n824), .ZN(n826) );
  INV_X1 U620 ( .A(KEYINPUT67), .ZN(n545) );
  NOR2_X1 U621 ( .A1(G651), .A2(G543), .ZN(n665) );
  XNOR2_X1 U622 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X2 U623 ( .A(G2104), .B(KEYINPUT65), .ZN(n547) );
  NAND2_X1 U624 ( .A1(G126), .A2(n632), .ZN(n549) );
  NAND2_X1 U625 ( .A1(n550), .A2(n549), .ZN(n555) );
  AND2_X1 U626 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U627 ( .A1(n891), .A2(G114), .ZN(n553) );
  NOR2_X1 U628 ( .A1(G2105), .A2(G2104), .ZN(n551) );
  XOR2_X1 U629 ( .A(KEYINPUT17), .B(n551), .Z(n634) );
  NAND2_X1 U630 ( .A1(n634), .A2(G138), .ZN(n552) );
  NAND2_X1 U631 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U632 ( .A1(G89), .A2(n665), .ZN(n557) );
  XNOR2_X1 U633 ( .A(n557), .B(KEYINPUT74), .ZN(n558) );
  XNOR2_X1 U634 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  XOR2_X1 U635 ( .A(G543), .B(KEYINPUT0), .Z(n653) );
  INV_X1 U636 ( .A(G651), .ZN(n562) );
  NOR2_X2 U637 ( .A1(n653), .A2(n562), .ZN(n668) );
  NAND2_X1 U638 ( .A1(G76), .A2(n668), .ZN(n559) );
  NAND2_X1 U639 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U640 ( .A(n561), .B(KEYINPUT5), .ZN(n568) );
  NOR2_X1 U641 ( .A1(G543), .A2(n562), .ZN(n563) );
  XOR2_X2 U642 ( .A(KEYINPUT1), .B(n563), .Z(n664) );
  NAND2_X1 U643 ( .A1(G63), .A2(n664), .ZN(n565) );
  NOR2_X2 U644 ( .A1(G651), .A2(n653), .ZN(n672) );
  NAND2_X1 U645 ( .A1(G51), .A2(n672), .ZN(n564) );
  NAND2_X1 U646 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U647 ( .A(KEYINPUT6), .B(n566), .Z(n567) );
  NAND2_X1 U648 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U649 ( .A(n569), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G72), .A2(n668), .ZN(n571) );
  NAND2_X1 U652 ( .A1(G85), .A2(n665), .ZN(n570) );
  NAND2_X1 U653 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U654 ( .A1(G60), .A2(n664), .ZN(n573) );
  NAND2_X1 U655 ( .A1(G47), .A2(n672), .ZN(n572) );
  NAND2_X1 U656 ( .A1(n573), .A2(n572), .ZN(n574) );
  OR2_X1 U657 ( .A1(n575), .A2(n574), .ZN(G290) );
  AND2_X1 U658 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U659 ( .A(G57), .ZN(G237) );
  NAND2_X1 U660 ( .A1(G77), .A2(n668), .ZN(n577) );
  NAND2_X1 U661 ( .A1(G90), .A2(n665), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U663 ( .A(KEYINPUT9), .B(n578), .ZN(n582) );
  NAND2_X1 U664 ( .A1(G64), .A2(n664), .ZN(n580) );
  NAND2_X1 U665 ( .A1(G52), .A2(n672), .ZN(n579) );
  AND2_X1 U666 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n582), .A2(n581), .ZN(G301) );
  NAND2_X1 U668 ( .A1(G137), .A2(n634), .ZN(n584) );
  NAND2_X1 U669 ( .A1(G113), .A2(n891), .ZN(n583) );
  NAND2_X1 U670 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U671 ( .A1(G7), .A2(G661), .ZN(n589) );
  XNOR2_X1 U672 ( .A(n589), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U673 ( .A(G223), .ZN(n845) );
  NAND2_X1 U674 ( .A1(n845), .A2(G567), .ZN(n590) );
  XOR2_X1 U675 ( .A(KEYINPUT11), .B(n590), .Z(G234) );
  XOR2_X1 U676 ( .A(G860), .B(KEYINPUT72), .Z(n622) );
  NAND2_X1 U677 ( .A1(n668), .A2(G68), .ZN(n591) );
  XNOR2_X1 U678 ( .A(n591), .B(KEYINPUT71), .ZN(n594) );
  NAND2_X1 U679 ( .A1(n665), .A2(G81), .ZN(n592) );
  XOR2_X1 U680 ( .A(KEYINPUT12), .B(n592), .Z(n593) );
  NOR2_X1 U681 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U682 ( .A(n595), .B(KEYINPUT13), .ZN(n597) );
  NAND2_X1 U683 ( .A1(G56), .A2(n664), .ZN(n596) );
  NOR2_X1 U684 ( .A1(n597), .A2(n544), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n672), .A2(G43), .ZN(n598) );
  NAND2_X1 U686 ( .A1(n599), .A2(n598), .ZN(n1024) );
  OR2_X1 U687 ( .A1(n622), .A2(n1024), .ZN(G153) );
  NAND2_X1 U688 ( .A1(G868), .A2(G301), .ZN(n609) );
  NAND2_X1 U689 ( .A1(G92), .A2(n665), .ZN(n606) );
  NAND2_X1 U690 ( .A1(G66), .A2(n664), .ZN(n601) );
  NAND2_X1 U691 ( .A1(G79), .A2(n668), .ZN(n600) );
  NAND2_X1 U692 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U693 ( .A1(G54), .A2(n672), .ZN(n602) );
  XNOR2_X1 U694 ( .A(KEYINPUT73), .B(n602), .ZN(n603) );
  NOR2_X1 U695 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U696 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X2 U697 ( .A(n607), .B(KEYINPUT15), .ZN(n912) );
  INV_X1 U698 ( .A(n912), .ZN(n1028) );
  INV_X1 U699 ( .A(G868), .ZN(n683) );
  NAND2_X1 U700 ( .A1(n1028), .A2(n683), .ZN(n608) );
  NAND2_X1 U701 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U702 ( .A1(G91), .A2(n665), .ZN(n610) );
  XNOR2_X1 U703 ( .A(n610), .B(KEYINPUT68), .ZN(n617) );
  NAND2_X1 U704 ( .A1(G65), .A2(n664), .ZN(n612) );
  NAND2_X1 U705 ( .A1(G78), .A2(n668), .ZN(n611) );
  NAND2_X1 U706 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U707 ( .A1(G53), .A2(n672), .ZN(n613) );
  XNOR2_X1 U708 ( .A(KEYINPUT69), .B(n613), .ZN(n614) );
  NOR2_X1 U709 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U710 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U711 ( .A(KEYINPUT70), .B(n618), .ZN(G299) );
  NOR2_X1 U712 ( .A1(G286), .A2(n683), .ZN(n620) );
  NOR2_X1 U713 ( .A1(G299), .A2(G868), .ZN(n619) );
  NOR2_X1 U714 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U715 ( .A(KEYINPUT75), .B(n621), .Z(G297) );
  NAND2_X1 U716 ( .A1(n622), .A2(G559), .ZN(n623) );
  NAND2_X1 U717 ( .A1(n623), .A2(n912), .ZN(n624) );
  XNOR2_X1 U718 ( .A(n624), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U719 ( .A1(G868), .A2(n1024), .ZN(n627) );
  NAND2_X1 U720 ( .A1(G868), .A2(n912), .ZN(n625) );
  NOR2_X1 U721 ( .A1(G559), .A2(n625), .ZN(n626) );
  NOR2_X1 U722 ( .A1(n627), .A2(n626), .ZN(G282) );
  NAND2_X1 U723 ( .A1(G111), .A2(n891), .ZN(n628) );
  XNOR2_X1 U724 ( .A(n628), .B(KEYINPUT76), .ZN(n631) );
  XOR2_X1 U725 ( .A(KEYINPUT77), .B(n629), .Z(n630) );
  NAND2_X1 U726 ( .A1(n631), .A2(n630), .ZN(n638) );
  NAND2_X1 U727 ( .A1(G123), .A2(n519), .ZN(n633) );
  XNOR2_X1 U728 ( .A(n633), .B(KEYINPUT18), .ZN(n636) );
  BUF_X1 U729 ( .A(n634), .Z(n896) );
  NAND2_X1 U730 ( .A1(G135), .A2(n896), .ZN(n635) );
  NAND2_X1 U731 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U732 ( .A1(n638), .A2(n637), .ZN(n963) );
  XNOR2_X1 U733 ( .A(n963), .B(G2096), .ZN(n639) );
  XNOR2_X1 U734 ( .A(n639), .B(KEYINPUT78), .ZN(n641) );
  INV_X1 U735 ( .A(G2100), .ZN(n640) );
  NAND2_X1 U736 ( .A1(n641), .A2(n640), .ZN(G156) );
  NAND2_X1 U737 ( .A1(G559), .A2(n912), .ZN(n642) );
  XNOR2_X1 U738 ( .A(n1024), .B(n642), .ZN(n681) );
  NOR2_X1 U739 ( .A1(n681), .A2(G860), .ZN(n649) );
  NAND2_X1 U740 ( .A1(G67), .A2(n664), .ZN(n644) );
  NAND2_X1 U741 ( .A1(G80), .A2(n668), .ZN(n643) );
  NAND2_X1 U742 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U743 ( .A1(G93), .A2(n665), .ZN(n646) );
  NAND2_X1 U744 ( .A1(G55), .A2(n672), .ZN(n645) );
  NAND2_X1 U745 ( .A1(n646), .A2(n645), .ZN(n647) );
  OR2_X1 U746 ( .A1(n648), .A2(n647), .ZN(n684) );
  XOR2_X1 U747 ( .A(n649), .B(n684), .Z(G145) );
  NAND2_X1 U748 ( .A1(G49), .A2(n672), .ZN(n651) );
  NAND2_X1 U749 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U750 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U751 ( .A1(n664), .A2(n652), .ZN(n655) );
  NAND2_X1 U752 ( .A1(n653), .A2(G87), .ZN(n654) );
  NAND2_X1 U753 ( .A1(n655), .A2(n654), .ZN(G288) );
  NAND2_X1 U754 ( .A1(G50), .A2(n672), .ZN(n656) );
  XNOR2_X1 U755 ( .A(n656), .B(KEYINPUT80), .ZN(n663) );
  NAND2_X1 U756 ( .A1(G75), .A2(n668), .ZN(n658) );
  NAND2_X1 U757 ( .A1(G88), .A2(n665), .ZN(n657) );
  NAND2_X1 U758 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U759 ( .A1(G62), .A2(n664), .ZN(n659) );
  XNOR2_X1 U760 ( .A(KEYINPUT79), .B(n659), .ZN(n660) );
  NOR2_X1 U761 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U762 ( .A1(n663), .A2(n662), .ZN(G303) );
  NAND2_X1 U763 ( .A1(G61), .A2(n664), .ZN(n667) );
  NAND2_X1 U764 ( .A1(G86), .A2(n665), .ZN(n666) );
  NAND2_X1 U765 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U766 ( .A1(n668), .A2(G73), .ZN(n669) );
  XOR2_X1 U767 ( .A(KEYINPUT2), .B(n669), .Z(n670) );
  NOR2_X1 U768 ( .A1(n671), .A2(n670), .ZN(n674) );
  NAND2_X1 U769 ( .A1(n672), .A2(G48), .ZN(n673) );
  NAND2_X1 U770 ( .A1(n674), .A2(n673), .ZN(G305) );
  XOR2_X1 U771 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n675) );
  XNOR2_X1 U772 ( .A(G288), .B(n675), .ZN(n678) );
  XNOR2_X1 U773 ( .A(G299), .B(G303), .ZN(n676) );
  XNOR2_X1 U774 ( .A(n676), .B(G305), .ZN(n677) );
  XNOR2_X1 U775 ( .A(n678), .B(n677), .ZN(n680) );
  XOR2_X1 U776 ( .A(G290), .B(n684), .Z(n679) );
  XNOR2_X1 U777 ( .A(n680), .B(n679), .ZN(n915) );
  XNOR2_X1 U778 ( .A(n915), .B(n681), .ZN(n682) );
  NOR2_X1 U779 ( .A1(n683), .A2(n682), .ZN(n686) );
  NOR2_X1 U780 ( .A1(G868), .A2(n684), .ZN(n685) );
  NOR2_X1 U781 ( .A1(n686), .A2(n685), .ZN(G295) );
  NAND2_X1 U782 ( .A1(G2084), .A2(G2078), .ZN(n687) );
  XOR2_X1 U783 ( .A(KEYINPUT20), .B(n687), .Z(n688) );
  NAND2_X1 U784 ( .A1(G2090), .A2(n688), .ZN(n689) );
  XNOR2_X1 U785 ( .A(KEYINPUT21), .B(n689), .ZN(n690) );
  NAND2_X1 U786 ( .A1(n690), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U787 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U788 ( .A1(G69), .A2(G120), .ZN(n691) );
  NOR2_X1 U789 ( .A1(G237), .A2(n691), .ZN(n692) );
  NAND2_X1 U790 ( .A1(G108), .A2(n692), .ZN(n851) );
  NAND2_X1 U791 ( .A1(G567), .A2(n851), .ZN(n693) );
  XNOR2_X1 U792 ( .A(KEYINPUT84), .B(n693), .ZN(n700) );
  XOR2_X1 U793 ( .A(KEYINPUT22), .B(KEYINPUT83), .Z(n695) );
  NAND2_X1 U794 ( .A1(G132), .A2(G82), .ZN(n694) );
  XNOR2_X1 U795 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U796 ( .A(n696), .B(KEYINPUT82), .ZN(n697) );
  NOR2_X1 U797 ( .A1(G218), .A2(n697), .ZN(n698) );
  NAND2_X1 U798 ( .A1(G96), .A2(n698), .ZN(n852) );
  NAND2_X1 U799 ( .A1(G2106), .A2(n852), .ZN(n699) );
  NAND2_X1 U800 ( .A1(n700), .A2(n699), .ZN(n871) );
  NAND2_X1 U801 ( .A1(G483), .A2(G661), .ZN(n701) );
  NOR2_X1 U802 ( .A1(n871), .A2(n701), .ZN(n848) );
  NAND2_X1 U803 ( .A1(n848), .A2(G36), .ZN(G176) );
  XOR2_X1 U804 ( .A(G1981), .B(KEYINPUT99), .Z(n702) );
  XNOR2_X1 U805 ( .A(G305), .B(n702), .ZN(n1014) );
  INV_X1 U806 ( .A(n1014), .ZN(n782) );
  NAND2_X1 U807 ( .A1(n805), .A2(n703), .ZN(n704) );
  NAND2_X1 U808 ( .A1(G2072), .A2(n708), .ZN(n705) );
  XNOR2_X1 U809 ( .A(n705), .B(KEYINPUT27), .ZN(n707) );
  INV_X1 U810 ( .A(G1956), .ZN(n1027) );
  NOR2_X1 U811 ( .A1(n708), .A2(n1027), .ZN(n706) );
  INV_X1 U812 ( .A(G299), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n721) );
  INV_X2 U814 ( .A(n708), .ZN(n736) );
  NAND2_X1 U815 ( .A1(n708), .A2(G1996), .ZN(n709) );
  XNOR2_X1 U816 ( .A(n709), .B(KEYINPUT26), .ZN(n714) );
  NOR2_X1 U817 ( .A1(n1024), .A2(n710), .ZN(n711) );
  NAND2_X1 U818 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U819 ( .A1(G2067), .A2(n736), .ZN(n716) );
  NOR2_X1 U820 ( .A1(G1348), .A2(n708), .ZN(n715) );
  NOR2_X1 U821 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U822 ( .A1(n718), .A2(n717), .ZN(n720) );
  XNOR2_X1 U823 ( .A(n725), .B(n724), .ZN(n730) );
  XOR2_X1 U824 ( .A(G2078), .B(KEYINPUT25), .Z(n939) );
  NAND2_X1 U825 ( .A1(n939), .A2(n708), .ZN(n727) );
  NAND2_X1 U826 ( .A1(n749), .A2(G1961), .ZN(n726) );
  NAND2_X1 U827 ( .A1(n727), .A2(n726), .ZN(n732) );
  NOR2_X1 U828 ( .A1(G301), .A2(n732), .ZN(n728) );
  XOR2_X1 U829 ( .A(KEYINPUT90), .B(n728), .Z(n729) );
  NAND2_X1 U830 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U831 ( .A(n731), .B(KEYINPUT92), .ZN(n745) );
  NAND2_X1 U832 ( .A1(G301), .A2(n732), .ZN(n733) );
  XNOR2_X1 U833 ( .A(n733), .B(KEYINPUT93), .ZN(n742) );
  NOR2_X1 U834 ( .A1(G1966), .A2(n747), .ZN(n735) );
  NOR2_X1 U835 ( .A1(n736), .A2(G2084), .ZN(n760) );
  INV_X1 U836 ( .A(n760), .ZN(n737) );
  NAND2_X1 U837 ( .A1(n737), .A2(G8), .ZN(n738) );
  XNOR2_X1 U838 ( .A(KEYINPUT30), .B(n739), .ZN(n740) );
  NOR2_X1 U839 ( .A1(n740), .A2(G168), .ZN(n741) );
  XOR2_X1 U840 ( .A(KEYINPUT31), .B(n743), .Z(n744) );
  NAND2_X1 U841 ( .A1(n745), .A2(n744), .ZN(n757) );
  NAND2_X1 U842 ( .A1(n757), .A2(G286), .ZN(n746) );
  XNOR2_X1 U843 ( .A(n746), .B(KEYINPUT94), .ZN(n754) );
  NOR2_X1 U844 ( .A1(G1971), .A2(n791), .ZN(n748) );
  XOR2_X1 U845 ( .A(KEYINPUT95), .B(n748), .Z(n751) );
  NOR2_X1 U846 ( .A1(n749), .A2(G2090), .ZN(n750) );
  NOR2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U848 ( .A1(n752), .A2(G303), .ZN(n753) );
  NAND2_X1 U849 ( .A1(n754), .A2(n753), .ZN(n755) );
  INV_X1 U850 ( .A(n757), .ZN(n758) );
  NOR2_X1 U851 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U852 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n783) );
  NOR2_X1 U854 ( .A1(G288), .A2(G1976), .ZN(n763) );
  XNOR2_X1 U855 ( .A(n763), .B(KEYINPUT96), .ZN(n773) );
  INV_X1 U856 ( .A(n791), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n773), .A2(n766), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n764), .A2(KEYINPUT33), .ZN(n774) );
  INV_X1 U859 ( .A(n774), .ZN(n769) );
  NAND2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n1016) );
  INV_X1 U861 ( .A(n1016), .ZN(n765) );
  NOR2_X1 U862 ( .A1(KEYINPUT33), .A2(n765), .ZN(n767) );
  AND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U864 ( .A1(n769), .A2(n768), .ZN(n771) );
  AND2_X1 U865 ( .A1(n783), .A2(n771), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n784), .A2(n770), .ZN(n779) );
  INV_X1 U867 ( .A(n771), .ZN(n777) );
  NOR2_X1 U868 ( .A1(G1971), .A2(G303), .ZN(n772) );
  NOR2_X1 U869 ( .A1(n773), .A2(n772), .ZN(n1017) );
  XOR2_X1 U870 ( .A(n1017), .B(KEYINPUT97), .Z(n775) );
  AND2_X1 U871 ( .A1(n775), .A2(n774), .ZN(n776) );
  OR2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n522), .ZN(n795) );
  NAND2_X1 U875 ( .A1(n517), .A2(n783), .ZN(n787) );
  NOR2_X1 U876 ( .A1(G2090), .A2(G303), .ZN(n785) );
  NAND2_X1 U877 ( .A1(G8), .A2(n785), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U879 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U880 ( .A(n789), .B(KEYINPUT88), .Z(n790) );
  XNOR2_X1 U881 ( .A(KEYINPUT24), .B(n790), .ZN(n792) );
  NOR2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U883 ( .A(KEYINPUT37), .B(G2067), .ZN(n827) );
  NAND2_X1 U884 ( .A1(G140), .A2(n896), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U886 ( .A(KEYINPUT34), .B(n798), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n891), .A2(G116), .ZN(n800) );
  NAND2_X1 U888 ( .A1(G128), .A2(n520), .ZN(n799) );
  NAND2_X1 U889 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U890 ( .A(KEYINPUT35), .B(n801), .Z(n802) );
  NOR2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U892 ( .A(KEYINPUT36), .B(n804), .ZN(n908) );
  NOR2_X1 U893 ( .A1(n827), .A2(n908), .ZN(n980) );
  NOR2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U895 ( .A(n807), .B(KEYINPUT86), .ZN(n839) );
  NAND2_X1 U896 ( .A1(n980), .A2(n839), .ZN(n836) );
  INV_X1 U897 ( .A(n836), .ZN(n825) );
  INV_X1 U898 ( .A(G1996), .ZN(n828) );
  NAND2_X1 U899 ( .A1(G141), .A2(n896), .ZN(n809) );
  NAND2_X1 U900 ( .A1(G117), .A2(n891), .ZN(n808) );
  NAND2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n810), .B(KEYINPUT38), .ZN(n812) );
  NAND2_X1 U903 ( .A1(G129), .A2(n520), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n904) );
  OR2_X1 U906 ( .A1(n828), .A2(n904), .ZN(n823) );
  NAND2_X1 U907 ( .A1(n891), .A2(G107), .ZN(n816) );
  NAND2_X1 U908 ( .A1(G119), .A2(n519), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n819) );
  NAND2_X1 U910 ( .A1(G131), .A2(n896), .ZN(n817) );
  XNOR2_X1 U911 ( .A(KEYINPUT87), .B(n817), .ZN(n818) );
  NOR2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n881) );
  NAND2_X1 U914 ( .A1(G1991), .A2(n881), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n967) );
  NAND2_X1 U916 ( .A1(n839), .A2(n967), .ZN(n832) );
  XNOR2_X1 U917 ( .A(G1986), .B(G290), .ZN(n1034) );
  NAND2_X1 U918 ( .A1(n827), .A2(n908), .ZN(n977) );
  NAND2_X1 U919 ( .A1(n904), .A2(n828), .ZN(n958) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n829) );
  XNOR2_X1 U921 ( .A(n829), .B(KEYINPUT101), .ZN(n831) );
  NOR2_X1 U922 ( .A1(G1991), .A2(n881), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT102), .B(n830), .Z(n965) );
  NAND2_X1 U924 ( .A1(n831), .A2(n965), .ZN(n833) );
  NAND2_X1 U925 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n958), .A2(n834), .ZN(n835) );
  XOR2_X1 U927 ( .A(KEYINPUT39), .B(n835), .Z(n837) );
  NAND2_X1 U928 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n977), .A2(n838), .ZN(n840) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U931 ( .A1(n842), .A2(n841), .ZN(n844) );
  XOR2_X1 U932 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n843) );
  XNOR2_X1 U933 ( .A(n844), .B(n843), .ZN(G329) );
  NAND2_X1 U934 ( .A1(n845), .A2(G2106), .ZN(n846) );
  XNOR2_X1 U935 ( .A(n846), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U937 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U939 ( .A1(n849), .A2(n848), .ZN(n850) );
  XOR2_X1 U940 ( .A(KEYINPUT107), .B(n850), .Z(G188) );
  NOR2_X1 U941 ( .A1(n852), .A2(n851), .ZN(G325) );
  XOR2_X1 U942 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U944 ( .A(G132), .ZN(G219) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  INV_X1 U947 ( .A(G82), .ZN(G220) );
  INV_X1 U948 ( .A(G69), .ZN(G235) );
  XOR2_X1 U949 ( .A(G2100), .B(G2096), .Z(n854) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(G2678), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U952 ( .A(KEYINPUT43), .B(G2090), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U956 ( .A(G2084), .B(G2078), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U958 ( .A(G1976), .B(G1956), .Z(n862) );
  XNOR2_X1 U959 ( .A(G1966), .B(G1961), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U961 ( .A(G1971), .B(G1986), .Z(n864) );
  XNOR2_X1 U962 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U964 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U965 ( .A(G2474), .B(KEYINPUT109), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n870) );
  XOR2_X1 U967 ( .A(G1981), .B(KEYINPUT41), .Z(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(G229) );
  INV_X1 U969 ( .A(n871), .ZN(G319) );
  NAND2_X1 U970 ( .A1(n520), .A2(G124), .ZN(n872) );
  XNOR2_X1 U971 ( .A(n872), .B(KEYINPUT44), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT110), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G112), .A2(n891), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G136), .A2(n896), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U977 ( .A1(n879), .A2(n878), .ZN(G162) );
  XOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n880) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(n890) );
  NAND2_X1 U980 ( .A1(n891), .A2(G118), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G130), .A2(n519), .ZN(n882) );
  NAND2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n888) );
  NAND2_X1 U983 ( .A1(G142), .A2(n896), .ZN(n885) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U985 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(n890), .B(n889), .Z(n903) );
  NAND2_X1 U988 ( .A1(n891), .A2(G115), .ZN(n893) );
  NAND2_X1 U989 ( .A1(G127), .A2(n520), .ZN(n892) );
  NAND2_X1 U990 ( .A1(n893), .A2(n892), .ZN(n895) );
  XOR2_X1 U991 ( .A(KEYINPUT112), .B(KEYINPUT47), .Z(n894) );
  XNOR2_X1 U992 ( .A(n895), .B(n894), .ZN(n901) );
  NAND2_X1 U993 ( .A1(G139), .A2(n896), .ZN(n898) );
  NAND2_X1 U994 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U995 ( .A(KEYINPUT111), .B(n899), .Z(n900) );
  NOR2_X1 U996 ( .A1(n901), .A2(n900), .ZN(n970) );
  XNOR2_X1 U997 ( .A(G164), .B(n970), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(n910) );
  XOR2_X1 U999 ( .A(n963), .B(G162), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G160), .B(n904), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n911), .ZN(G395) );
  INV_X1 U1005 ( .A(G301), .ZN(G171) );
  XOR2_X1 U1006 ( .A(KEYINPUT113), .B(G286), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G171), .B(n912), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n917) );
  XOR2_X1 U1009 ( .A(n1024), .B(n915), .Z(n916) );
  XNOR2_X1 U1010 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n918), .ZN(G397) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n920) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n933) );
  XNOR2_X1 U1015 ( .A(G2443), .B(G2427), .ZN(n930) );
  XOR2_X1 U1016 ( .A(G2430), .B(KEYINPUT105), .Z(n922) );
  XNOR2_X1 U1017 ( .A(G2454), .B(G2435), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(n922), .B(n921), .ZN(n926) );
  XOR2_X1 U1019 ( .A(G2438), .B(KEYINPUT104), .Z(n924) );
  XNOR2_X1 U1020 ( .A(G1341), .B(G1348), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n924), .B(n923), .ZN(n925) );
  XOR2_X1 U1022 ( .A(n926), .B(n925), .Z(n928) );
  XNOR2_X1 U1023 ( .A(G2451), .B(G2446), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n928), .B(n927), .ZN(n929) );
  XNOR2_X1 U1025 ( .A(n930), .B(n929), .ZN(n931) );
  NAND2_X1 U1026 ( .A1(n931), .A2(G14), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(G319), .A2(n936), .ZN(n932) );
  NOR2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1029 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  INV_X1 U1032 ( .A(G303), .ZN(G166) );
  INV_X1 U1033 ( .A(G108), .ZN(G238) );
  INV_X1 U1034 ( .A(n936), .ZN(G401) );
  XNOR2_X1 U1035 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n983) );
  XNOR2_X1 U1036 ( .A(G2084), .B(G34), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT54), .ZN(n954) );
  XNOR2_X1 U1038 ( .A(G2090), .B(G35), .ZN(n951) );
  XOR2_X1 U1039 ( .A(G1991), .B(G25), .Z(n938) );
  NAND2_X1 U1040 ( .A1(n938), .A2(G28), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(G1996), .B(G32), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(n939), .B(G27), .ZN(n940) );
  NOR2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(KEYINPUT120), .B(n942), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n949), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(n952), .B(KEYINPUT121), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1054 ( .A(n983), .B(n955), .Z(n957) );
  XNOR2_X1 U1055 ( .A(KEYINPUT122), .B(G29), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n1045) );
  INV_X1 U1057 ( .A(G29), .ZN(n986) );
  XNOR2_X1 U1058 ( .A(KEYINPUT117), .B(KEYINPUT52), .ZN(n982) );
  XNOR2_X1 U1059 ( .A(G2090), .B(G162), .ZN(n959) );
  NAND2_X1 U1060 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1061 ( .A(n960), .B(KEYINPUT51), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G2084), .B(G160), .ZN(n961) );
  XNOR2_X1 U1063 ( .A(KEYINPUT115), .B(n961), .ZN(n962) );
  NOR2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1065 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n976) );
  XOR2_X1 U1068 ( .A(G2072), .B(n970), .Z(n972) );
  XOR2_X1 U1069 ( .A(G164), .B(G2078), .Z(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1071 ( .A(KEYINPUT116), .B(n973), .Z(n974) );
  XNOR2_X1 U1072 ( .A(KEYINPUT50), .B(n974), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n982), .B(n981), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT119), .B(n987), .ZN(n1043) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT59), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n988), .B(G4), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(G1341), .B(G19), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(G6), .B(G1981), .ZN(n989) );
  NOR2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1086 ( .A(G20), .B(G1956), .Z(n993) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n993), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(KEYINPUT60), .B(n996), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1966), .B(G21), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(G5), .B(G1961), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1002) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1003) );
  NAND2_X1 U1098 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1102 ( .A(n1009), .B(KEYINPUT61), .ZN(n1011) );
  INV_X1 U1103 ( .A(G16), .ZN(n1010) );
  NAND2_X1 U1104 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1105 ( .A1(G11), .A2(n1012), .ZN(n1041) );
  XNOR2_X1 U1106 ( .A(G16), .B(KEYINPUT56), .ZN(n1038) );
  XOR2_X1 U1107 ( .A(G168), .B(G1966), .Z(n1013) );
  NOR2_X1 U1108 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1109 ( .A(KEYINPUT57), .B(n1015), .Z(n1023) );
  NAND2_X1 U1110 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  INV_X1 U1111 ( .A(G1971), .ZN(n1018) );
  NOR2_X1 U1112 ( .A1(G166), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1113 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1114 ( .A(KEYINPUT123), .B(n1021), .Z(n1022) );
  NAND2_X1 U1115 ( .A1(n1023), .A2(n1022), .ZN(n1026) );
  XNOR2_X1 U1116 ( .A(G1341), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1117 ( .A1(n1026), .A2(n1025), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(G299), .B(n1027), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(G301), .B(G1961), .ZN(n1030) );
  XNOR2_X1 U1120 ( .A(n1028), .B(G1348), .ZN(n1029) );
  NOR2_X1 U1121 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1122 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1123 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1124 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1125 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1126 ( .A(KEYINPUT124), .B(n1039), .Z(n1040) );
  NOR2_X1 U1127 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  NAND2_X1 U1128 ( .A1(n1043), .A2(n1042), .ZN(n1044) );
  NOR2_X1 U1129 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  XOR2_X1 U1130 ( .A(KEYINPUT127), .B(n1046), .Z(n1047) );
  XNOR2_X1 U1131 ( .A(KEYINPUT62), .B(n1047), .ZN(G311) );
  INV_X1 U1132 ( .A(G311), .ZN(G150) );
endmodule

