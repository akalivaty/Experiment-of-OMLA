

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  INV_X1 U325 ( .A(KEYINPUT32), .ZN(n426) );
  XNOR2_X1 U326 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U327 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n514) );
  XNOR2_X1 U328 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U329 ( .A(n515), .B(n514), .ZN(n548) );
  NOR2_X1 U330 ( .A1(n552), .A2(n551), .ZN(n573) );
  AND2_X1 U331 ( .A1(n558), .A2(n557), .ZN(n568) );
  XOR2_X1 U332 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n454) );
  XNOR2_X1 U333 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n293), .B(KEYINPUT17), .ZN(n294) );
  XOR2_X1 U335 ( .A(n294), .B(KEYINPUT18), .Z(n296) );
  XNOR2_X1 U336 ( .A(G169GAT), .B(G176GAT), .ZN(n295) );
  XOR2_X1 U337 ( .A(n296), .B(n295), .Z(n319) );
  XOR2_X1 U338 ( .A(KEYINPUT89), .B(KEYINPUT65), .Z(n298) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(KEYINPUT90), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U341 ( .A(n319), .B(n299), .Z(n309) );
  XOR2_X1 U342 ( .A(G127GAT), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U343 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n339) );
  XOR2_X1 U345 ( .A(G43GAT), .B(G134GAT), .Z(n383) );
  XOR2_X1 U346 ( .A(n339), .B(n383), .Z(n307) );
  XOR2_X1 U347 ( .A(G113GAT), .B(G15GAT), .Z(n445) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G71GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n302), .B(G120GAT), .ZN(n425) );
  XOR2_X1 U350 ( .A(n425), .B(KEYINPUT20), .Z(n304) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n445), .B(n305), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U355 ( .A(n309), .B(n308), .Z(n557) );
  INV_X1 U356 ( .A(n557), .ZN(n495) );
  XOR2_X1 U357 ( .A(n495), .B(KEYINPUT91), .Z(n362) );
  XOR2_X1 U358 ( .A(G8GAT), .B(KEYINPUT80), .Z(n404) );
  XOR2_X1 U359 ( .A(KEYINPUT98), .B(n404), .Z(n311) );
  NAND2_X1 U360 ( .A1(G226GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n313) );
  XNOR2_X1 U362 ( .A(G36GAT), .B(G190GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n312), .B(KEYINPUT79), .ZN(n379) );
  XOR2_X1 U364 ( .A(n313), .B(n379), .Z(n318) );
  XOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT21), .Z(n315) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n352) );
  XNOR2_X1 U368 ( .A(G204GAT), .B(G92GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n316), .B(G64GAT), .ZN(n422) );
  XNOR2_X1 U370 ( .A(n352), .B(n422), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n321) );
  INV_X1 U372 ( .A(n319), .ZN(n320) );
  XOR2_X1 U373 ( .A(n321), .B(n320), .Z(n492) );
  INV_X1 U374 ( .A(n492), .ZN(n546) );
  XOR2_X1 U375 ( .A(n546), .B(KEYINPUT99), .Z(n322) );
  XNOR2_X1 U376 ( .A(n322), .B(KEYINPUT27), .ZN(n364) );
  XOR2_X1 U377 ( .A(G162GAT), .B(G148GAT), .Z(n324) );
  XNOR2_X1 U378 ( .A(G29GAT), .B(G134GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U380 ( .A(KEYINPUT4), .B(G155GAT), .Z(n326) );
  XNOR2_X1 U381 ( .A(G113GAT), .B(G120GAT), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U383 ( .A(n328), .B(n327), .Z(n333) );
  XOR2_X1 U384 ( .A(KEYINPUT1), .B(KEYINPUT96), .Z(n330) );
  NAND2_X1 U385 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U387 ( .A(G1GAT), .B(n331), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U389 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n335) );
  XNOR2_X1 U390 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U392 ( .A(n337), .B(n336), .Z(n341) );
  XNOR2_X1 U393 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n338), .B(KEYINPUT2), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n339), .B(n343), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n489) );
  XNOR2_X1 U397 ( .A(G85GAT), .B(n489), .ZN(n478) );
  INV_X1 U398 ( .A(n478), .ZN(n552) );
  NAND2_X1 U399 ( .A1(n364), .A2(n552), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n342), .B(KEYINPUT100), .ZN(n516) );
  XOR2_X1 U401 ( .A(G50GAT), .B(G162GAT), .Z(n382) );
  XOR2_X1 U402 ( .A(n382), .B(n343), .Z(n345) );
  NAND2_X1 U403 ( .A1(G228GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n356) );
  XOR2_X1 U405 ( .A(G204GAT), .B(KEYINPUT23), .Z(n347) );
  XNOR2_X1 U406 ( .A(KEYINPUT94), .B(KEYINPUT22), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U408 ( .A(n348), .B(KEYINPUT24), .Z(n350) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U410 ( .A(n401), .B(KEYINPUT92), .ZN(n349) );
  XNOR2_X1 U411 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U412 ( .A(n351), .B(KEYINPUT95), .Z(n354) );
  XNOR2_X1 U413 ( .A(n352), .B(KEYINPUT93), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(G148GAT), .B(G106GAT), .Z(n358) );
  XNOR2_X1 U417 ( .A(KEYINPUT75), .B(G78GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U419 ( .A(KEYINPUT74), .B(n359), .Z(n416) );
  XOR2_X1 U420 ( .A(n360), .B(n416), .Z(n553) );
  XNOR2_X1 U421 ( .A(KEYINPUT28), .B(n553), .ZN(n500) );
  INV_X1 U422 ( .A(n500), .ZN(n519) );
  NOR2_X1 U423 ( .A1(n516), .A2(n519), .ZN(n361) );
  NAND2_X1 U424 ( .A1(n362), .A2(n361), .ZN(n371) );
  NOR2_X1 U425 ( .A1(n553), .A2(n557), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n363), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U427 ( .A1(n572), .A2(n364), .ZN(n368) );
  NAND2_X1 U428 ( .A1(n557), .A2(n546), .ZN(n365) );
  NAND2_X1 U429 ( .A1(n553), .A2(n365), .ZN(n366) );
  XOR2_X1 U430 ( .A(KEYINPUT25), .B(n366), .Z(n367) );
  NAND2_X1 U431 ( .A1(n368), .A2(n367), .ZN(n369) );
  NAND2_X1 U432 ( .A1(n369), .A2(n478), .ZN(n370) );
  NAND2_X1 U433 ( .A1(n371), .A2(n370), .ZN(n463) );
  XOR2_X1 U434 ( .A(KEYINPUT66), .B(KEYINPUT78), .Z(n373) );
  XNOR2_X1 U435 ( .A(G85GAT), .B(KEYINPUT77), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n391) );
  XOR2_X1 U437 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n375) );
  NAND2_X1 U438 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U440 ( .A(n376), .B(KEYINPUT11), .Z(n381) );
  XOR2_X1 U441 ( .A(G29GAT), .B(KEYINPUT7), .Z(n378) );
  XNOR2_X1 U442 ( .A(KEYINPUT70), .B(KEYINPUT8), .ZN(n377) );
  XNOR2_X1 U443 ( .A(n378), .B(n377), .ZN(n442) );
  XNOR2_X1 U444 ( .A(n442), .B(n379), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n387) );
  XOR2_X1 U446 ( .A(n382), .B(G218GAT), .Z(n385) );
  XNOR2_X1 U447 ( .A(n383), .B(G106GAT), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U449 ( .A(n387), .B(n386), .Z(n389) );
  XNOR2_X1 U450 ( .A(G99GAT), .B(G92GAT), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n569) );
  INV_X1 U453 ( .A(n569), .ZN(n543) );
  XOR2_X1 U454 ( .A(G127GAT), .B(G71GAT), .Z(n393) );
  XNOR2_X1 U455 ( .A(G15GAT), .B(G183GAT), .ZN(n392) );
  XNOR2_X1 U456 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U457 ( .A(KEYINPUT14), .B(KEYINPUT81), .Z(n395) );
  XNOR2_X1 U458 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n394) );
  XNOR2_X1 U459 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U460 ( .A(n397), .B(n396), .Z(n403) );
  XOR2_X1 U461 ( .A(KEYINPUT86), .B(KEYINPUT12), .Z(n399) );
  NAND2_X1 U462 ( .A1(G231GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U464 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U465 ( .A(n403), .B(n402), .ZN(n408) );
  XOR2_X1 U466 ( .A(G57GAT), .B(KEYINPUT13), .Z(n421) );
  XOR2_X1 U467 ( .A(n404), .B(n421), .Z(n406) );
  XNOR2_X1 U468 ( .A(G78GAT), .B(G211GAT), .ZN(n405) );
  XNOR2_X1 U469 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U470 ( .A(n408), .B(n407), .Z(n413) );
  XOR2_X1 U471 ( .A(G1GAT), .B(KEYINPUT71), .Z(n440) );
  XOR2_X1 U472 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n410) );
  XNOR2_X1 U473 ( .A(KEYINPUT82), .B(KEYINPUT84), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n440), .B(n411), .ZN(n412) );
  XOR2_X1 U476 ( .A(n413), .B(n412), .Z(n584) );
  INV_X1 U477 ( .A(n584), .ZN(n566) );
  NAND2_X1 U478 ( .A1(n543), .A2(n566), .ZN(n414) );
  XOR2_X1 U479 ( .A(KEYINPUT16), .B(n414), .Z(n415) );
  AND2_X1 U480 ( .A1(n463), .A2(n415), .ZN(n477) );
  INV_X1 U481 ( .A(n416), .ZN(n420) );
  XOR2_X1 U482 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n418) );
  XNOR2_X1 U483 ( .A(G176GAT), .B(G85GAT), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U485 ( .A(n420), .B(n419), .Z(n431) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n424) );
  AND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n425), .B(KEYINPUT33), .ZN(n427) );
  XOR2_X1 U490 ( .A(n431), .B(n430), .Z(n580) );
  XOR2_X1 U491 ( .A(G8GAT), .B(G141GAT), .Z(n433) );
  XNOR2_X1 U492 ( .A(G169GAT), .B(G22GAT), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U494 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n435) );
  XNOR2_X1 U495 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n434) );
  XNOR2_X1 U496 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n450) );
  XOR2_X1 U498 ( .A(G197GAT), .B(G43GAT), .Z(n439) );
  XNOR2_X1 U499 ( .A(G36GAT), .B(G50GAT), .ZN(n438) );
  XNOR2_X1 U500 ( .A(n439), .B(n438), .ZN(n441) );
  XOR2_X1 U501 ( .A(n441), .B(n440), .Z(n448) );
  XOR2_X1 U502 ( .A(n442), .B(KEYINPUT72), .Z(n444) );
  NAND2_X1 U503 ( .A1(G229GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U506 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U507 ( .A(n450), .B(n449), .Z(n559) );
  AND2_X1 U508 ( .A1(n580), .A2(n559), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n451), .B(KEYINPUT76), .ZN(n466) );
  NAND2_X1 U510 ( .A1(n477), .A2(n466), .ZN(n452) );
  XNOR2_X1 U511 ( .A(KEYINPUT101), .B(n452), .ZN(n461) );
  NAND2_X1 U512 ( .A1(n461), .A2(n552), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U514 ( .A(G1GAT), .B(n455), .Z(G1324GAT) );
  XOR2_X1 U515 ( .A(G8GAT), .B(KEYINPUT103), .Z(n457) );
  NAND2_X1 U516 ( .A1(n461), .A2(n546), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n457), .B(n456), .ZN(G1325GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT35), .B(KEYINPUT104), .Z(n459) );
  NAND2_X1 U519 ( .A1(n461), .A2(n557), .ZN(n458) );
  XNOR2_X1 U520 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U521 ( .A(G15GAT), .B(n460), .ZN(G1326GAT) );
  NAND2_X1 U522 ( .A1(n519), .A2(n461), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n462), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U524 ( .A(KEYINPUT36), .B(n543), .Z(n587) );
  NAND2_X1 U525 ( .A1(n587), .A2(n463), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n566), .A2(n464), .ZN(n465) );
  XOR2_X1 U527 ( .A(KEYINPUT37), .B(n465), .Z(n487) );
  NAND2_X1 U528 ( .A1(n466), .A2(n487), .ZN(n467) );
  XNOR2_X1 U529 ( .A(n467), .B(KEYINPUT38), .ZN(n468) );
  XNOR2_X1 U530 ( .A(KEYINPUT105), .B(n468), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n552), .A2(n475), .ZN(n470) );
  XOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT39), .Z(n469) );
  XNOR2_X1 U533 ( .A(n470), .B(n469), .ZN(G1328GAT) );
  NAND2_X1 U534 ( .A1(n475), .A2(n546), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n471), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n473) );
  NAND2_X1 U537 ( .A1(n475), .A2(n557), .ZN(n472) );
  XNOR2_X1 U538 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U539 ( .A(G43GAT), .B(n474), .Z(G1330GAT) );
  NAND2_X1 U540 ( .A1(n475), .A2(n519), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n476), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U542 ( .A(n580), .B(KEYINPUT41), .Z(n537) );
  NOR2_X1 U543 ( .A1(n559), .A2(n537), .ZN(n486) );
  NAND2_X1 U544 ( .A1(n477), .A2(n486), .ZN(n483) );
  NOR2_X1 U545 ( .A1(n478), .A2(n483), .ZN(n479) );
  XOR2_X1 U546 ( .A(G57GAT), .B(n479), .Z(n480) );
  XNOR2_X1 U547 ( .A(KEYINPUT42), .B(n480), .ZN(G1332GAT) );
  NOR2_X1 U548 ( .A1(n492), .A2(n483), .ZN(n481) );
  XOR2_X1 U549 ( .A(G64GAT), .B(n481), .Z(G1333GAT) );
  NOR2_X1 U550 ( .A1(n495), .A2(n483), .ZN(n482) );
  XOR2_X1 U551 ( .A(G71GAT), .B(n482), .Z(G1334GAT) );
  NOR2_X1 U552 ( .A1(n500), .A2(n483), .ZN(n485) );
  XNOR2_X1 U553 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n484) );
  XNOR2_X1 U554 ( .A(n485), .B(n484), .ZN(G1335GAT) );
  NAND2_X1 U555 ( .A1(n487), .A2(n486), .ZN(n499) );
  INV_X1 U556 ( .A(n499), .ZN(n488) );
  NAND2_X1 U557 ( .A1(n489), .A2(n488), .ZN(n491) );
  NAND2_X1 U558 ( .A1(G85GAT), .A2(n499), .ZN(n490) );
  NAND2_X1 U559 ( .A1(n491), .A2(n490), .ZN(G1336GAT) );
  NOR2_X1 U560 ( .A1(n492), .A2(n499), .ZN(n494) );
  XNOR2_X1 U561 ( .A(G92GAT), .B(KEYINPUT107), .ZN(n493) );
  XNOR2_X1 U562 ( .A(n494), .B(n493), .ZN(G1337GAT) );
  NOR2_X1 U563 ( .A1(n495), .A2(n499), .ZN(n497) );
  XNOR2_X1 U564 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n496) );
  XNOR2_X1 U565 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U566 ( .A(G99GAT), .B(n498), .ZN(G1338GAT) );
  NOR2_X1 U567 ( .A1(n500), .A2(n499), .ZN(n502) );
  XNOR2_X1 U568 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n501) );
  XNOR2_X1 U569 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U570 ( .A(G106GAT), .B(n503), .Z(G1339GAT) );
  INV_X1 U571 ( .A(n559), .ZN(n574) );
  NOR2_X1 U572 ( .A1(n574), .A2(n537), .ZN(n504) );
  XOR2_X1 U573 ( .A(n504), .B(KEYINPUT46), .Z(n506) );
  NOR2_X1 U574 ( .A1(n566), .A2(n569), .ZN(n505) );
  NAND2_X1 U575 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n507), .B(KEYINPUT47), .ZN(n513) );
  XOR2_X1 U577 ( .A(KEYINPUT67), .B(KEYINPUT45), .Z(n509) );
  NAND2_X1 U578 ( .A1(n566), .A2(n587), .ZN(n508) );
  XNOR2_X1 U579 ( .A(n509), .B(n508), .ZN(n511) );
  NAND2_X1 U580 ( .A1(n574), .A2(n580), .ZN(n510) );
  NOR2_X1 U581 ( .A1(n511), .A2(n510), .ZN(n512) );
  NOR2_X1 U582 ( .A1(n513), .A2(n512), .ZN(n515) );
  NOR2_X1 U583 ( .A1(n548), .A2(n516), .ZN(n535) );
  NAND2_X1 U584 ( .A1(n535), .A2(n557), .ZN(n517) );
  XOR2_X1 U585 ( .A(KEYINPUT111), .B(n517), .Z(n518) );
  NOR2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n559), .A2(n532), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(KEYINPUT112), .ZN(n521) );
  XNOR2_X1 U589 ( .A(G113GAT), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n523) );
  INV_X1 U591 ( .A(n537), .ZN(n561) );
  NAND2_X1 U592 ( .A1(n532), .A2(n561), .ZN(n522) );
  XNOR2_X1 U593 ( .A(n523), .B(n522), .ZN(n525) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT113), .Z(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n527) );
  NAND2_X1 U597 ( .A1(n532), .A2(n566), .ZN(n526) );
  XNOR2_X1 U598 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n530) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n529) );
  XNOR2_X1 U602 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U603 ( .A(KEYINPUT116), .B(n531), .Z(n534) );
  NAND2_X1 U604 ( .A1(n532), .A2(n569), .ZN(n533) );
  XNOR2_X1 U605 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n535), .A2(n572), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n574), .A2(n542), .ZN(n536) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n536), .Z(G1344GAT) );
  NOR2_X1 U609 ( .A1(n537), .A2(n542), .ZN(n539) );
  XNOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n538) );
  XNOR2_X1 U611 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(n540), .ZN(G1345GAT) );
  NOR2_X1 U613 ( .A1(n584), .A2(n542), .ZN(n541) );
  XOR2_X1 U614 ( .A(G155GAT), .B(n541), .Z(G1346GAT) );
  NOR2_X1 U615 ( .A1(n543), .A2(n542), .ZN(n545) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n544) );
  XNOR2_X1 U617 ( .A(n545), .B(n544), .ZN(G1347GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n555) );
  INV_X1 U619 ( .A(KEYINPUT54), .ZN(n550) );
  XOR2_X1 U620 ( .A(n546), .B(KEYINPUT120), .Z(n547) );
  NOR2_X1 U621 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U622 ( .A(n550), .B(n549), .ZN(n551) );
  NAND2_X1 U623 ( .A1(n573), .A2(n553), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n556), .B(KEYINPUT55), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n568), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(G176GAT), .B(KEYINPUT57), .Z(n563) );
  NAND2_X1 U629 ( .A1(n568), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(n571), .ZN(G1351GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n586) );
  NOR2_X1 U639 ( .A1(n574), .A2(n586), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(KEYINPUT124), .B(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n586), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n586), .ZN(n585) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n585), .Z(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n590) );
  INV_X1 U652 ( .A(n586), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

