//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n207), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n218), .B(new_n219), .C1(new_n214), .C2(KEYINPUT64), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n209), .B(new_n213), .C1(new_n215), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  NOR4_X1   g021(.A1(new_n212), .A2(new_n205), .A3(new_n222), .A4(new_n208), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT24), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n225), .B2(new_n224), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n218), .A3(new_n219), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n221), .A2(new_n222), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n230));
  AOI21_X1  g029(.A(G190gat), .B1(new_n230), .B2(KEYINPUT66), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT27), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT67), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT27), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n233), .A2(new_n236), .A3(KEYINPUT67), .A4(new_n217), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT28), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT68), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n233), .A2(new_n236), .A3(new_n217), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n243), .A2(new_n244), .A3(new_n238), .A4(new_n237), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(KEYINPUT28), .A3(new_n217), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n240), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(new_n208), .A2(KEYINPUT26), .A3(new_n204), .ZN(new_n249));
  INV_X1    g048(.A(new_n224), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n204), .A2(KEYINPUT26), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n229), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n203), .B1(new_n253), .B2(KEYINPUT29), .ZN(new_n254));
  INV_X1    g053(.A(new_n252), .ZN(new_n255));
  INV_X1    g054(.A(new_n247), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n243), .A2(new_n238), .A3(new_n237), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT68), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n255), .B1(new_n258), .B2(new_n245), .ZN(new_n259));
  OAI211_X1 g058(.A(G226gat), .B(G233gat), .C1(new_n259), .C2(new_n229), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n262));
  OR2_X1    g061(.A1(G197gat), .A2(G204gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(G197gat), .A2(G204gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT73), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n265), .B2(new_n266), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT74), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n265), .A2(new_n271), .A3(new_n266), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n271), .B1(new_n265), .B2(new_n266), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n268), .B(new_n270), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT37), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n254), .A2(new_n275), .A3(new_n260), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n277), .A2(KEYINPUT85), .A3(new_n279), .A4(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n254), .A2(new_n275), .A3(new_n260), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n275), .B1(new_n254), .B2(new_n260), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT37), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G8gat), .B(G36gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G64gat), .B(G92gat), .ZN(new_n289));
  XOR2_X1   g088(.A(new_n288), .B(new_n289), .Z(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n202), .B1(new_n284), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(new_n202), .A3(new_n291), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(new_n282), .B2(new_n283), .ZN(new_n296));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n297), .B(KEYINPUT77), .Z(new_n298));
  INV_X1    g097(.A(G120gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G113gat), .ZN(new_n300));
  INV_X1    g099(.A(G113gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(G120gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT69), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n301), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n305));
  INV_X1    g104(.A(G134gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G127gat), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n305), .A2(new_n307), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT1), .B1(new_n300), .B2(new_n302), .ZN(new_n312));
  XNOR2_X1  g111(.A(G127gat), .B(G134gat), .ZN(new_n313));
  OAI22_X1  g112(.A1(new_n304), .A2(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI221_X1 g115(.A(KEYINPUT76), .B1(new_n312), .B2(new_n313), .C1(new_n304), .C2(new_n311), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT2), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n318), .A2(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n319));
  INV_X1    g118(.A(G155gat), .ZN(new_n320));
  INV_X1    g119(.A(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G141gat), .B(G148gat), .Z(new_n324));
  AOI21_X1  g123(.A(new_n318), .B1(G155gat), .B2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G141gat), .B(G148gat), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n322), .B(new_n319), .C1(new_n328), .C2(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n316), .A2(new_n317), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT78), .A4(new_n330), .ZN(new_n334));
  INV_X1    g133(.A(new_n330), .ZN(new_n335));
  INV_X1    g134(.A(new_n311), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n300), .A2(new_n302), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n310), .ZN(new_n339));
  INV_X1    g138(.A(new_n313), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n336), .A2(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n298), .B1(new_n333), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n341), .A2(new_n345), .A3(new_n327), .A4(new_n329), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT4), .B1(new_n330), .B2(new_n314), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n327), .A2(new_n329), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n349), .A2(new_n316), .A3(new_n317), .A4(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n298), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n348), .A2(new_n352), .A3(KEYINPUT5), .A4(new_n353), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n344), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n344), .A2(new_n356), .A3(KEYINPUT84), .A4(new_n357), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n360), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT6), .B1(new_n358), .B2(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n358), .A2(new_n365), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT6), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n277), .A2(new_n279), .A3(new_n290), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n294), .A2(new_n296), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n274), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n267), .B1(new_n376), .B2(new_n272), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n350), .B1(new_n377), .B2(KEYINPUT29), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n351), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n378), .A2(new_n330), .B1(new_n276), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(G228gat), .A2(G233gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT81), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT3), .B1(new_n275), .B2(new_n379), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n335), .ZN(new_n387));
  INV_X1    g186(.A(new_n382), .ZN(new_n388));
  INV_X1    g187(.A(new_n380), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(new_n275), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n385), .A2(new_n391), .A3(KEYINPUT82), .A4(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n394));
  OAI22_X1  g193(.A1(new_n381), .A2(new_n384), .B1(new_n387), .B2(new_n390), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(G22gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(G22gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n393), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT31), .B(G50gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT80), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n392), .A3(new_n391), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n401), .B1(new_n395), .B2(G22gat), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n398), .A2(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n348), .A2(new_n352), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n298), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n365), .B1(new_n408), .B2(KEYINPUT39), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n334), .A2(new_n342), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n331), .A2(new_n332), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n353), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n411), .A2(KEYINPUT83), .A3(new_n353), .A4(new_n412), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n408), .A2(KEYINPUT39), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT40), .B(new_n410), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT40), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n415), .B2(new_n416), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n409), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n422), .A3(new_n368), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n291), .B1(new_n285), .B2(new_n286), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n373), .A3(KEYINPUT30), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n277), .A2(new_n426), .A3(new_n279), .A4(new_n290), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n406), .B1(new_n423), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT86), .B1(new_n375), .B2(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n370), .A2(new_n372), .A3(new_n373), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n287), .A2(new_n202), .A3(new_n291), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n284), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n292), .B1(new_n282), .B2(new_n283), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n431), .B(new_n433), .C1(new_n434), .C2(new_n202), .ZN(new_n435));
  INV_X1    g234(.A(new_n428), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n419), .A2(new_n368), .A3(new_n422), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n405), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n369), .B1(new_n365), .B2(new_n358), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n372), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n428), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(new_n405), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT34), .ZN(new_n445));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT71), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n341), .B1(new_n259), .B2(new_n229), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n248), .A2(new_n252), .ZN(new_n451));
  INV_X1    g250(.A(new_n229), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n314), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n449), .B1(new_n454), .B2(new_n446), .ZN(new_n455));
  INV_X1    g254(.A(new_n446), .ZN(new_n456));
  AOI211_X1 g255(.A(new_n456), .B(new_n448), .C1(new_n450), .C2(new_n453), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n453), .A3(new_n456), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT32), .ZN(new_n460));
  XOR2_X1   g259(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g261(.A(G15gat), .B(G43gat), .Z(new_n463));
  XNOR2_X1  g262(.A(G71gat), .B(G99gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n465), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n459), .B(KEYINPUT32), .C1(new_n461), .C2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT72), .B(new_n458), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n446), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n448), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n446), .A3(new_n449), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT72), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT72), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n455), .B2(new_n457), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n474), .A2(new_n476), .A3(new_n468), .A4(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n470), .A2(new_n478), .A3(KEYINPUT36), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(new_n478), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n444), .A2(new_n479), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n430), .A2(new_n440), .A3(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n406), .A2(new_n428), .A3(new_n480), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT35), .B1(new_n370), .B2(new_n372), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n406), .A2(new_n480), .A3(new_n442), .A4(new_n428), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(KEYINPUT35), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G134gat), .B(G162gat), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  INV_X1    g293(.A(KEYINPUT99), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(KEYINPUT15), .ZN(new_n498));
  NAND2_X1  g297(.A1(G29gat), .A2(G36gat), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT90), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT14), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT91), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n502), .B(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n501), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n497), .A2(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n497), .A2(KEYINPUT89), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n510), .A2(KEYINPUT15), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n500), .B2(new_n506), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(KEYINPUT17), .A3(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT93), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT92), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT17), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(new_n520), .A3(new_n514), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT96), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g322(.A(G85gat), .ZN(new_n524));
  INV_X1    g323(.A(G92gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n523), .A2(new_n526), .ZN(new_n528));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529));
  AOI22_X1  g328(.A1(KEYINPUT8), .A2(new_n529), .B1(new_n524), .B2(new_n525), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G99gat), .B(G106gat), .Z(new_n532));
  OR2_X1    g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(KEYINPUT97), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT97), .B1(new_n533), .B2(new_n534), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n516), .B(new_n522), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n537), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n518), .A2(new_n521), .A3(new_n535), .A4(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT98), .ZN(new_n541));
  NAND3_X1  g340(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G190gat), .B(G218gat), .Z(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n546), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n538), .B(new_n548), .C1(new_n543), .C2(new_n544), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n496), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n494), .A2(new_n495), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n547), .A2(new_n549), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G57gat), .B(G64gat), .Z(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n560), .A2(new_n556), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n555), .B(new_n558), .C1(new_n561), .C2(KEYINPUT94), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n558), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n556), .A2(new_n560), .B1(new_n558), .B2(KEYINPUT94), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G127gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT16), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n572), .B2(G1gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n573), .B1(G1gat), .B2(new_n571), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G8gat), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(KEYINPUT21), .B2(new_n566), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT95), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n570), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(new_n320), .ZN(new_n580));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n578), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n533), .A2(new_n534), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n566), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n533), .A2(new_n562), .A3(new_n565), .A4(new_n534), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(G230gat), .ZN(new_n588));
  INV_X1    g387(.A(G233gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n566), .A2(KEYINPUT10), .ZN(new_n592));
  NOR3_X1   g391(.A1(new_n536), .A2(new_n537), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT10), .B1(new_n585), .B2(new_n586), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n591), .B1(new_n595), .B2(new_n590), .ZN(new_n596));
  XOR2_X1   g395(.A(G120gat), .B(G148gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT100), .ZN(new_n598));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  NOR2_X1   g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n600), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n554), .A2(new_n583), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n575), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n516), .A2(new_n607), .A3(new_n522), .ZN(new_n608));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n518), .A2(new_n521), .A3(new_n575), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n518), .A2(new_n521), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n607), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n610), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n609), .B(KEYINPUT13), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n608), .A2(KEYINPUT18), .A3(new_n609), .A4(new_n610), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n613), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G169gat), .B(G197gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT88), .ZN(new_n622));
  XOR2_X1   g421(.A(G113gat), .B(G141gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n620), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n618), .A3(new_n627), .A4(new_n619), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n606), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n491), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n442), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT101), .B(G1gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1324gat));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  NAND4_X1  g438(.A1(new_n634), .A2(KEYINPUT42), .A3(new_n436), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(new_n436), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT102), .ZN(new_n642));
  INV_X1    g441(.A(new_n639), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n642), .A2(KEYINPUT103), .A3(G8gat), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT103), .B1(new_n642), .B2(G8gat), .ZN(new_n646));
  OAI221_X1 g445(.A(new_n640), .B1(new_n644), .B2(KEYINPUT42), .C1(new_n645), .C2(new_n646), .ZN(G1325gat));
  AOI21_X1  g446(.A(G15gat), .B1(new_n634), .B2(new_n480), .ZN(new_n648));
  INV_X1    g447(.A(new_n482), .ZN(new_n649));
  INV_X1    g448(.A(new_n479), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(G15gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT104), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n648), .B1(new_n654), .B2(new_n634), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT105), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n634), .A2(new_n405), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT43), .B(G22gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  AOI21_X1  g458(.A(new_n554), .B1(new_n485), .B2(new_n490), .ZN(new_n660));
  INV_X1    g459(.A(new_n583), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n631), .A2(new_n661), .A3(new_n605), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n664), .A2(G29gat), .A3(new_n442), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT45), .Z(new_n666));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n435), .A2(new_n438), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n483), .B1(new_n668), .B2(KEYINPUT86), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n489), .B1(new_n669), .B2(new_n440), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n670), .B2(new_n554), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n491), .A2(KEYINPUT44), .A3(new_n553), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n662), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G29gat), .B1(new_n675), .B2(new_n442), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n666), .A2(new_n676), .ZN(G1328gat));
  OAI21_X1  g476(.A(G36gat), .B1(new_n675), .B2(new_n428), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n664), .A2(G36gat), .A3(new_n428), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT46), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(G1329gat));
  NAND2_X1  g480(.A1(new_n674), .A2(new_n652), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G43gat), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT106), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT47), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n480), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n664), .A2(G43gat), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  OAI211_X1 g488(.A(new_n683), .B(new_n687), .C1(new_n684), .C2(KEYINPUT47), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  INV_X1    g490(.A(KEYINPUT48), .ZN(new_n692));
  INV_X1    g491(.A(new_n664), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n406), .A2(G50gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT107), .Z(new_n696));
  NAND4_X1  g495(.A1(new_n671), .A2(new_n672), .A3(new_n405), .A4(new_n663), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n697), .A2(G50gat), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n692), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(G50gat), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n701), .B2(new_n697), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n695), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n693), .A2(KEYINPUT108), .A3(new_n694), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n692), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n703), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n708), .B1(new_n703), .B2(new_n707), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n699), .B1(new_n709), .B2(new_n710), .ZN(G1331gat));
  NOR4_X1   g510(.A1(new_n553), .A2(new_n631), .A3(new_n661), .A4(new_n605), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n491), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n635), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g514(.A1(new_n713), .A2(new_n436), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n652), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n686), .A2(G71gat), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n721), .A2(G71gat), .B1(new_n713), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n713), .A2(new_n405), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(new_n631), .B2(new_n583), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n661), .A2(KEYINPUT111), .A3(new_n629), .A4(new_n630), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT112), .B1(new_n730), .B2(new_n604), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n732), .B(new_n605), .C1(new_n728), .C2(new_n729), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n673), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n442), .ZN(new_n736));
  AND3_X1   g535(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n439), .B1(new_n435), .B2(new_n438), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n737), .A2(new_n738), .A3(new_n483), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT113), .B(new_n553), .C1(new_n739), .C2(new_n489), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n730), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n660), .A2(KEYINPUT113), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT51), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n730), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n660), .B2(KEYINPUT113), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n670), .B2(new_n554), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n604), .A2(new_n524), .A3(new_n635), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n736), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  NOR3_X1   g551(.A1(new_n605), .A2(G92gat), .A3(new_n428), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n743), .A2(new_n749), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n731), .A2(new_n733), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n671), .A2(new_n755), .A3(new_n672), .A4(new_n436), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT52), .B1(new_n756), .B2(G92gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT116), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n754), .A2(new_n760), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g561(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n730), .A2(new_n748), .A3(new_n740), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n745), .B2(new_n748), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n753), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n756), .A2(G92gat), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT115), .B1(new_n768), .B2(KEYINPUT52), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  AOI211_X1 g570(.A(new_n770), .B(new_n771), .C1(new_n766), .C2(new_n767), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n762), .B1(new_n769), .B2(new_n772), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n735), .B2(new_n651), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n686), .A2(new_n605), .A3(G99gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n750), .B2(new_n775), .ZN(G1338gat));
  NAND2_X1  g575(.A1(new_n734), .A2(new_n405), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n764), .A2(new_n765), .ZN(new_n779));
  OR3_X1    g578(.A1(new_n605), .A2(new_n406), .A3(G106gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n777), .B2(G106gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n750), .B2(new_n780), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(G1339gat));
  INV_X1    g585(.A(KEYINPUT119), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n539), .A2(KEYINPUT10), .A3(new_n566), .A4(new_n535), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n587), .B2(KEYINPUT10), .ZN(new_n790));
  INV_X1    g589(.A(new_n590), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n788), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n595), .B2(new_n590), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT118), .A4(new_n791), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n791), .B1(new_n593), .B2(new_n594), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n600), .B1(new_n797), .B2(KEYINPUT54), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n602), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT118), .B1(new_n790), .B2(new_n791), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n595), .A2(new_n793), .A3(new_n590), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n798), .B1(new_n805), .B2(new_n792), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(KEYINPUT55), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n787), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n601), .B1(new_n806), .B2(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n800), .A2(new_n801), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(KEYINPUT119), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n811), .A3(new_n631), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n616), .A2(new_n617), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n626), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n630), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n604), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n553), .B1(new_n812), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n808), .A2(new_n553), .A3(new_n811), .A4(new_n816), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n661), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n606), .A2(new_n631), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n442), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n486), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n632), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(new_n301), .ZN(G1340gat));
  NOR2_X1   g626(.A1(new_n825), .A2(new_n605), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(new_n299), .ZN(G1341gat));
  AOI21_X1  g628(.A(new_n661), .B1(KEYINPUT120), .B2(new_n308), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n824), .A2(new_n486), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n308), .A2(KEYINPUT120), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(G1342gat));
  NOR2_X1   g632(.A1(new_n686), .A2(new_n405), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n554), .A2(new_n436), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n824), .A2(new_n306), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT56), .Z(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n825), .B2(new_n554), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(G1343gat));
  NAND3_X1  g638(.A1(new_n651), .A2(new_n635), .A3(new_n428), .ZN(new_n840));
  XNOR2_X1  g639(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n809), .B1(new_n806), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n817), .B1(new_n632), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n554), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n583), .B1(new_n844), .B2(new_n819), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n405), .B1(new_n845), .B2(new_n822), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n840), .B1(new_n846), .B2(KEYINPUT57), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n406), .B1(new_n821), .B2(new_n823), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n632), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n652), .A2(new_n406), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n824), .A2(new_n428), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(G141gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n631), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT58), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n852), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1344gat));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n863), .B(G148gat), .C1(new_n851), .C2(new_n605), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n553), .A2(new_n816), .A3(new_n809), .A4(new_n810), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n583), .B1(new_n844), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n849), .B(new_n405), .C1(new_n867), .C2(new_n822), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n840), .A2(new_n605), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n868), .B(new_n869), .C1(new_n848), .C2(new_n849), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(G148gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n865), .B1(new_n871), .B2(KEYINPUT59), .ZN(new_n872));
  AOI211_X1 g671(.A(KEYINPUT122), .B(new_n863), .C1(new_n870), .C2(G148gat), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n864), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR3_X1    g673(.A1(new_n854), .A2(G148gat), .A3(new_n605), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1345gat));
  OAI21_X1  g675(.A(G155gat), .B1(new_n851), .B2(new_n661), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n320), .A3(new_n583), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n851), .B2(new_n554), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n824), .A2(new_n321), .A3(new_n835), .A4(new_n853), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n635), .A2(new_n428), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n821), .B2(new_n823), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n834), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n631), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(G169gat), .ZN(G1348gat));
  AOI21_X1  g687(.A(new_n605), .B1(KEYINPUT123), .B2(new_n207), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n207), .A2(KEYINPUT123), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(G1349gat));
  NAND3_X1  g691(.A1(new_n885), .A2(new_n834), .A3(new_n583), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT124), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n885), .A2(new_n895), .A3(new_n834), .A4(new_n583), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(G183gat), .A3(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT60), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n885), .A2(new_n246), .A3(new_n834), .A4(new_n583), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(KEYINPUT60), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n897), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n899), .B1(new_n897), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(G1350gat));
  NOR2_X1   g704(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n886), .B2(new_n553), .ZN(new_n907));
  NAND2_X1  g706(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n907), .B(new_n908), .Z(G1351gat));
  AND2_X1   g708(.A1(new_n885), .A2(new_n853), .ZN(new_n910));
  XNOR2_X1  g709(.A(KEYINPUT126), .B(G197gat), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n631), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n652), .A2(new_n884), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n868), .B(new_n913), .C1(new_n848), .C2(new_n849), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(new_n632), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n911), .ZN(G1352gat));
  INV_X1    g715(.A(G204gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n910), .A2(new_n917), .A3(new_n604), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n919));
  OAI21_X1  g718(.A(G204gat), .B1(new_n914), .B2(new_n605), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(KEYINPUT62), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(G1353gat));
  INV_X1    g721(.A(G211gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n910), .A2(new_n923), .A3(new_n583), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G211gat), .B1(new_n914), .B2(new_n661), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT63), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(KEYINPUT63), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n928), .A3(new_n929), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n914), .B2(new_n554), .ZN(new_n931));
  INV_X1    g730(.A(G218gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n910), .A2(new_n932), .A3(new_n553), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1355gat));
endmodule


