//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT92), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  OR3_X1    g003(.A1(new_n204), .A2(KEYINPUT94), .A3(G1gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT93), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n207), .A2(G1gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT94), .B1(new_n204), .B2(G1gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n205), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G8gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n204), .A2(G1gat), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n204), .A2(new_n208), .B1(new_n206), .B2(G8gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g017(.A(G43gat), .B(G50gat), .Z(new_n219));
  INV_X1    g018(.A(KEYINPUT15), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n219), .A2(new_n220), .B1(G29gat), .B2(G36gat), .ZN(new_n221));
  NOR3_X1   g020(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n222));
  XOR2_X1   g021(.A(new_n222), .B(KEYINPUT91), .Z(new_n223));
  OAI21_X1  g022(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  OAI221_X1 g024(.A(new_n221), .B1(new_n220), .B2(new_n219), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n219), .A2(new_n220), .ZN(new_n227));
  INV_X1    g026(.A(G29gat), .ZN(new_n228));
  INV_X1    g027(.A(G36gat), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n225), .A2(new_n222), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n218), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n234), .B(KEYINPUT13), .Z(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(KEYINPUT95), .A3(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n218), .A2(new_n232), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n212), .A2(new_n217), .B1(new_n231), .B2(new_n226), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n235), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT95), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n236), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n232), .B(KEYINPUT17), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n211), .A2(G8gat), .B1(new_n216), .B2(new_n215), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n218), .A2(new_n232), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n234), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT18), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n245), .A2(new_n246), .A3(new_n249), .A4(new_n234), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G113gat), .B(G141gat), .ZN(new_n252));
  INV_X1    g051(.A(G197gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT11), .B(G169gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n256), .B(KEYINPUT12), .Z(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n242), .A2(new_n251), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n242), .B2(new_n251), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G71gat), .A2(G78gat), .ZN(new_n262));
  OR2_X1    g061(.A1(G71gat), .A2(G78gat), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT9), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(G57gat), .B(G64gat), .Z(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT96), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(KEYINPUT9), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n262), .A3(new_n263), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT21), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n272), .A2(new_n273), .ZN(new_n277));
  OAI21_X1  g076(.A(G183gat), .B1(new_n218), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n277), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n244), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n278), .B2(new_n281), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n276), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G127gat), .B(G155gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G231gat), .A2(G233gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n278), .A2(new_n281), .ZN(new_n290));
  INV_X1    g089(.A(new_n282), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(new_n283), .A3(new_n275), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n286), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n289), .B1(new_n286), .B2(new_n293), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT97), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT7), .ZN(new_n299));
  NAND2_X1  g098(.A1(G85gat), .A2(G92gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(G99gat), .A2(G106gat), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n299), .A2(new_n300), .B1(KEYINPUT8), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT97), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n298), .A2(KEYINPUT7), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n304), .A2(new_n305), .A3(G85gat), .A4(G92gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n302), .B(new_n306), .C1(G85gat), .C2(G92gat), .ZN(new_n307));
  XOR2_X1   g106(.A(G99gat), .B(G106gat), .Z(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n243), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n311));
  INV_X1    g110(.A(new_n309), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n232), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G134gat), .B(G162gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(KEYINPUT98), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n310), .A2(new_n318), .A3(new_n311), .A4(new_n313), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G190gat), .B(G218gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n317), .A2(new_n323), .A3(new_n319), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT99), .B1(new_n297), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n286), .A2(new_n293), .ZN(new_n329));
  INV_X1    g128(.A(new_n289), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(new_n294), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT99), .ZN(new_n333));
  INV_X1    g132(.A(new_n327), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n272), .A2(new_n309), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n272), .A2(new_n309), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G230gat), .A2(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT10), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n336), .A2(new_n341), .A3(new_n337), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT100), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n336), .A2(new_n341), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n336), .A2(KEYINPUT100), .A3(new_n341), .A4(new_n337), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n340), .B1(new_n347), .B2(new_n339), .ZN(new_n348));
  XNOR2_X1  g147(.A(G120gat), .B(G148gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT101), .ZN(new_n350));
  XNOR2_X1  g149(.A(G176gat), .B(G204gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT102), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n348), .B2(new_n353), .ZN(new_n355));
  INV_X1    g154(.A(new_n348), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(KEYINPUT102), .A3(new_n352), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n328), .A2(new_n335), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT84), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT82), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  XNOR2_X1  g161(.A(G141gat), .B(G148gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT2), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n363), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT75), .ZN(new_n370));
  INV_X1    g169(.A(G141gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n371), .A2(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n373), .A2(G141gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n366), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n364), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(new_n365), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n370), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(G141gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n371), .A2(G148gat), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT2), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G155gat), .B(G162gat), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n362), .B(new_n369), .C1(new_n378), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT76), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT75), .B1(new_n381), .B2(new_n382), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n377), .B(new_n370), .C1(new_n363), .C2(KEYINPUT2), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n368), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT76), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n362), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G211gat), .A2(G218gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT22), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G197gat), .B(G204gat), .ZN(new_n395));
  OR2_X1    g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT72), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n392), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n397), .B1(new_n396), .B2(new_n392), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n394), .B(new_n395), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n392), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n395), .A2(new_n394), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n404), .A3(new_n398), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT73), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n361), .B1(new_n391), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n386), .A2(new_n387), .ZN(new_n412));
  AND4_X1   g211(.A1(new_n389), .A2(new_n412), .A3(new_n362), .A4(new_n369), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n389), .B1(new_n388), .B2(new_n362), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n406), .A2(new_n408), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT82), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(new_n369), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n401), .B2(new_n405), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(KEYINPUT3), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n410), .A2(new_n417), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G228gat), .A2(G233gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n385), .A2(new_n390), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n409), .B1(new_n424), .B2(new_n411), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n411), .B1(new_n406), .B2(new_n408), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n388), .B1(new_n426), .B2(new_n362), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n425), .A2(new_n427), .A3(new_n422), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(G22gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n422), .B2(new_n421), .ZN(new_n433));
  INV_X1    g232(.A(new_n431), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(KEYINPUT31), .B(G50gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n437), .B(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT81), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n360), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n423), .A2(new_n434), .A3(new_n429), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n434), .B1(new_n423), .B2(new_n429), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n360), .B(new_n440), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n446));
  INV_X1    g245(.A(G22gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n433), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n430), .A2(KEYINPUT85), .A3(G22gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n439), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n442), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n435), .A2(KEYINPUT86), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI22_X1  g253(.A1(new_n441), .A2(new_n445), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT25), .ZN(new_n456));
  INV_X1    g255(.A(G190gat), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n457), .A2(KEYINPUT65), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(KEYINPUT65), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n279), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT24), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n456), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT23), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n467), .A2(G169gat), .A3(G176gat), .ZN(new_n468));
  NOR2_X1   g267(.A1(G169gat), .A2(G176gat), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G169gat), .ZN(new_n471));
  INV_X1    g270(.A(G176gat), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT23), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n468), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n470), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(KEYINPUT23), .ZN(new_n476));
  NOR2_X1   g275(.A1(G183gat), .A2(G190gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n463), .A2(new_n464), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n466), .A2(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT26), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n482), .B1(new_n471), .B2(new_n472), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n469), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n461), .B1(new_n470), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G183gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT65), .B(G190gat), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT28), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n489), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n487), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n486), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(G226gat), .A2(G233gat), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n481), .A2(new_n494), .B1(KEYINPUT29), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n460), .A2(new_n465), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT25), .A3(new_n474), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n478), .A2(new_n477), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n467), .B1(G169gat), .B2(G176gat), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n476), .B1(new_n500), .B2(new_n469), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n480), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n495), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n486), .A2(new_n490), .A3(new_n493), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n496), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n416), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n409), .A2(new_n496), .A3(new_n506), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G8gat), .B(G36gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(G64gat), .B(G92gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(KEYINPUT74), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n514), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n513), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n515), .A2(KEYINPUT74), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G1gat), .B(G29gat), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT0), .B(G57gat), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G120gat), .ZN(new_n527));
  INV_X1    g326(.A(G113gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT68), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G113gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n527), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n528), .A2(G120gat), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT69), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT69), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n527), .A2(G113gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT68), .B(G113gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n535), .B(new_n536), .C1(new_n537), .C2(new_n527), .ZN(new_n538));
  NOR2_X1   g337(.A1(G127gat), .A2(G134gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G127gat), .A2(G134gat), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT1), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n534), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n528), .A2(G120gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT67), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT1), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n536), .A2(new_n544), .A3(KEYINPUT67), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n551), .B1(new_n540), .B2(new_n541), .ZN(new_n552));
  INV_X1    g351(.A(new_n541), .ZN(new_n553));
  NOR3_X1   g352(.A1(new_n553), .A2(new_n539), .A3(KEYINPUT66), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n388), .A2(new_n543), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT4), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n388), .A2(new_n543), .A3(new_n556), .A4(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(KEYINPUT77), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n418), .A2(KEYINPUT3), .B1(new_n543), .B2(new_n556), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n562), .B1(new_n414), .B2(new_n413), .ZN(new_n563));
  NAND2_X1  g362(.A1(G225gat), .A2(G233gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n557), .A2(new_n565), .A3(KEYINPUT4), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n561), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n543), .A2(new_n556), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n418), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n569), .A2(new_n557), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n567), .B(KEYINPUT5), .C1(new_n564), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n558), .A2(KEYINPUT78), .A3(new_n560), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n573), .A3(KEYINPUT4), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n564), .ZN(new_n577));
  AOI211_X1 g376(.A(KEYINPUT5), .B(new_n577), .C1(new_n424), .C2(new_n562), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT79), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT5), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n580), .A3(new_n564), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT79), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n581), .A2(new_n575), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n526), .B(new_n571), .C1(new_n579), .C2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n571), .B1(new_n579), .B2(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n525), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT79), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n582), .B1(new_n581), .B2(new_n575), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n592), .A2(KEYINPUT80), .A3(new_n526), .A4(new_n571), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(KEYINPUT6), .A3(new_n525), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n520), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n568), .B1(new_n481), .B2(new_n494), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n503), .A2(new_n543), .A3(new_n556), .A4(new_n505), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n599), .A2(G227gat), .A3(G233gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G15gat), .B(G43gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G71gat), .B(G99gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT34), .ZN(new_n607));
  NAND2_X1  g406(.A1(G227gat), .A2(G233gat), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n597), .A2(new_n598), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT71), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT70), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n608), .B1(new_n599), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT70), .B1(new_n597), .B2(new_n598), .ZN(new_n613));
  OAI21_X1  g412(.A(KEYINPUT34), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n600), .A2(KEYINPUT32), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n610), .B2(new_n614), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n606), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n610), .A2(new_n614), .ZN(new_n619));
  INV_X1    g418(.A(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n606), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n455), .A2(new_n596), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT35), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n618), .A2(new_n624), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT90), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n618), .A2(new_n624), .A3(KEYINPUT90), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n520), .A2(KEYINPUT35), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n525), .B(KEYINPUT87), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n587), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n586), .A2(new_n636), .A3(new_n589), .A4(new_n593), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n595), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n455), .A2(new_n632), .A3(new_n633), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n509), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n641), .A2(KEYINPUT88), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT88), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n508), .B1(new_n509), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT37), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT37), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n508), .A2(new_n647), .A3(new_n509), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n645), .A2(new_n646), .A3(new_n513), .A4(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n409), .B1(new_n496), .B2(new_n506), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT37), .B1(new_n641), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n648), .A3(new_n513), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n652), .A2(KEYINPUT89), .A3(KEYINPUT38), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT89), .B1(new_n652), .B2(KEYINPUT38), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n649), .B(new_n514), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n656), .A2(new_n595), .A3(new_n637), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n576), .A2(new_n563), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n577), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n570), .A2(new_n564), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n660), .A2(KEYINPUT39), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n634), .B1(new_n660), .B2(KEYINPUT39), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n658), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n660), .A2(KEYINPUT39), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n666), .A2(KEYINPUT40), .A3(new_n634), .A4(new_n662), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n520), .A2(new_n665), .A3(new_n636), .A4(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n455), .A2(new_n657), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n448), .A2(new_n449), .A3(new_n439), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n430), .A2(KEYINPUT86), .A3(new_n431), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n451), .B1(new_n433), .B2(new_n434), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n671), .A2(new_n444), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n594), .A2(new_n595), .ZN(new_n677));
  INV_X1    g476(.A(new_n520), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n625), .B(KEYINPUT36), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n669), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  AOI211_X1 g481(.A(new_n261), .B(new_n359), .C1(new_n640), .C2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n677), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n520), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT16), .B(G8gat), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(G8gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(G1325gat));
  INV_X1    g492(.A(new_n681), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n683), .A2(G15gat), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n683), .A2(new_n632), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n695), .B1(new_n696), .B2(G15gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT103), .Z(G1326gat));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n676), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  AOI21_X1  g500(.A(new_n334), .B1(new_n640), .B2(new_n682), .ZN(new_n702));
  INV_X1    g501(.A(new_n358), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n703), .A2(new_n261), .A3(new_n332), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n228), .A3(new_n684), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT35), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n671), .A2(new_n444), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n672), .A2(new_n675), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n628), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n708), .B1(new_n711), .B2(new_n596), .ZN(new_n712));
  AND4_X1   g511(.A1(new_n455), .A2(new_n633), .A3(new_n632), .A4(new_n638), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n682), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n327), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n704), .ZN(new_n720));
  OAI21_X1  g519(.A(G29gat), .B1(new_n720), .B2(new_n677), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n707), .A2(new_n721), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n229), .A3(new_n520), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT46), .Z(new_n724));
  OAI21_X1  g523(.A(G36gat), .B1(new_n720), .B2(new_n678), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1329gat));
  NAND2_X1  g525(.A1(new_n705), .A2(new_n632), .ZN(new_n727));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n694), .A2(G43gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n720), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT47), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n729), .B(new_n733), .C1(new_n720), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(G1330gat));
  NAND4_X1  g534(.A1(new_n719), .A2(G50gat), .A3(new_n676), .A4(new_n704), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n705), .A2(new_n676), .ZN(new_n737));
  INV_X1    g536(.A(G50gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g540(.A1(new_n328), .A2(new_n261), .A3(new_n335), .A4(new_n703), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT104), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n714), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n677), .B(KEYINPUT105), .Z(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n744), .A2(new_n520), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n749), .B(new_n750), .Z(G1333gat));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n743), .A2(new_n632), .A3(new_n714), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n743), .A2(new_n755), .A3(new_n632), .A4(new_n714), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G71gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n744), .B2(new_n694), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n752), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(G71gat), .B1(new_n754), .B2(new_n756), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n763), .A2(KEYINPUT50), .A3(new_n760), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n762), .A2(new_n764), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n744), .A2(new_n676), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n242), .A2(new_n251), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n257), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n242), .A2(new_n251), .A3(new_n258), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n332), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n716), .B2(new_n718), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n775), .A2(G85gat), .A3(new_n684), .A4(new_n703), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n714), .A2(new_n327), .A3(new_n773), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n714), .A2(KEYINPUT51), .A3(new_n327), .A4(new_n773), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n358), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n684), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n768), .B(new_n776), .C1(new_n782), .C2(G85gat), .ZN(new_n783));
  AOI21_X1  g582(.A(G85gat), .B1(new_n781), .B2(new_n684), .ZN(new_n784));
  AOI211_X1 g583(.A(KEYINPUT44), .B(new_n334), .C1(new_n640), .C2(new_n682), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n717), .B1(new_n714), .B2(new_n327), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n703), .B(new_n773), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n787), .A2(new_n522), .A3(new_n677), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT107), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n789), .ZN(G1336gat));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n678), .A2(G92gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n781), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(G92gat), .B1(new_n787), .B2(new_n678), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT52), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n794), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n787), .B2(new_n681), .ZN(new_n800));
  INV_X1    g599(.A(G99gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n703), .A2(new_n632), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT109), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT51), .B1(new_n702), .B2(new_n773), .ZN(new_n804));
  AND4_X1   g603(.A1(KEYINPUT51), .A2(new_n714), .A3(new_n327), .A4(new_n773), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n800), .A2(new_n806), .ZN(G1338gat));
  OAI211_X1 g606(.A(new_n703), .B(new_n676), .C1(new_n804), .C2(new_n805), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n676), .A2(G106gat), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n775), .A2(KEYINPUT110), .A3(new_n703), .A4(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n811), .B2(new_n813), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(G1339gat));
  NAND2_X1  g616(.A1(new_n455), .A2(new_n632), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n348), .A2(new_n353), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n347), .A2(new_n339), .ZN(new_n820));
  INV_X1    g619(.A(new_n339), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n344), .A2(new_n821), .A3(new_n345), .A4(new_n346), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n347), .A2(new_n824), .A3(new_n339), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n352), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n820), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n352), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n772), .A2(new_n819), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n233), .A2(new_n235), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n234), .B1(new_n245), .B2(new_n246), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n256), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n355), .A2(new_n771), .A3(new_n357), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n327), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n830), .A2(new_n819), .A3(new_n826), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n327), .A2(new_n771), .A3(new_n834), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n297), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n328), .A2(new_n261), .A3(new_n335), .A4(new_n358), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n818), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n677), .A2(new_n520), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n772), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n846), .A2(KEYINPUT112), .A3(G113gat), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT112), .B1(new_n846), .B2(G113gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n835), .B1(new_n837), .B2(new_n261), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n839), .B1(new_n849), .B2(new_n334), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n841), .B1(new_n850), .B2(new_n332), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n745), .ZN(new_n852));
  INV_X1    g651(.A(new_n711), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT113), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT113), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n851), .A2(new_n855), .A3(new_n711), .A4(new_n745), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n678), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n261), .A2(new_n537), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n847), .A2(new_n848), .B1(new_n858), .B2(new_n859), .ZN(G1340gat));
  OAI21_X1  g659(.A(G120gat), .B1(new_n844), .B2(new_n358), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n854), .A2(new_n527), .A3(new_n678), .A4(new_n856), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n358), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT114), .ZN(G1341gat));
  NAND3_X1  g663(.A1(new_n845), .A2(G127gat), .A3(new_n332), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n845), .A2(KEYINPUT115), .A3(G127gat), .A4(new_n332), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n857), .A2(new_n332), .A3(new_n678), .ZN(new_n870));
  INV_X1    g669(.A(G127gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(G1342gat));
  NOR2_X1   g671(.A1(new_n334), .A2(G134gat), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n854), .A2(new_n678), .A3(new_n856), .A4(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n844), .B2(new_n334), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  OR2_X1    g677(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n851), .A2(new_n676), .ZN(new_n880));
  NAND2_X1  g679(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n681), .A2(new_n843), .ZN(new_n884));
  OR2_X1    g683(.A1(KEYINPUT116), .A2(KEYINPUT57), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n851), .A2(new_n676), .A3(new_n881), .A4(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n883), .A2(new_n772), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G141gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n681), .A2(new_n676), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n520), .B1(new_n890), .B2(KEYINPUT117), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(KEYINPUT117), .ZN(new_n893));
  NOR4_X1   g692(.A1(new_n852), .A2(G141gat), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n772), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n879), .A2(new_n888), .A3(new_n889), .A4(new_n895), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n887), .A2(G141gat), .B1(new_n894), .B2(new_n772), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n879), .B1(new_n897), .B2(new_n889), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n896), .A2(new_n898), .ZN(G1344gat));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n455), .B2(KEYINPUT119), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n851), .A2(new_n676), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n851), .B2(new_n676), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n703), .A3(new_n884), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n900), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT59), .B(new_n373), .C1(new_n908), .C2(new_n703), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n852), .A2(new_n893), .A3(new_n892), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n703), .A2(new_n373), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n907), .A2(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1345gat));
  NOR2_X1   g711(.A1(new_n910), .A2(new_n297), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n908), .A2(new_n332), .ZN(new_n914));
  MUX2_X1   g713(.A(new_n913), .B(new_n914), .S(G155gat), .Z(G1346gat));
  NOR2_X1   g714(.A1(new_n910), .A2(new_n334), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n908), .A2(new_n327), .ZN(new_n917));
  MUX2_X1   g716(.A(new_n916), .B(new_n917), .S(G162gat), .Z(G1347gat));
  NAND2_X1  g717(.A1(new_n851), .A2(new_n677), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n851), .A2(KEYINPUT120), .A3(new_n677), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n853), .A2(new_n678), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n471), .A3(new_n772), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n745), .A2(new_n678), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n842), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n261), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(new_n929), .ZN(G1348gat));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n472), .A3(new_n358), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n925), .A2(new_n703), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n472), .ZN(G1349gat));
  NOR2_X1   g732(.A1(new_n297), .A2(new_n488), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n924), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n936));
  OAI21_X1  g735(.A(G183gat), .B1(new_n928), .B2(new_n297), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(KEYINPUT121), .A2(KEYINPUT60), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(new_n939), .ZN(G1350gat));
  INV_X1    g739(.A(KEYINPUT122), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n941), .A3(new_n327), .A4(new_n491), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n491), .A3(new_n924), .ZN(new_n943));
  OAI21_X1  g742(.A(KEYINPUT122), .B1(new_n943), .B2(new_n334), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n842), .A2(new_n327), .A3(new_n927), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n946), .A2(G190gat), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n949), .B(new_n950), .Z(new_n951));
  NAND2_X1  g750(.A1(new_n945), .A2(new_n951), .ZN(G1351gat));
  NOR3_X1   g751(.A1(new_n745), .A2(new_n678), .A3(new_n694), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n905), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n772), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(G197gat), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n890), .A2(new_n678), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n923), .A2(new_n253), .A3(new_n772), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1352gat));
  INV_X1    g758(.A(new_n922), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT120), .B1(new_n851), .B2(new_n677), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n703), .B(new_n957), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT62), .B1(new_n962), .B2(G204gat), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OR3_X1    g764(.A1(new_n962), .A2(KEYINPUT62), .A3(G204gat), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n905), .A2(new_n703), .A3(new_n953), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G204gat), .ZN(new_n968));
  OAI211_X1 g767(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n962), .C2(G204gat), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n965), .A2(new_n966), .A3(new_n968), .A4(new_n969), .ZN(G1353gat));
  OAI211_X1 g769(.A(new_n332), .B(new_n953), .C1(new_n903), .C2(new_n904), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT63), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n971), .A2(G211gat), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n972), .A2(new_n973), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n297), .A2(G211gat), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n957), .B(new_n978), .C1(new_n960), .C2(new_n961), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n975), .A2(new_n976), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n977), .A2(new_n981), .A3(new_n982), .ZN(G1354gat));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n923), .A2(new_n327), .A3(new_n957), .ZN(new_n985));
  INV_X1    g784(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n984), .B1(new_n986), .B2(G218gat), .ZN(new_n987));
  INV_X1    g786(.A(G218gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n985), .A2(KEYINPUT127), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n334), .A2(new_n988), .ZN(new_n990));
  AOI22_X1  g789(.A1(new_n987), .A2(new_n989), .B1(new_n954), .B2(new_n990), .ZN(G1355gat));
endmodule


