// Benchmark "locked_c2670" written by ABC on Sat Dec 16 10:59:07 2023

module locked_c2670 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6,
    G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26,
    G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48,
    G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64,
    G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80,
    G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140,
    G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184,
    G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
    G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210,
    G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245,
    G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
    G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273,
    G274, G275, G276, G277, G278, G279, G452, G483, G543, G559, G567, G651,
    G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966,
    G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078,
    G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435,
    G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3,
    G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24,
    G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44,
    G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62,
    G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78,
    G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94,
    G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138,
    G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196,
    G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208,
    G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243,
    G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255,
    G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271,
    G272, G273, G274, G275, G276, G277, G278, G279, G452, G483, G543, G559,
    G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961,
    G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072,
    G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430,
    G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n372, new_n383, new_n387, new_n388, new_n389, new_n390, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n407, new_n408, new_n409,
    new_n410, new_n411, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n435, new_n436, new_n437, new_n438, new_n439, new_n440, new_n441,
    new_n442, new_n443, new_n446, new_n447, new_n448, new_n449, new_n451,
    new_n452, new_n453, new_n454, new_n455, new_n456, new_n457, new_n458,
    new_n460, new_n462, new_n463, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n478, new_n479, new_n480, new_n482, new_n483, new_n485, new_n486,
    new_n487, new_n488, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n501, new_n504, new_n506,
    new_n507, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n915, new_n916;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n372));
  INV_X1    g011(.A(new_n372), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n383));
  XOR2_X1   g022(.A(new_n383), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n372), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n387));
  XNOR2_X1  g026(.A(new_n387), .B(KEYINPUT2), .ZN(new_n388));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n389));
  INV_X1    g028(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g029(.A1(new_n388), .A2(new_n390), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n388), .A2(G2106), .B1(G567), .B2(new_n390), .ZN(G319));
  NAND2_X1  g032(.A1(G101), .A2(G2104), .ZN(new_n394));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n395));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n396));
  NOR2_X1   g035(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g036(.A(G137), .ZN(new_n398));
  OAI21_X1  g037(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g038(.A(G2105), .ZN(new_n400));
  NAND2_X1  g039(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n402));
  INV_X1    g041(.A(G125), .ZN(new_n403));
  OAI21_X1  g042(.A(new_n402), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g043(.A1(new_n404), .A2(G2105), .ZN(new_n405));
  AND2_X1   g044(.A1(new_n401), .A2(new_n405), .ZN(G160));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n407));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n408));
  NAND2_X1  g047(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI22_X1  g048(.A1(new_n409), .A2(G124), .B1(G112), .B2(G2104), .ZN(new_n410));
  AOI22_X1  g049(.A1(new_n409), .A2(G136), .B1(G100), .B2(G2104), .ZN(new_n411));
  MUX2_X1   g050(.A(new_n410), .B(new_n411), .S(new_n400), .Z(G162));
  AND2_X1   g051(.A1(G126), .A2(G2105), .ZN(new_n413));
  OAI21_X1  g052(.A(new_n413), .B1(new_n395), .B2(new_n396), .ZN(new_n414));
  NAND3_X1  g053(.A1(G114), .A2(G2104), .A3(G2105), .ZN(new_n415));
  NAND3_X1  g054(.A1(new_n400), .A2(G102), .A3(G2104), .ZN(new_n416));
  NAND3_X1  g055(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g056(.A(G2105), .B1(new_n407), .B2(new_n408), .ZN(new_n418));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n419));
  NAND3_X1  g058(.A1(new_n418), .A2(new_n419), .A3(G138), .ZN(new_n420));
  OAI211_X1 g059(.A(G138), .B(new_n400), .C1(new_n395), .C2(new_n396), .ZN(new_n421));
  NAND2_X1  g060(.A1(new_n421), .A2(KEYINPUT4), .ZN(new_n422));
  AOI21_X1  g061(.A(new_n417), .B1(new_n420), .B2(new_n422), .ZN(G164));
  XNOR2_X1  g062(.A(KEYINPUT5), .B(G543), .ZN(new_n424));
  AOI22_X1  g063(.A1(new_n424), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n425));
  AND2_X1   g064(.A1(KEYINPUT6), .A2(G651), .ZN(new_n426));
  NOR2_X1   g065(.A1(KEYINPUT6), .A2(G651), .ZN(new_n427));
  NOR2_X1   g066(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g067(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g068(.A1(new_n424), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n430));
  INV_X1    g069(.A(G651), .ZN(new_n431));
  NOR2_X1   g070(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OR2_X1    g071(.A1(new_n429), .A2(new_n432), .ZN(G303));
  INV_X1    g072(.A(G303), .ZN(G166));
  NAND2_X1  g073(.A1(G51), .A2(G543), .ZN(new_n435));
  XOR2_X1   g074(.A(KEYINPUT5), .B(G543), .Z(new_n436));
  INV_X1    g075(.A(G89), .ZN(new_n437));
  OAI21_X1  g076(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g077(.A(new_n428), .ZN(new_n439));
  NAND2_X1  g078(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g079(.A1(new_n424), .A2(G63), .A3(G651), .ZN(new_n441));
  NAND3_X1  g080(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n442));
  XNOR2_X1  g081(.A(new_n442), .B(KEYINPUT7), .ZN(new_n443));
  NAND3_X1  g082(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(G286));
  INV_X1    g083(.A(G286), .ZN(G168));
  AOI22_X1  g084(.A1(new_n424), .A2(G90), .B1(G52), .B2(G543), .ZN(new_n446));
  NOR2_X1   g085(.A1(new_n446), .A2(new_n428), .ZN(new_n447));
  AOI22_X1  g086(.A1(new_n424), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n448));
  NOR2_X1   g087(.A1(new_n448), .A2(new_n431), .ZN(new_n449));
  NOR2_X1   g088(.A1(new_n447), .A2(new_n449), .ZN(G171));
  AOI22_X1  g089(.A1(new_n439), .A2(G81), .B1(G56), .B2(G651), .ZN(new_n451));
  OR2_X1    g090(.A1(new_n451), .A2(new_n436), .ZN(new_n452));
  NAND2_X1  g091(.A1(G68), .A2(G651), .ZN(new_n453));
  INV_X1    g092(.A(G43), .ZN(new_n454));
  OAI21_X1  g093(.A(new_n453), .B1(new_n428), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g094(.A1(new_n455), .A2(G543), .ZN(new_n456));
  NAND2_X1  g095(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g096(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g097(.A1(new_n458), .A2(G860), .ZN(G153));
  AND3_X1   g098(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n460));
  NAND2_X1  g099(.A1(new_n460), .A2(G36), .ZN(G176));
  NAND2_X1  g100(.A1(G1), .A2(G3), .ZN(new_n462));
  XNOR2_X1  g101(.A(new_n462), .B(KEYINPUT8), .ZN(new_n463));
  NAND2_X1  g102(.A1(new_n460), .A2(new_n463), .ZN(G188));
  INV_X1    g103(.A(KEYINPUT9), .ZN(new_n465));
  AND2_X1   g104(.A1(G53), .A2(G543), .ZN(new_n466));
  NAND3_X1  g105(.A1(new_n439), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g106(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g107(.A(new_n465), .B1(new_n439), .B2(new_n466), .ZN(new_n469));
  NOR2_X1   g108(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g109(.A1(new_n439), .A2(G91), .A3(new_n424), .ZN(new_n471));
  NAND3_X1  g110(.A1(G78), .A2(G543), .A3(G651), .ZN(new_n472));
  NAND3_X1  g111(.A1(new_n424), .A2(G65), .A3(G651), .ZN(new_n473));
  NAND3_X1  g112(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g113(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g114(.A(new_n475), .ZN(G299));
  INV_X1    g115(.A(G171), .ZN(G301));
  OR2_X1    g116(.A1(new_n424), .A2(G74), .ZN(new_n478));
  NAND2_X1  g117(.A1(new_n478), .A2(G651), .ZN(new_n479));
  AOI22_X1  g118(.A1(new_n424), .A2(G87), .B1(G49), .B2(G543), .ZN(new_n480));
  OAI21_X1  g119(.A(new_n479), .B1(new_n480), .B2(new_n428), .ZN(G288));
  AOI22_X1  g120(.A1(new_n424), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n482));
  AOI22_X1  g121(.A1(new_n424), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n483));
  OAI22_X1  g122(.A1(new_n431), .A2(new_n482), .B1(new_n483), .B2(new_n428), .ZN(G305));
  AOI22_X1  g123(.A1(new_n424), .A2(G85), .B1(G47), .B2(G543), .ZN(new_n485));
  OR2_X1    g124(.A1(new_n485), .A2(new_n428), .ZN(new_n486));
  AOI22_X1  g125(.A1(new_n424), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n487));
  OR2_X1    g126(.A1(new_n487), .A2(new_n431), .ZN(new_n488));
  NAND2_X1  g127(.A1(new_n486), .A2(new_n488), .ZN(G290));
  NAND2_X1  g128(.A1(G301), .A2(G868), .ZN(new_n490));
  NAND3_X1  g129(.A1(new_n439), .A2(G92), .A3(new_n424), .ZN(new_n491));
  INV_X1    g130(.A(KEYINPUT10), .ZN(new_n492));
  XNOR2_X1  g131(.A(new_n491), .B(new_n492), .ZN(new_n493));
  AOI22_X1  g132(.A1(new_n424), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n494));
  OR2_X1    g133(.A1(new_n494), .A2(new_n431), .ZN(new_n495));
  NAND3_X1  g134(.A1(new_n439), .A2(G54), .A3(G543), .ZN(new_n496));
  NAND3_X1  g135(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g136(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g137(.A(new_n490), .B1(new_n498), .B2(G868), .ZN(G284));
  OAI21_X1  g138(.A(new_n490), .B1(new_n498), .B2(G868), .ZN(G321));
  NAND2_X1  g139(.A1(G286), .A2(G868), .ZN(new_n501));
  OAI21_X1  g140(.A(new_n501), .B1(new_n475), .B2(G868), .ZN(G297));
  OAI21_X1  g141(.A(new_n501), .B1(new_n475), .B2(G868), .ZN(G280));
  INV_X1    g142(.A(G559), .ZN(new_n504));
  OAI21_X1  g143(.A(new_n498), .B1(new_n504), .B2(G860), .ZN(G148));
  NAND2_X1  g144(.A1(new_n498), .A2(new_n504), .ZN(new_n506));
  NAND2_X1  g145(.A1(new_n506), .A2(G868), .ZN(new_n507));
  OAI21_X1  g146(.A(new_n507), .B1(G868), .B2(new_n458), .ZN(G323));
  XNOR2_X1  g147(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g148(.A1(new_n409), .A2(G135), .B1(G99), .B2(G2104), .ZN(new_n510));
  OR2_X1    g149(.A1(new_n510), .A2(G2105), .ZN(new_n511));
  AOI22_X1  g150(.A1(new_n409), .A2(G123), .B1(G111), .B2(G2104), .ZN(new_n512));
  OR2_X1    g151(.A1(new_n512), .A2(new_n400), .ZN(new_n513));
  NAND2_X1  g152(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g153(.A(new_n514), .B(G2096), .Z(new_n515));
  NAND3_X1  g154(.A1(new_n400), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n516));
  XOR2_X1   g155(.A(new_n516), .B(KEYINPUT12), .Z(new_n517));
  XOR2_X1   g156(.A(KEYINPUT13), .B(G2100), .Z(new_n518));
  XNOR2_X1  g157(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND2_X1  g158(.A1(new_n515), .A2(new_n519), .ZN(G156));
  XNOR2_X1  g159(.A(G2427), .B(G2430), .ZN(new_n521));
  XNOR2_X1  g160(.A(new_n521), .B(KEYINPUT15), .ZN(new_n522));
  XNOR2_X1  g161(.A(new_n522), .B(G2435), .ZN(new_n523));
  XOR2_X1   g162(.A(new_n523), .B(G2438), .Z(new_n524));
  NAND2_X1  g163(.A1(new_n524), .A2(KEYINPUT14), .ZN(new_n525));
  XNOR2_X1  g164(.A(G2451), .B(G2454), .ZN(new_n526));
  XNOR2_X1  g165(.A(new_n526), .B(KEYINPUT16), .ZN(new_n527));
  XNOR2_X1  g166(.A(G1341), .B(G1348), .ZN(new_n528));
  XNOR2_X1  g167(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g168(.A(G2443), .B(G2446), .ZN(new_n530));
  XOR2_X1   g169(.A(new_n529), .B(new_n530), .Z(new_n531));
  XNOR2_X1  g170(.A(new_n525), .B(new_n531), .ZN(new_n532));
  AND2_X1   g171(.A1(new_n532), .A2(G14), .ZN(G401));
  XOR2_X1   g172(.A(G2067), .B(G2678), .Z(new_n534));
  INV_X1    g173(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g174(.A(G2072), .B(G2078), .ZN(new_n536));
  XOR2_X1   g175(.A(G2084), .B(G2090), .Z(new_n537));
  NAND3_X1  g176(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  XOR2_X1   g177(.A(new_n538), .B(KEYINPUT18), .Z(new_n539));
  XNOR2_X1  g178(.A(new_n536), .B(KEYINPUT17), .ZN(new_n540));
  OR3_X1    g179(.A1(new_n540), .A2(new_n537), .A3(new_n534), .ZN(new_n541));
  AOI21_X1  g180(.A(new_n535), .B1(new_n540), .B2(new_n537), .ZN(new_n542));
  OAI21_X1  g181(.A(new_n542), .B1(new_n536), .B2(new_n537), .ZN(new_n543));
  NAND3_X1  g182(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g183(.A(new_n544), .B(G2096), .ZN(new_n545));
  XNOR2_X1  g184(.A(new_n545), .B(G2100), .ZN(new_n546));
  INV_X1    g185(.A(new_n546), .ZN(G227));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n548));
  XNOR2_X1  g187(.A(G1971), .B(G1976), .ZN(new_n549));
  XOR2_X1   g188(.A(new_n549), .B(KEYINPUT19), .Z(new_n550));
  XOR2_X1   g189(.A(G1961), .B(G1966), .Z(new_n551));
  INV_X1    g190(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g191(.A(new_n548), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g192(.A1(new_n550), .A2(new_n552), .ZN(new_n554));
  XOR2_X1   g193(.A(G1956), .B(G2474), .Z(new_n555));
  INV_X1    g194(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g195(.A(new_n553), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g196(.A(new_n550), .B1(new_n548), .B2(new_n552), .ZN(new_n558));
  OAI21_X1  g197(.A(new_n555), .B1(new_n551), .B2(KEYINPUT20), .ZN(new_n559));
  OAI21_X1  g198(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g199(.A(new_n554), .ZN(new_n561));
  OAI21_X1  g200(.A(new_n560), .B1(new_n561), .B2(new_n555), .ZN(new_n562));
  XOR2_X1   g201(.A(G1991), .B(G1996), .Z(new_n563));
  XNOR2_X1  g202(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g203(.A(G1981), .B(G1986), .Z(new_n565));
  XNOR2_X1  g204(.A(new_n565), .B(KEYINPUT21), .ZN(new_n566));
  XNOR2_X1  g205(.A(new_n566), .B(KEYINPUT22), .ZN(new_n567));
  XNOR2_X1  g206(.A(new_n564), .B(new_n567), .ZN(G229));
  INV_X1    g207(.A(G16), .ZN(new_n569));
  NAND2_X1  g208(.A1(new_n569), .A2(G22), .ZN(new_n570));
  OAI21_X1  g209(.A(new_n570), .B1(G166), .B2(new_n569), .ZN(new_n571));
  XOR2_X1   g210(.A(new_n571), .B(G1971), .Z(new_n572));
  NAND2_X1  g211(.A1(new_n569), .A2(G23), .ZN(new_n573));
  INV_X1    g212(.A(G288), .ZN(new_n574));
  OAI21_X1  g213(.A(new_n573), .B1(new_n574), .B2(new_n569), .ZN(new_n575));
  XNOR2_X1  g214(.A(KEYINPUT33), .B(G1976), .ZN(new_n576));
  XNOR2_X1  g215(.A(new_n575), .B(new_n576), .ZN(new_n577));
  MUX2_X1   g216(.A(G6), .B(G305), .S(G16), .Z(new_n578));
  XOR2_X1   g217(.A(KEYINPUT32), .B(G1981), .Z(new_n579));
  XNOR2_X1  g218(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND3_X1  g219(.A1(new_n572), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  OR2_X1    g220(.A1(new_n581), .A2(KEYINPUT34), .ZN(new_n582));
  NAND2_X1  g221(.A1(new_n569), .A2(G24), .ZN(new_n583));
  INV_X1    g222(.A(G290), .ZN(new_n584));
  OAI21_X1  g223(.A(new_n583), .B1(new_n584), .B2(new_n569), .ZN(new_n585));
  INV_X1    g224(.A(G1986), .ZN(new_n586));
  XNOR2_X1  g225(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g226(.A1(new_n581), .A2(KEYINPUT34), .ZN(new_n588));
  INV_X1    g227(.A(G29), .ZN(new_n589));
  NAND2_X1  g228(.A1(new_n589), .A2(G25), .ZN(new_n590));
  AOI22_X1  g229(.A1(new_n409), .A2(G119), .B1(G107), .B2(G2104), .ZN(new_n591));
  AOI22_X1  g230(.A1(new_n409), .A2(G131), .B1(G95), .B2(G2104), .ZN(new_n592));
  MUX2_X1   g231(.A(new_n591), .B(new_n592), .S(new_n400), .Z(new_n593));
  OAI21_X1  g232(.A(new_n590), .B1(new_n593), .B2(new_n589), .ZN(new_n594));
  XOR2_X1   g233(.A(KEYINPUT35), .B(G1991), .Z(new_n595));
  XNOR2_X1  g234(.A(new_n594), .B(new_n595), .ZN(new_n596));
  NAND4_X1  g235(.A1(new_n582), .A2(new_n587), .A3(new_n588), .A4(new_n596), .ZN(new_n597));
  XNOR2_X1  g236(.A(new_n597), .B(KEYINPUT36), .ZN(new_n598));
  NAND2_X1  g237(.A1(new_n589), .A2(G32), .ZN(new_n599));
  NAND3_X1  g238(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n600));
  XNOR2_X1  g239(.A(new_n600), .B(KEYINPUT26), .ZN(new_n601));
  INV_X1    g240(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g241(.A1(new_n409), .A2(G129), .A3(G2105), .ZN(new_n603));
  AOI22_X1  g242(.A1(new_n409), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n604));
  OAI211_X1 g243(.A(new_n602), .B(new_n603), .C1(new_n604), .C2(G2105), .ZN(new_n605));
  INV_X1    g244(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g245(.A(new_n599), .B1(new_n606), .B2(new_n589), .ZN(new_n607));
  XOR2_X1   g246(.A(new_n607), .B(KEYINPUT27), .Z(new_n608));
  XNOR2_X1  g247(.A(new_n608), .B(G1996), .ZN(new_n609));
  INV_X1    g248(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g249(.A1(new_n498), .A2(new_n569), .ZN(new_n611));
  AOI21_X1  g250(.A(new_n611), .B1(G4), .B2(new_n569), .ZN(new_n612));
  INV_X1    g251(.A(G1348), .ZN(new_n613));
  INV_X1    g252(.A(G2078), .ZN(new_n614));
  NAND2_X1  g253(.A1(new_n589), .A2(G27), .ZN(new_n615));
  OAI21_X1  g254(.A(new_n615), .B1(G164), .B2(new_n589), .ZN(new_n616));
  INV_X1    g255(.A(new_n616), .ZN(new_n617));
  OAI22_X1  g256(.A1(new_n612), .A2(new_n613), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  XNOR2_X1  g257(.A(KEYINPUT31), .B(G11), .ZN(new_n619));
  XNOR2_X1  g258(.A(KEYINPUT30), .B(G28), .ZN(new_n620));
  NAND2_X1  g259(.A1(new_n620), .A2(new_n589), .ZN(new_n621));
  OAI211_X1 g260(.A(new_n619), .B(new_n621), .C1(new_n514), .C2(new_n589), .ZN(new_n622));
  NAND2_X1  g261(.A1(new_n569), .A2(G5), .ZN(new_n623));
  OAI21_X1  g262(.A(new_n623), .B1(G171), .B2(new_n569), .ZN(new_n624));
  XNOR2_X1  g263(.A(new_n624), .B(G1961), .ZN(new_n625));
  NAND3_X1  g264(.A1(new_n400), .A2(G103), .A3(G2104), .ZN(new_n626));
  XOR2_X1   g265(.A(new_n626), .B(KEYINPUT25), .Z(new_n627));
  NAND3_X1  g266(.A1(G115), .A2(G2104), .A3(G2105), .ZN(new_n628));
  NAND2_X1  g267(.A1(new_n418), .A2(G139), .ZN(new_n629));
  NAND3_X1  g268(.A1(new_n409), .A2(G127), .A3(G2105), .ZN(new_n630));
  NAND4_X1  g269(.A1(new_n627), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(new_n631));
  MUX2_X1   g270(.A(G33), .B(new_n631), .S(G29), .Z(new_n632));
  XNOR2_X1  g271(.A(new_n632), .B(G2072), .ZN(new_n633));
  NOR4_X1   g272(.A1(new_n618), .A2(new_n622), .A3(new_n625), .A4(new_n633), .ZN(new_n634));
  OAI21_X1  g273(.A(new_n634), .B1(G2078), .B2(new_n616), .ZN(new_n635));
  NAND2_X1  g274(.A1(new_n569), .A2(G19), .ZN(new_n636));
  OAI21_X1  g275(.A(new_n636), .B1(new_n458), .B2(new_n569), .ZN(new_n637));
  NOR2_X1   g276(.A1(new_n637), .A2(G1341), .ZN(new_n638));
  NAND2_X1  g277(.A1(new_n612), .A2(new_n613), .ZN(new_n639));
  OR2_X1    g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n640));
  NAND2_X1  g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n641));
  NAND3_X1  g280(.A1(new_n640), .A2(new_n589), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g281(.A(new_n642), .B1(G160), .B2(new_n589), .ZN(new_n643));
  INV_X1    g282(.A(G2084), .ZN(new_n644));
  XNOR2_X1  g283(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g284(.A1(G286), .A2(G16), .ZN(new_n646));
  NAND2_X1  g285(.A1(new_n569), .A2(G21), .ZN(new_n647));
  AND2_X1   g286(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g287(.A(new_n648), .ZN(new_n649));
  AOI22_X1  g288(.A1(new_n649), .A2(G1966), .B1(new_n637), .B2(G1341), .ZN(new_n650));
  NAND3_X1  g289(.A1(new_n639), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g290(.A(KEYINPUT28), .B1(new_n589), .B2(G26), .ZN(new_n652));
  AND3_X1   g291(.A1(new_n589), .A2(KEYINPUT28), .A3(G26), .ZN(new_n653));
  AOI22_X1  g292(.A1(new_n409), .A2(G140), .B1(G104), .B2(G2104), .ZN(new_n654));
  NOR2_X1   g293(.A1(new_n654), .A2(G2105), .ZN(new_n655));
  AOI22_X1  g294(.A1(new_n409), .A2(G128), .B1(G116), .B2(G2104), .ZN(new_n656));
  NOR2_X1   g295(.A1(new_n656), .A2(new_n400), .ZN(new_n657));
  NOR2_X1   g296(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g297(.A(new_n658), .ZN(new_n659));
  AOI211_X1 g298(.A(new_n652), .B(new_n653), .C1(new_n659), .C2(G29), .ZN(new_n660));
  INV_X1    g299(.A(G2067), .ZN(new_n661));
  XNOR2_X1  g300(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g301(.A(G1966), .ZN(new_n663));
  AOI21_X1  g302(.A(new_n662), .B1(new_n663), .B2(new_n648), .ZN(new_n664));
  AOI21_X1  g303(.A(KEYINPUT23), .B1(new_n569), .B2(G20), .ZN(new_n665));
  AND3_X1   g304(.A1(new_n569), .A2(KEYINPUT23), .A3(G20), .ZN(new_n666));
  AOI211_X1 g305(.A(new_n665), .B(new_n666), .C1(G299), .C2(G16), .ZN(new_n667));
  XNOR2_X1  g306(.A(new_n667), .B(G1956), .ZN(new_n668));
  NAND2_X1  g307(.A1(new_n589), .A2(G35), .ZN(new_n669));
  OAI21_X1  g308(.A(new_n669), .B1(G162), .B2(new_n589), .ZN(new_n670));
  XOR2_X1   g309(.A(KEYINPUT29), .B(G2090), .Z(new_n671));
  XNOR2_X1  g310(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND3_X1  g311(.A1(new_n664), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NOR4_X1   g312(.A1(new_n635), .A2(new_n638), .A3(new_n651), .A4(new_n673), .ZN(new_n674));
  AND3_X1   g313(.A1(new_n598), .A2(new_n610), .A3(new_n674), .ZN(G311));
  NAND3_X1  g314(.A1(new_n598), .A2(new_n610), .A3(new_n674), .ZN(G150));
  AOI22_X1  g315(.A1(new_n424), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n677));
  AOI22_X1  g316(.A1(new_n424), .A2(G93), .B1(G55), .B2(G543), .ZN(new_n678));
  OAI22_X1  g317(.A1(new_n431), .A2(new_n677), .B1(new_n678), .B2(new_n428), .ZN(new_n679));
  NAND2_X1  g318(.A1(new_n679), .A2(G860), .ZN(new_n680));
  XOR2_X1   g319(.A(new_n680), .B(KEYINPUT37), .Z(new_n681));
  NOR2_X1   g320(.A1(new_n497), .A2(new_n504), .ZN(new_n682));
  XNOR2_X1  g321(.A(new_n682), .B(new_n679), .ZN(new_n683));
  XNOR2_X1  g322(.A(new_n683), .B(KEYINPUT39), .ZN(new_n684));
  XNOR2_X1  g323(.A(new_n457), .B(KEYINPUT38), .ZN(new_n685));
  XNOR2_X1  g324(.A(new_n684), .B(new_n685), .ZN(new_n686));
  OAI21_X1  g325(.A(new_n681), .B1(new_n686), .B2(G860), .ZN(G145));
  AOI22_X1  g326(.A1(new_n409), .A2(G130), .B1(G118), .B2(G2104), .ZN(new_n688));
  AOI22_X1  g327(.A1(new_n409), .A2(G142), .B1(G106), .B2(G2104), .ZN(new_n689));
  MUX2_X1   g328(.A(new_n688), .B(new_n689), .S(new_n400), .Z(new_n690));
  XOR2_X1   g329(.A(new_n593), .B(new_n690), .Z(new_n691));
  XNOR2_X1  g330(.A(new_n691), .B(new_n606), .ZN(new_n692));
  XNOR2_X1  g331(.A(G160), .B(G162), .ZN(new_n693));
  INV_X1    g332(.A(new_n517), .ZN(new_n694));
  NAND2_X1  g333(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g334(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g335(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  OAI21_X1  g336(.A(new_n514), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g337(.A(new_n697), .ZN(new_n699));
  INV_X1    g338(.A(new_n514), .ZN(new_n700));
  NAND3_X1  g339(.A1(new_n699), .A2(new_n700), .A3(new_n695), .ZN(new_n701));
  AOI21_X1  g340(.A(new_n692), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  INV_X1    g341(.A(new_n702), .ZN(new_n703));
  AND3_X1   g342(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n704));
  AOI21_X1  g343(.A(new_n419), .B1(new_n418), .B2(G138), .ZN(new_n705));
  NOR2_X1   g344(.A1(new_n421), .A2(KEYINPUT4), .ZN(new_n706));
  OAI21_X1  g345(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g346(.A(new_n631), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g347(.A(new_n708), .B(new_n659), .ZN(new_n709));
  NAND3_X1  g348(.A1(new_n698), .A2(new_n701), .A3(new_n692), .ZN(new_n710));
  NAND3_X1  g349(.A1(new_n703), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g350(.A(new_n709), .ZN(new_n712));
  INV_X1    g351(.A(new_n710), .ZN(new_n713));
  OAI21_X1  g352(.A(new_n712), .B1(new_n713), .B2(new_n702), .ZN(new_n714));
  INV_X1    g353(.A(G37), .ZN(new_n715));
  NAND3_X1  g354(.A1(new_n711), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g355(.A(new_n716), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g356(.A1(new_n679), .A2(G868), .ZN(new_n718));
  XOR2_X1   g357(.A(new_n457), .B(new_n679), .Z(new_n719));
  XNOR2_X1  g358(.A(new_n719), .B(new_n506), .ZN(new_n720));
  NAND2_X1  g359(.A1(new_n498), .A2(new_n475), .ZN(new_n721));
  NAND2_X1  g360(.A1(G299), .A2(new_n497), .ZN(new_n722));
  NAND2_X1  g361(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g362(.A(KEYINPUT41), .ZN(new_n724));
  NAND2_X1  g363(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g364(.A(new_n497), .B(new_n475), .ZN(new_n726));
  NAND2_X1  g365(.A1(new_n726), .A2(KEYINPUT41), .ZN(new_n727));
  NAND2_X1  g366(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g367(.A1(new_n720), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g368(.A(new_n457), .B(new_n679), .ZN(new_n730));
  XNOR2_X1  g369(.A(new_n730), .B(new_n506), .ZN(new_n731));
  NAND2_X1  g370(.A1(new_n731), .A2(new_n723), .ZN(new_n732));
  NAND2_X1  g371(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g372(.A1(new_n733), .A2(KEYINPUT42), .ZN(new_n734));
  INV_X1    g373(.A(KEYINPUT42), .ZN(new_n735));
  NAND3_X1  g374(.A1(new_n729), .A2(new_n735), .A3(new_n732), .ZN(new_n736));
  NAND2_X1  g375(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g376(.A(G290), .B(G305), .ZN(new_n738));
  OR2_X1    g377(.A1(new_n738), .A2(G303), .ZN(new_n739));
  NAND2_X1  g378(.A1(new_n738), .A2(G303), .ZN(new_n740));
  NAND2_X1  g379(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g380(.A1(new_n741), .A2(G288), .ZN(new_n742));
  NAND3_X1  g381(.A1(new_n739), .A2(new_n574), .A3(new_n740), .ZN(new_n743));
  AND2_X1   g382(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g383(.A(new_n737), .B(new_n744), .ZN(new_n745));
  AOI21_X1  g384(.A(new_n718), .B1(new_n745), .B2(G868), .ZN(G295));
  AOI21_X1  g385(.A(new_n718), .B1(new_n745), .B2(G868), .ZN(G331));
  XOR2_X1   g386(.A(G171), .B(G286), .Z(new_n748));
  XNOR2_X1  g387(.A(new_n730), .B(new_n748), .ZN(new_n749));
  NAND3_X1  g388(.A1(new_n749), .A2(new_n725), .A3(new_n727), .ZN(new_n750));
  AND2_X1   g389(.A1(new_n719), .A2(new_n748), .ZN(new_n751));
  NOR2_X1   g390(.A1(new_n719), .A2(new_n748), .ZN(new_n752));
  OAI21_X1  g391(.A(new_n726), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g392(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g393(.A1(new_n754), .A2(new_n744), .ZN(new_n755));
  NAND2_X1  g394(.A1(new_n742), .A2(new_n743), .ZN(new_n756));
  NAND3_X1  g395(.A1(new_n756), .A2(new_n750), .A3(new_n753), .ZN(new_n757));
  NAND3_X1  g396(.A1(new_n755), .A2(new_n715), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g397(.A1(new_n758), .A2(KEYINPUT43), .ZN(new_n759));
  INV_X1    g398(.A(KEYINPUT43), .ZN(new_n760));
  NAND4_X1  g399(.A1(new_n755), .A2(new_n760), .A3(new_n715), .A4(new_n757), .ZN(new_n761));
  NAND2_X1  g400(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g401(.A(KEYINPUT44), .ZN(new_n763));
  NAND2_X1  g402(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g403(.A1(new_n759), .A2(KEYINPUT44), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g404(.A1(new_n764), .A2(new_n765), .ZN(G397));
  AND3_X1   g405(.A1(new_n401), .A2(new_n405), .A3(G40), .ZN(new_n767));
  INV_X1    g406(.A(KEYINPUT45), .ZN(new_n768));
  OAI211_X1 g407(.A(new_n767), .B(new_n768), .C1(G1384), .C2(G164), .ZN(new_n769));
  INV_X1    g408(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g409(.A1(new_n659), .A2(G2067), .ZN(new_n771));
  NOR2_X1   g410(.A1(new_n658), .A2(new_n661), .ZN(new_n772));
  OAI21_X1  g411(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g412(.A1(new_n769), .A2(new_n606), .ZN(new_n774));
  NOR2_X1   g413(.A1(new_n769), .A2(G1996), .ZN(new_n775));
  NOR2_X1   g414(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g415(.A(new_n776), .B1(new_n605), .B2(new_n775), .ZN(new_n777));
  NAND3_X1  g416(.A1(new_n401), .A2(new_n405), .A3(G40), .ZN(new_n778));
  INV_X1    g417(.A(G1384), .ZN(new_n779));
  AOI211_X1 g418(.A(KEYINPUT45), .B(new_n778), .C1(new_n779), .C2(new_n707), .ZN(new_n780));
  NAND2_X1  g419(.A1(new_n780), .A2(new_n595), .ZN(new_n781));
  OR2_X1    g420(.A1(new_n769), .A2(new_n593), .ZN(new_n782));
  XNOR2_X1  g421(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g422(.A1(G290), .A2(G1986), .ZN(new_n784));
  NAND2_X1  g423(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  INV_X1    g424(.A(new_n785), .ZN(new_n786));
  OR2_X1    g425(.A1(new_n786), .A2(KEYINPUT48), .ZN(new_n787));
  NAND2_X1  g426(.A1(new_n786), .A2(KEYINPUT48), .ZN(new_n788));
  NAND3_X1  g427(.A1(new_n783), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g428(.A1(new_n782), .A2(new_n595), .A3(new_n780), .ZN(new_n790));
  AOI21_X1  g429(.A(new_n777), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g430(.A(new_n775), .B(KEYINPUT46), .ZN(new_n792));
  INV_X1    g431(.A(KEYINPUT47), .ZN(new_n793));
  NOR3_X1   g432(.A1(new_n792), .A2(new_n793), .A3(new_n774), .ZN(new_n794));
  OAI21_X1  g433(.A(new_n773), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g434(.A(new_n773), .B1(new_n606), .B2(new_n769), .ZN(new_n796));
  OAI21_X1  g435(.A(new_n793), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g436(.A1(new_n780), .A2(new_n771), .ZN(new_n798));
  AND3_X1   g437(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g438(.A1(new_n767), .A2(new_n779), .A3(new_n707), .ZN(new_n800));
  NAND2_X1  g439(.A1(new_n800), .A2(G8), .ZN(new_n801));
  XNOR2_X1  g440(.A(KEYINPUT49), .B(G1981), .ZN(new_n802));
  XNOR2_X1  g441(.A(G305), .B(new_n802), .ZN(new_n803));
  NOR4_X1   g442(.A1(new_n801), .A2(new_n803), .A3(G1976), .A4(G288), .ZN(new_n804));
  NOR3_X1   g443(.A1(new_n801), .A2(G1981), .A3(G305), .ZN(new_n805));
  NOR2_X1   g444(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR3_X1    g445(.A1(new_n801), .A2(G1976), .A3(new_n574), .ZN(new_n807));
  INV_X1    g446(.A(new_n801), .ZN(new_n808));
  NAND2_X1  g447(.A1(new_n574), .A2(G1976), .ZN(new_n809));
  NAND3_X1  g448(.A1(new_n808), .A2(KEYINPUT52), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g449(.A1(new_n809), .A2(new_n800), .A3(G8), .ZN(new_n811));
  INV_X1    g450(.A(KEYINPUT52), .ZN(new_n812));
  NAND2_X1  g451(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g452(.A1(new_n807), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g453(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n815));
  INV_X1    g454(.A(KEYINPUT50), .ZN(new_n816));
  NAND3_X1  g455(.A1(new_n707), .A2(new_n816), .A3(new_n779), .ZN(new_n817));
  NAND4_X1  g456(.A1(new_n815), .A2(new_n817), .A3(new_n644), .A4(new_n767), .ZN(new_n818));
  OAI21_X1  g457(.A(KEYINPUT45), .B1(G164), .B2(G1384), .ZN(new_n819));
  NAND3_X1  g458(.A1(new_n707), .A2(new_n768), .A3(new_n779), .ZN(new_n820));
  AOI21_X1  g459(.A(new_n778), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g460(.A(new_n818), .B1(new_n821), .B2(G1966), .ZN(new_n822));
  NAND4_X1  g461(.A1(new_n814), .A2(G8), .A3(G168), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g462(.A1(G303), .A2(G8), .ZN(new_n824));
  XNOR2_X1  g463(.A(new_n824), .B(KEYINPUT55), .ZN(new_n825));
  INV_X1    g464(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g465(.A1(new_n815), .A2(new_n817), .A3(new_n767), .ZN(new_n827));
  OAI22_X1  g466(.A1(new_n821), .A2(G1971), .B1(new_n827), .B2(G2090), .ZN(new_n828));
  NAND3_X1  g467(.A1(new_n826), .A2(G8), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g468(.A1(new_n828), .A2(G8), .ZN(new_n830));
  NAND2_X1  g469(.A1(new_n830), .A2(new_n825), .ZN(new_n831));
  NAND2_X1  g470(.A1(new_n808), .A2(new_n803), .ZN(new_n832));
  NAND3_X1  g471(.A1(new_n829), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g472(.A1(new_n823), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g473(.A1(new_n834), .A2(KEYINPUT63), .ZN(new_n835));
  INV_X1    g474(.A(KEYINPUT63), .ZN(new_n836));
  NOR3_X1   g475(.A1(new_n823), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g476(.A(new_n806), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g477(.A1(new_n821), .A2(new_n614), .ZN(new_n839));
  INV_X1    g478(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g479(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g480(.A(G1961), .ZN(new_n842));
  NAND2_X1  g481(.A1(new_n827), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g482(.A1(new_n821), .A2(KEYINPUT53), .A3(new_n614), .ZN(new_n844));
  NAND3_X1  g483(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AND3_X1   g484(.A1(new_n829), .A2(new_n831), .A3(new_n845), .ZN(new_n846));
  OAI211_X1 g485(.A(G168), .B(new_n818), .C1(new_n821), .C2(G1966), .ZN(new_n847));
  NAND2_X1  g486(.A1(new_n847), .A2(G8), .ZN(new_n848));
  INV_X1    g487(.A(KEYINPUT51), .ZN(new_n849));
  NAND2_X1  g488(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g489(.A1(new_n847), .A2(KEYINPUT51), .A3(G8), .ZN(new_n851));
  NAND2_X1  g490(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g491(.A1(new_n822), .A2(G8), .A3(G286), .ZN(new_n853));
  AOI21_X1  g492(.A(KEYINPUT62), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g493(.A1(new_n847), .A2(KEYINPUT51), .A3(G8), .ZN(new_n855));
  AOI21_X1  g494(.A(KEYINPUT51), .B1(new_n847), .B2(G8), .ZN(new_n856));
  OAI211_X1 g495(.A(KEYINPUT62), .B(new_n853), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  INV_X1    g496(.A(new_n857), .ZN(new_n858));
  OAI211_X1 g497(.A(G171), .B(new_n846), .C1(new_n854), .C2(new_n858), .ZN(new_n859));
  INV_X1    g498(.A(KEYINPUT61), .ZN(new_n860));
  XNOR2_X1  g499(.A(KEYINPUT56), .B(G2072), .ZN(new_n861));
  INV_X1    g500(.A(G1956), .ZN(new_n862));
  AOI22_X1  g501(.A1(new_n821), .A2(new_n861), .B1(new_n827), .B2(new_n862), .ZN(new_n863));
  INV_X1    g502(.A(new_n474), .ZN(new_n864));
  INV_X1    g503(.A(KEYINPUT57), .ZN(new_n865));
  OAI211_X1 g504(.A(new_n864), .B(new_n865), .C1(new_n469), .C2(new_n468), .ZN(new_n866));
  OAI21_X1  g505(.A(KEYINPUT57), .B1(new_n470), .B2(new_n474), .ZN(new_n867));
  AND2_X1   g506(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g507(.A(new_n860), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g508(.A1(new_n821), .A2(new_n861), .ZN(new_n870));
  NAND2_X1  g509(.A1(new_n827), .A2(new_n862), .ZN(new_n871));
  AND4_X1   g510(.A1(new_n860), .A2(new_n870), .A3(new_n868), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g511(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  AOI211_X1 g512(.A(G1996), .B(new_n778), .C1(new_n819), .C2(new_n820), .ZN(new_n874));
  NOR3_X1   g513(.A1(new_n778), .A2(G1384), .A3(G164), .ZN(new_n875));
  XOR2_X1   g514(.A(KEYINPUT58), .B(G1341), .Z(new_n876));
  INV_X1    g515(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g516(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g517(.A(new_n458), .B1(new_n874), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g518(.A1(new_n879), .A2(KEYINPUT59), .ZN(new_n880));
  INV_X1    g519(.A(KEYINPUT59), .ZN(new_n881));
  OAI211_X1 g520(.A(new_n881), .B(new_n458), .C1(new_n874), .C2(new_n878), .ZN(new_n882));
  NAND2_X1  g521(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g522(.A1(new_n827), .A2(new_n613), .ZN(new_n884));
  NAND2_X1  g523(.A1(new_n875), .A2(new_n661), .ZN(new_n885));
  AND3_X1   g524(.A1(new_n884), .A2(new_n497), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g525(.A(new_n497), .B1(new_n884), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g526(.A(KEYINPUT60), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g527(.A1(new_n497), .A2(KEYINPUT60), .ZN(new_n889));
  NAND3_X1  g528(.A1(new_n884), .A2(new_n889), .A3(new_n885), .ZN(new_n890));
  NAND4_X1  g529(.A1(new_n873), .A2(new_n883), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  INV_X1    g530(.A(new_n863), .ZN(new_n892));
  INV_X1    g531(.A(new_n868), .ZN(new_n893));
  OAI21_X1  g532(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g533(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  AND3_X1   g534(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g535(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n897));
  INV_X1    g536(.A(KEYINPUT54), .ZN(new_n898));
  NAND4_X1  g537(.A1(new_n841), .A2(new_n898), .A3(new_n843), .A4(new_n844), .ZN(new_n899));
  NAND2_X1  g538(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g539(.A1(new_n900), .A2(G301), .ZN(new_n901));
  AND2_X1   g540(.A1(new_n829), .A2(new_n831), .ZN(new_n902));
  NAND2_X1  g541(.A1(new_n852), .A2(new_n853), .ZN(new_n903));
  NAND3_X1  g542(.A1(new_n897), .A2(G171), .A3(new_n899), .ZN(new_n904));
  NAND4_X1  g543(.A1(new_n901), .A2(new_n902), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  OAI211_X1 g544(.A(new_n859), .B(new_n829), .C1(new_n896), .C2(new_n905), .ZN(new_n906));
  AND2_X1   g545(.A1(new_n814), .A2(new_n832), .ZN(new_n907));
  AOI21_X1  g546(.A(new_n838), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g547(.A(new_n777), .ZN(new_n909));
  NOR2_X1   g548(.A1(new_n584), .A2(new_n586), .ZN(new_n910));
  OAI21_X1  g549(.A(new_n770), .B1(new_n784), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g550(.A1(new_n909), .A2(new_n783), .A3(new_n773), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g551(.A(new_n799), .B1(new_n908), .B2(new_n912), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g552(.A1(new_n716), .A2(G319), .ZN(new_n915));
  NOR2_X1   g553(.A1(G229), .A2(G401), .ZN(new_n916));
  AND4_X1   g554(.A1(new_n546), .A2(new_n762), .A3(new_n915), .A4(new_n916), .ZN(G308));
  NAND4_X1  g555(.A1(new_n762), .A2(new_n915), .A3(new_n546), .A4(new_n916), .ZN(G225));
endmodule


