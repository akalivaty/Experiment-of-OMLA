//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n187), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(KEYINPUT75), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT75), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n199), .A3(new_n195), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NOR2_X1   g015(.A1(G237), .A2(G953), .ZN(new_n202));
  AOI21_X1  g016(.A(G143), .B1(new_n202), .B2(G214), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(G143), .A3(G214), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT17), .A3(G131), .ZN(new_n207));
  INV_X1    g021(.A(new_n205), .ZN(new_n208));
  OAI21_X1  g022(.A(G131), .B1(new_n208), .B2(new_n203), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n210), .A3(new_n205), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n201), .A2(new_n207), .A3(new_n213), .ZN(new_n214));
  XOR2_X1   g028(.A(G113), .B(G122), .Z(new_n215));
  XOR2_X1   g029(.A(KEYINPUT92), .B(G104), .Z(new_n216));
  XOR2_X1   g030(.A(new_n215), .B(new_n216), .Z(new_n217));
  NAND3_X1  g031(.A1(new_n206), .A2(KEYINPUT18), .A3(G131), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n193), .A2(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n190), .A2(new_n192), .A3(new_n195), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT18), .A2(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n204), .A2(new_n205), .A3(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n218), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n217), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT93), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n213), .A2(new_n207), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n229), .B2(new_n201), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT93), .B1(new_n230), .B2(new_n217), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n193), .B(KEYINPUT19), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n197), .B1(new_n232), .B2(G146), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT91), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n209), .A2(new_n211), .ZN(new_n236));
  OAI211_X1 g050(.A(KEYINPUT91), .B(new_n197), .C1(new_n232), .C2(G146), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n238), .A2(new_n225), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n228), .A2(new_n231), .B1(new_n217), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n241));
  NOR2_X1   g055(.A1(G475), .A2(G902), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n217), .B1(new_n238), .B2(new_n225), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n226), .A2(new_n227), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n230), .A2(KEYINPUT93), .A3(new_n217), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n242), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT20), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G952), .ZN(new_n251));
  AOI211_X1 g065(.A(G953), .B(new_n251), .C1(G234), .C2(G237), .ZN(new_n252));
  NAND2_X1  g066(.A1(G234), .A2(G237), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(G902), .A3(G953), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n254), .B(KEYINPUT96), .Z(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT21), .B(G898), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G478), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT15), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G116), .B(G122), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT14), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G116), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(KEYINPUT14), .A3(G122), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(G107), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT95), .ZN(new_n268));
  INV_X1    g082(.A(G107), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G143), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G128), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G143), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n275), .A2(new_n276), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n270), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n268), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT13), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n274), .B1(new_n272), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT13), .B1(new_n271), .B2(G128), .ZN(new_n285));
  OAI21_X1  g099(.A(G134), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(KEYINPUT94), .ZN(new_n287));
  INV_X1    g101(.A(new_n270), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n262), .A2(new_n269), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n277), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT9), .B(G234), .ZN(new_n293));
  INV_X1    g107(.A(G217), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(new_n294), .A3(G953), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n295), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n281), .B2(new_n291), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n261), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  AOI211_X1 g115(.A(G902), .B(new_n260), .C1(new_n296), .C2(new_n298), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n230), .A2(new_n217), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(new_n245), .B2(new_n246), .ZN(new_n305));
  OAI21_X1  g119(.A(G475), .B1(new_n305), .B2(G902), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n250), .A2(new_n258), .A3(new_n303), .A4(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT97), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n228), .A2(new_n231), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n300), .B1(new_n309), .B2(new_n304), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n243), .A2(new_n249), .B1(new_n310), .B2(G475), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT97), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n311), .A2(new_n312), .A3(new_n258), .A4(new_n303), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n308), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT64), .B1(new_n276), .B2(G137), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT11), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT11), .ZN(new_n317));
  OAI211_X1 g131(.A(KEYINPUT64), .B(new_n317), .C1(new_n276), .C2(G137), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n276), .A2(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(KEYINPUT65), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n315), .A2(KEYINPUT11), .B1(new_n276), .B2(G137), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n318), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n195), .A2(G143), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n271), .A2(G146), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n329), .A2(KEYINPUT1), .A3(new_n273), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n329), .A2(new_n273), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n271), .A2(KEYINPUT1), .A3(G146), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(G128), .B1(new_n327), .B2(new_n328), .ZN(new_n336));
  INV_X1    g150(.A(new_n334), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n336), .A2(KEYINPUT67), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n331), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT10), .ZN(new_n340));
  OR2_X1    g154(.A1(KEYINPUT79), .A2(G104), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT79), .A2(G104), .ZN(new_n342));
  AOI21_X1  g156(.A(G107), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n269), .A2(G104), .ZN(new_n344));
  OAI21_X1  g158(.A(G101), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT82), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(G101), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n350));
  AND2_X1   g164(.A1(KEYINPUT79), .A2(G104), .ZN(new_n351));
  NOR2_X1   g165(.A1(KEYINPUT79), .A2(G104), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n269), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n269), .A3(G104), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT80), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n357), .A2(new_n354), .A3(new_n269), .A4(G104), .ZN(new_n358));
  AOI22_X1  g172(.A1(KEYINPUT3), .A2(new_n353), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n351), .A2(new_n352), .ZN(new_n360));
  AOI21_X1  g174(.A(G101), .B1(new_n360), .B2(G107), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n350), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n353), .A2(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n358), .ZN(new_n364));
  AND4_X1   g178(.A1(new_n350), .A2(new_n361), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n349), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT81), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n359), .A2(new_n350), .A3(new_n361), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT83), .A3(new_n349), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n340), .B1(new_n368), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n360), .A2(G107), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n359), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n377), .B2(G101), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n372), .ZN(new_n379));
  OR2_X1    g193(.A1(KEYINPUT0), .A2(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT0), .A2(G128), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n327), .A2(new_n328), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n327), .A2(new_n328), .A3(new_n381), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G101), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n359), .B2(new_n376), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n386), .B2(new_n375), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n331), .A2(new_n333), .A3(new_n334), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n349), .B(new_n389), .C1(new_n362), .C2(new_n365), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT10), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n326), .B1(new_n374), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g208(.A1(new_n379), .A2(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n395));
  INV_X1    g209(.A(new_n326), .ZN(new_n396));
  AOI221_X4 g210(.A(new_n367), .B1(new_n346), .B2(new_n348), .C1(new_n370), .C2(new_n371), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT83), .B1(new_n372), .B2(new_n349), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n395), .B(new_n396), .C1(new_n399), .C2(new_n340), .ZN(new_n400));
  XNOR2_X1  g214(.A(G110), .B(G140), .ZN(new_n401));
  INV_X1    g215(.A(G227), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(G953), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n401), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n394), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT67), .B1(new_n336), .B2(new_n337), .ZN(new_n407));
  XNOR2_X1  g221(.A(G143), .B(G146), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n334), .B(new_n332), .C1(new_n408), .C2(G128), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n330), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n368), .A2(new_n410), .A3(new_n373), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n390), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT12), .B1(new_n412), .B2(new_n326), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT12), .ZN(new_n414));
  AOI211_X1 g228(.A(new_n414), .B(new_n396), .C1(new_n411), .C2(new_n390), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n400), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n406), .B1(new_n416), .B2(new_n404), .ZN(new_n417));
  OAI21_X1  g231(.A(G469), .B1(new_n417), .B2(G902), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n400), .B(new_n405), .C1(new_n413), .C2(new_n415), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n394), .A2(new_n400), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n404), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT84), .B(G469), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n314), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  INV_X1    g243(.A(G953), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n429), .A2(new_n430), .A3(G210), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n428), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT26), .B(G101), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n432), .B(new_n433), .Z(new_n434));
  OR2_X1    g248(.A1(new_n382), .A2(new_n383), .ZN(new_n435));
  AND4_X1   g249(.A1(new_n318), .A2(new_n316), .A3(new_n319), .A4(new_n321), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n321), .B1(new_n324), .B2(new_n318), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G116), .B(G119), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(KEYINPUT69), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT2), .B(G113), .Z(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n316), .A2(new_n210), .A3(new_n318), .A4(new_n319), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n276), .B2(G137), .ZN(new_n445));
  INV_X1    g259(.A(G137), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT66), .A3(G134), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n319), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G131), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n438), .B(new_n442), .C1(new_n410), .C2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT28), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT68), .ZN(new_n453));
  INV_X1    g267(.A(new_n450), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n339), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT68), .B1(new_n410), .B2(new_n450), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n438), .ZN(new_n457));
  INV_X1    g271(.A(new_n442), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n434), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT31), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n407), .A2(new_n409), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n450), .B1(new_n462), .B2(new_n331), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n384), .B1(new_n323), .B2(new_n325), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n442), .B(new_n466), .C1(new_n465), .C2(new_n457), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n451), .A2(new_n434), .A3(KEYINPUT71), .ZN(new_n468));
  AOI21_X1  g282(.A(KEYINPUT71), .B1(new_n451), .B2(new_n434), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n461), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n451), .A2(new_n434), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT71), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n451), .A2(new_n434), .A3(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n457), .A2(new_n465), .ZN(new_n477));
  INV_X1    g291(.A(new_n466), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n458), .A3(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT31), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n460), .B1(new_n471), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(G472), .A2(G902), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT72), .Z(new_n483));
  OAI21_X1  g297(.A(KEYINPUT32), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n460), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT31), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT31), .B1(new_n476), .B2(new_n479), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT32), .ZN(new_n489));
  INV_X1    g303(.A(new_n483), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n484), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G472), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n452), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n434), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(G902), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n452), .A2(new_n459), .A3(new_n434), .ZN(new_n500));
  INV_X1    g314(.A(new_n451), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n466), .B1(new_n457), .B2(new_n465), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n458), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n500), .B(new_n497), .C1(new_n503), .C2(new_n434), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n493), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT73), .B1(new_n492), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT73), .ZN(new_n508));
  AOI211_X1 g322(.A(new_n508), .B(new_n505), .C1(new_n484), .C2(new_n491), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G214), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G113), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n265), .A2(G119), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n439), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n441), .A2(new_n439), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n368), .B2(new_n373), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n442), .B1(new_n375), .B2(new_n386), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n379), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT86), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n520), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n397), .B2(new_n398), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT86), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  XNOR2_X1  g343(.A(G110), .B(G122), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT87), .Z(new_n531));
  INV_X1    g345(.A(KEYINPUT6), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n525), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT88), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n525), .A2(new_n529), .A3(new_n536), .A4(new_n533), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n525), .A2(new_n529), .A3(new_n531), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n521), .A2(new_n524), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n532), .B1(new_n540), .B2(new_n530), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n384), .A2(G125), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT89), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n544), .B1(new_n191), .B2(new_n410), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n430), .A2(G224), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n538), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n540), .A2(new_n530), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n530), .B(KEYINPUT8), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT5), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n516), .B1(new_n551), .B2(new_n517), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n519), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n368), .B2(new_n373), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n526), .B1(new_n372), .B2(new_n349), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n546), .A2(KEYINPUT7), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n410), .A2(new_n191), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n543), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n545), .B2(new_n557), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n549), .A2(new_n556), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n300), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n548), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G210), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g383(.A1(new_n535), .A2(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n562), .B1(new_n570), .B2(new_n547), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n567), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n512), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n294), .B1(G234), .B2(new_n300), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n273), .A2(G119), .ZN(new_n577));
  INV_X1    g391(.A(G119), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G128), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT24), .B(G110), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n273), .A2(KEYINPUT23), .A3(G119), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n578), .A2(G128), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(new_n579), .C1(new_n584), .C2(KEYINPUT23), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n585), .B2(G110), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT76), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(new_n197), .A3(new_n220), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n580), .A2(new_n581), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n590), .A2(KEYINPUT74), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(KEYINPUT74), .ZN(new_n592));
  AOI22_X1  g406(.A1(new_n591), .A2(new_n592), .B1(G110), .B2(new_n585), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n200), .A3(new_n198), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT22), .B(G137), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n430), .A2(G221), .A3(G234), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n589), .A2(new_n594), .A3(new_n598), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n300), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n576), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n603), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n600), .A2(new_n300), .A3(new_n601), .A4(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n575), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n574), .A2(G902), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n600), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OR3_X1    g424(.A1(new_n607), .A2(KEYINPUT78), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT78), .B1(new_n607), .B2(new_n610), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n427), .A2(new_n510), .A3(new_n573), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  INV_X1    g429(.A(KEYINPUT98), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n511), .B1(new_n571), .B2(new_n566), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n565), .B(new_n562), .C1(new_n570), .C2(new_n547), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n512), .B1(new_n564), .B2(new_n565), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n571), .A2(new_n566), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(KEYINPUT98), .A3(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n311), .ZN(new_n623));
  AOI21_X1  g437(.A(G478), .B1(new_n299), .B2(new_n300), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n299), .A2(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n282), .A2(new_n292), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n297), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n296), .A2(new_n629), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n627), .B(KEYINPUT99), .C1(new_n629), .C2(new_n297), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n626), .B1(new_n634), .B2(KEYINPUT33), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n259), .A2(G902), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n625), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n623), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n619), .A2(new_n622), .A3(new_n258), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n611), .A2(new_n612), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n481), .A2(G902), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n493), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n481), .A2(new_n483), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n426), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n418), .B2(new_n424), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT34), .B(G104), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NOR3_X1   g466(.A1(new_n617), .A2(new_n616), .A3(new_n618), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT98), .B1(new_n620), .B2(new_n621), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n303), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n311), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n655), .A2(new_n258), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(new_n649), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n644), .A2(new_n645), .ZN(new_n663));
  INV_X1    g477(.A(new_n607), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n589), .A2(new_n594), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n665), .B1(new_n589), .B2(new_n594), .ZN(new_n668));
  OAI22_X1  g482(.A1(new_n667), .A2(new_n668), .B1(KEYINPUT36), .B2(new_n599), .ZN(new_n669));
  INV_X1    g483(.A(new_n668), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n599), .A2(KEYINPUT36), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n670), .A2(new_n671), .A3(new_n666), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n608), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT102), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT102), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n673), .A2(new_n676), .A3(new_n608), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n664), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n427), .A2(new_n573), .A3(new_n663), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT37), .B(G110), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G12));
  NOR3_X1   g495(.A1(new_n481), .A2(KEYINPUT32), .A3(new_n483), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n506), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n508), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n492), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n686));
  AND4_X1   g500(.A1(new_n685), .A2(new_n648), .A3(new_n686), .A4(new_n678), .ZN(new_n687));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n252), .B1(new_n255), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n657), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n687), .A2(new_n619), .A3(new_n622), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  XOR2_X1   g506(.A(new_n689), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n648), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT40), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n569), .A2(new_n572), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n434), .B1(new_n494), .B2(new_n451), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n476), .B2(new_n479), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n492), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n311), .A2(new_n303), .ZN(new_n703));
  INV_X1    g517(.A(new_n678), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n511), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n695), .A2(new_n698), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT104), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G143), .ZN(G45));
  INV_X1    g522(.A(new_n689), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n623), .A2(new_n638), .A3(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n687), .A2(new_n619), .A3(new_n622), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NAND3_X1  g527(.A1(new_n685), .A2(new_n613), .A3(new_n686), .ZN(new_n714));
  INV_X1    g528(.A(G469), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n424), .B(new_n426), .C1(new_n422), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n655), .A2(new_n258), .A3(new_n640), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND4_X1  g534(.A1(new_n655), .A2(new_n258), .A3(new_n658), .A4(new_n717), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n723));
  INV_X1    g537(.A(new_n716), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n619), .A2(new_n622), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n510), .A2(new_n314), .A3(new_n678), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n723), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n619), .A2(new_n622), .A3(new_n724), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n726), .A3(KEYINPUT105), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n578), .ZN(G21));
  NOR2_X1   g546(.A1(new_n607), .A2(new_n610), .ZN(new_n733));
  OAI22_X1  g547(.A1(new_n486), .A2(new_n487), .B1(new_n434), .B2(new_n495), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n490), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n733), .B(new_n735), .C1(new_n643), .C2(new_n493), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n716), .A2(new_n736), .A3(new_n257), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n619), .A3(new_n622), .A4(new_n703), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  OAI211_X1 g553(.A(new_n678), .B(new_n735), .C1(new_n493), .C2(new_n643), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n710), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n619), .A2(new_n622), .A3(new_n724), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  INV_X1    g557(.A(new_n696), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n505), .B1(new_n484), .B2(new_n491), .ZN(new_n745));
  INV_X1    g559(.A(new_n733), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n710), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n744), .A2(new_n747), .A3(new_n511), .A4(new_n648), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n648), .A2(new_n511), .A3(new_n569), .A4(new_n572), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n714), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n751));
  AOI22_X1  g565(.A1(KEYINPUT42), .A2(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G131), .ZN(G33));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n690), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n638), .A2(new_n311), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT43), .Z(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT106), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT106), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  AOI211_X1 g574(.A(new_n704), .B(new_n663), .C1(KEYINPUT107), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(KEYINPUT107), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(G469), .B1(new_n417), .B2(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(KEYINPUT45), .B2(new_n417), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n715), .A2(new_n300), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n424), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n771), .B1(new_n768), .B2(new_n769), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n647), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n569), .A2(new_n572), .A3(new_n511), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT108), .Z(new_n775));
  NAND4_X1  g589(.A1(new_n764), .A2(new_n693), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G137), .ZN(G39));
  XOR2_X1   g591(.A(new_n773), .B(KEYINPUT47), .Z(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n774), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n510), .A2(new_n613), .A3(new_n710), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  AND2_X1   g597(.A1(new_n757), .A2(new_n252), .ZN(new_n784));
  INV_X1    g598(.A(new_n736), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n251), .B(G953), .C1(new_n786), .C2(new_n725), .ZN(new_n787));
  INV_X1    g601(.A(new_n702), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n613), .A3(new_n252), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n789), .A2(new_n774), .A3(new_n716), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT116), .Z(new_n791));
  NAND3_X1  g605(.A1(new_n784), .A2(new_n724), .A3(new_n780), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n792), .A2(new_n745), .A3(new_n746), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT48), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT118), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n794), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT117), .ZN(new_n798));
  OAI221_X1 g612(.A(new_n787), .B1(new_n639), .B2(new_n791), .C1(new_n796), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT119), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n786), .A2(new_n512), .A3(new_n698), .A4(new_n724), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT50), .Z(new_n802));
  OR3_X1    g616(.A1(new_n791), .A2(new_n623), .A3(new_n638), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n802), .B(new_n803), .C1(new_n740), .C2(new_n792), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n786), .A2(new_n775), .ZN(new_n806));
  INV_X1    g620(.A(new_n422), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n771), .B1(G469), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n647), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n806), .B1(new_n778), .B2(new_n809), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n804), .A2(new_n805), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n809), .B(KEYINPUT115), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n806), .B1(new_n778), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n805), .B1(new_n804), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n800), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT111), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n648), .A2(new_n704), .A3(new_n709), .A4(new_n702), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(new_n619), .A3(new_n622), .A4(new_n703), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n691), .A2(new_n712), .A3(new_n742), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n816), .B1(new_n819), .B2(KEYINPUT52), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n691), .A2(new_n712), .A3(new_n818), .A4(new_n742), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n821), .A2(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT112), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT111), .B1(new_n821), .B2(new_n823), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n780), .A2(new_n648), .A3(new_n741), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n623), .A2(new_n656), .A3(new_n689), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n744), .A2(KEYINPUT110), .A3(new_n511), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  INV_X1    g650(.A(new_n834), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n836), .B1(new_n774), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n838), .A3(new_n687), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n752), .A2(new_n754), .A3(new_n833), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n257), .B1(new_n639), .B2(new_n657), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n573), .A2(new_n646), .A3(new_n648), .A4(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n614), .A2(new_n679), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n718), .A3(new_n721), .A4(new_n738), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n840), .A2(new_n844), .A3(new_n731), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n826), .A2(new_n831), .A3(new_n832), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n691), .A2(new_n742), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n712), .A2(new_n818), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT52), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n827), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n844), .A2(new_n731), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n748), .A2(KEYINPUT42), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n750), .A2(new_n751), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n754), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n839), .A2(new_n833), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT53), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n846), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n857), .B2(new_n832), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n826), .A2(new_n831), .A3(KEYINPUT53), .A4(new_n845), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n730), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT105), .B1(new_n729), .B2(new_n726), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n641), .A2(new_n714), .A3(new_n716), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n738), .A2(new_n614), .A3(new_n679), .A4(new_n842), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n856), .A2(new_n721), .A3(new_n868), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n828), .A2(new_n830), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n820), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n862), .A3(KEYINPUT53), .A4(new_n831), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT54), .B1(new_n865), .B2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT114), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n861), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n865), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n860), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT114), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n815), .A2(new_n882), .B1(G952), .B2(G953), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n756), .A2(new_n746), .A3(new_n512), .A4(new_n647), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT109), .Z(new_n885));
  XNOR2_X1  g699(.A(new_n808), .B(KEYINPUT49), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n698), .A3(new_n788), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(G75));
  NOR2_X1   g702(.A1(new_n430), .A2(G952), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT121), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n865), .A2(new_n875), .A3(G210), .A4(G902), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n570), .B(new_n547), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n891), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n892), .A2(KEYINPUT120), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n892), .B2(KEYINPUT120), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n897), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT122), .ZN(G51));
  XNOR2_X1  g716(.A(new_n879), .B(new_n860), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n767), .B(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n419), .A2(new_n421), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n879), .A2(new_n300), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n766), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n889), .B1(new_n907), .B2(new_n909), .ZN(G54));
  NAND3_X1  g724(.A1(new_n908), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(new_n247), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n911), .A2(new_n247), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n913), .A3(new_n889), .ZN(G60));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n915));
  INV_X1    g729(.A(new_n635), .ZN(new_n916));
  NAND2_X1  g730(.A1(G478), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT59), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n916), .B1(new_n882), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n635), .A2(new_n918), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n879), .A2(new_n860), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(new_n876), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n890), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n915), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n891), .B1(new_n903), .B2(new_n921), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n918), .B1(new_n878), .B2(new_n881), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n926), .B(KEYINPUT123), .C1(new_n916), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n928), .ZN(G63));
  NAND2_X1  g743(.A1(new_n600), .A2(new_n601), .ZN(new_n930));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT60), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n879), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n932), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n865), .A2(new_n875), .A3(new_n673), .A4(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n890), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(KEYINPUT125), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n938), .B1(new_n939), .B2(new_n936), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT125), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n256), .B2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT126), .Z(new_n945));
  INV_X1    g759(.A(new_n851), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n946), .B2(new_n430), .ZN(new_n947));
  INV_X1    g761(.A(G898), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n570), .B1(new_n948), .B2(G953), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n947), .B(new_n949), .ZN(G69));
  AOI21_X1  g764(.A(new_n694), .B1(new_n639), .B2(new_n657), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n780), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n782), .B(new_n776), .C1(new_n714), .C2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n847), .A2(new_n712), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n707), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n953), .B1(new_n955), .B2(KEYINPUT62), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n956), .B(new_n430), .C1(KEYINPUT62), .C2(new_n955), .ZN(new_n957));
  NAND3_X1  g771(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n502), .B(new_n232), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n776), .A2(new_n752), .A3(new_n754), .ZN(new_n961));
  AND4_X1   g775(.A1(new_n684), .A2(new_n655), .A3(new_n733), .A4(new_n703), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n773), .A3(new_n693), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n961), .A2(new_n782), .A3(new_n954), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n430), .ZN(new_n965));
  INV_X1    g779(.A(new_n959), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n402), .A2(G900), .A3(G953), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n960), .A2(new_n968), .ZN(G72));
  OAI21_X1  g783(.A(new_n434), .B1(new_n467), .B2(new_n501), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n946), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n956), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  AOI21_X1  g789(.A(new_n970), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n964), .B2(new_n946), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n977), .A2(new_n496), .A3(new_n503), .ZN(new_n978));
  INV_X1    g792(.A(new_n975), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n503), .A2(new_n434), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n479), .B2(new_n476), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n859), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NOR4_X1   g796(.A1(new_n976), .A2(new_n978), .A3(new_n889), .A4(new_n982), .ZN(G57));
endmodule


