

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795;

  AND2_X1 U384 ( .A1(n525), .A2(n611), .ZN(n524) );
  XNOR2_X1 U385 ( .A(n363), .B(n518), .ZN(n773) );
  XNOR2_X1 U386 ( .A(n564), .B(n451), .ZN(n363) );
  INV_X4 U387 ( .A(G953), .ZN(n784) );
  NAND2_X1 U388 ( .A1(n399), .A2(n421), .ZN(n605) );
  NAND2_X2 U389 ( .A1(n404), .A2(n680), .ZN(n446) );
  XNOR2_X2 U390 ( .A(n499), .B(n607), .ZN(n610) );
  INV_X2 U391 ( .A(KEYINPUT67), .ZN(n447) );
  XOR2_X1 U392 ( .A(n371), .B(n560), .Z(n364) );
  XNOR2_X2 U393 ( .A(n781), .B(n506), .ZN(n601) );
  XNOR2_X2 U394 ( .A(n579), .B(n389), .ZN(n781) );
  NAND2_X1 U395 ( .A1(n430), .A2(n431), .ZN(n429) );
  NOR2_X1 U396 ( .A1(n705), .A2(n674), .ZN(n675) );
  NOR2_X1 U397 ( .A1(n386), .A2(n461), .ZN(n401) );
  XNOR2_X1 U398 ( .A(n402), .B(KEYINPUT32), .ZN(n791) );
  XNOR2_X1 U399 ( .A(n473), .B(n376), .ZN(n793) );
  AND2_X1 U400 ( .A1(n407), .A2(n718), .ZN(n621) );
  AND2_X1 U401 ( .A1(n459), .A2(n458), .ZN(n386) );
  XNOR2_X1 U402 ( .A(n489), .B(n408), .ZN(n407) );
  XNOR2_X1 U403 ( .A(n390), .B(KEYINPUT92), .ZN(n399) );
  XNOR2_X1 U404 ( .A(n500), .B(KEYINPUT110), .ZN(n656) );
  XNOR2_X1 U405 ( .A(n503), .B(n377), .ZN(n502) );
  NOR2_X1 U406 ( .A1(n632), .A2(n633), .ZN(n666) );
  OR2_X1 U407 ( .A1(n630), .A2(n450), .ZN(n719) );
  XNOR2_X1 U408 ( .A(n594), .B(n373), .ZN(n630) );
  XNOR2_X1 U409 ( .A(n755), .B(n754), .ZN(n756) );
  NAND2_X1 U410 ( .A1(n428), .A2(n675), .ZN(n427) );
  BUF_X1 U411 ( .A(n672), .Z(n488) );
  XNOR2_X2 U412 ( .A(n477), .B(KEYINPUT4), .ZN(n389) );
  XNOR2_X2 U413 ( .A(n466), .B(n551), .ZN(n672) );
  XNOR2_X2 U414 ( .A(n446), .B(KEYINPUT64), .ZN(n514) );
  NAND2_X1 U415 ( .A1(n415), .A2(KEYINPUT75), .ZN(n414) );
  NAND2_X1 U416 ( .A1(n417), .A2(n429), .ZN(n416) );
  NOR2_X1 U417 ( .A1(G237), .A2(G902), .ZN(n542) );
  XNOR2_X1 U418 ( .A(G902), .B(KEYINPUT15), .ZN(n678) );
  XNOR2_X1 U419 ( .A(n426), .B(G140), .ZN(n589) );
  INV_X1 U420 ( .A(G137), .ZN(n426) );
  NAND2_X1 U421 ( .A1(G953), .A2(G902), .ZN(n624) );
  XNOR2_X1 U422 ( .A(n578), .B(G134), .ZN(n579) );
  INV_X1 U423 ( .A(KEYINPUT73), .ZN(n522) );
  AND2_X1 U424 ( .A1(n438), .A2(n675), .ZN(n430) );
  NAND2_X1 U425 ( .A1(n486), .A2(KEYINPUT48), .ZN(n433) );
  INV_X1 U426 ( .A(KEYINPUT42), .ZN(n464) );
  INV_X1 U427 ( .A(n630), .ZN(n487) );
  NAND2_X1 U428 ( .A1(G234), .A2(G237), .ZN(n541) );
  XNOR2_X1 U429 ( .A(n566), .B(n490), .ZN(n612) );
  XNOR2_X1 U430 ( .A(n565), .B(n491), .ZN(n490) );
  INV_X1 U431 ( .A(G475), .ZN(n491) );
  XNOR2_X1 U432 ( .A(n596), .B(n475), .ZN(n474) );
  XNOR2_X1 U433 ( .A(G137), .B(KEYINPUT5), .ZN(n596) );
  XNOR2_X1 U434 ( .A(G113), .B(G116), .ZN(n475) );
  XNOR2_X1 U435 ( .A(n393), .B(n397), .ZN(n392) );
  INV_X1 U436 ( .A(KEYINPUT76), .ZN(n397) );
  XNOR2_X1 U437 ( .A(KEYINPUT24), .B(G128), .ZN(n393) );
  XNOR2_X1 U438 ( .A(n396), .B(n395), .ZN(n394) );
  XNOR2_X1 U439 ( .A(G119), .B(KEYINPUT93), .ZN(n396) );
  XNOR2_X1 U440 ( .A(G110), .B(KEYINPUT23), .ZN(n395) );
  XNOR2_X1 U441 ( .A(n508), .B(n507), .ZN(n592) );
  INV_X1 U442 ( .A(KEYINPUT8), .ZN(n507) );
  NAND2_X1 U443 ( .A1(n784), .A2(G234), .ZN(n508) );
  XNOR2_X1 U444 ( .A(n591), .B(n590), .ZN(n780) );
  NOR2_X1 U445 ( .A1(G953), .A2(G237), .ZN(n597) );
  XNOR2_X1 U446 ( .A(n558), .B(KEYINPUT10), .ZN(n591) );
  XNOR2_X1 U447 ( .A(n422), .B(KEYINPUT71), .ZN(n575) );
  XNOR2_X1 U448 ( .A(G110), .B(KEYINPUT72), .ZN(n422) );
  XNOR2_X1 U449 ( .A(n589), .B(n424), .ZN(n423) );
  XNOR2_X1 U450 ( .A(G104), .B(n425), .ZN(n424) );
  INV_X1 U451 ( .A(KEYINPUT77), .ZN(n425) );
  INV_X1 U452 ( .A(G107), .ZN(n495) );
  XNOR2_X1 U453 ( .A(n581), .B(n580), .ZN(n506) );
  INV_X1 U454 ( .A(G146), .ZN(n580) );
  INV_X1 U455 ( .A(KEYINPUT41), .ZN(n405) );
  NAND2_X1 U456 ( .A1(n715), .A2(n711), .ZN(n406) );
  XNOR2_X1 U457 ( .A(KEYINPUT34), .B(KEYINPUT79), .ZN(n604) );
  INV_X1 U458 ( .A(KEYINPUT22), .ZN(n408) );
  XNOR2_X1 U459 ( .A(n492), .B(KEYINPUT103), .ZN(n496) );
  XNOR2_X1 U460 ( .A(n513), .B(n510), .ZN(n761) );
  XNOR2_X1 U461 ( .A(n511), .B(n568), .ZN(n510) );
  XNOR2_X1 U462 ( .A(n567), .B(n571), .ZN(n513) );
  XOR2_X1 U463 ( .A(G122), .B(KEYINPUT7), .Z(n568) );
  NAND2_X1 U464 ( .A1(n440), .A2(n662), .ZN(n439) );
  XNOR2_X1 U465 ( .A(n441), .B(KEYINPUT96), .ZN(n440) );
  NAND2_X1 U466 ( .A1(n442), .A2(n443), .ZN(n441) );
  NOR2_X1 U467 ( .A1(n793), .A2(n454), .ZN(n453) );
  INV_X1 U468 ( .A(n658), .ZN(n432) );
  NOR2_X1 U469 ( .A1(n411), .A2(n410), .ZN(n409) );
  NAND2_X1 U470 ( .A1(n414), .A2(n677), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n509), .B(G107), .ZN(n569) );
  INV_X1 U472 ( .A(G116), .ZN(n509) );
  XNOR2_X1 U473 ( .A(G146), .B(G125), .ZN(n558) );
  XNOR2_X1 U474 ( .A(n366), .B(KEYINPUT91), .ZN(n482) );
  XOR2_X1 U475 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n547) );
  NAND2_X1 U476 ( .A1(n526), .A2(n545), .ZN(n480) );
  INV_X1 U477 ( .A(KEYINPUT65), .ZN(n484) );
  NAND2_X1 U478 ( .A1(n710), .A2(n721), .ZN(n492) );
  XNOR2_X1 U479 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U480 ( .A(n569), .B(n519), .ZN(n518) );
  INV_X1 U481 ( .A(KEYINPUT16), .ZN(n519) );
  XNOR2_X1 U482 ( .A(n570), .B(KEYINPUT9), .ZN(n512) );
  INV_X1 U483 ( .A(KEYINPUT99), .ZN(n570) );
  XNOR2_X1 U484 ( .A(n481), .B(n478), .ZN(n745) );
  NAND2_X1 U485 ( .A1(n480), .A2(n479), .ZN(n478) );
  XNOR2_X1 U486 ( .A(n773), .B(n482), .ZN(n481) );
  NAND2_X1 U487 ( .A1(n544), .A2(n543), .ZN(n479) );
  XOR2_X1 U488 ( .A(n603), .B(KEYINPUT33), .Z(n717) );
  XNOR2_X1 U489 ( .A(n676), .B(KEYINPUT87), .ZN(n403) );
  NAND2_X1 U490 ( .A1(n656), .A2(n464), .ZN(n462) );
  NAND2_X1 U491 ( .A1(n448), .A2(n468), .ZN(n673) );
  NAND2_X1 U492 ( .A1(n470), .A2(n469), .ZN(n468) );
  AND2_X1 U493 ( .A1(n472), .A2(n471), .ZN(n448) );
  NAND2_X1 U494 ( .A1(n378), .A2(n623), .ZN(n517) );
  NOR2_X1 U495 ( .A1(n640), .A2(n719), .ZN(n647) );
  XNOR2_X1 U496 ( .A(n601), .B(n600), .ZN(n681) );
  XNOR2_X1 U497 ( .A(n394), .B(n392), .ZN(n536) );
  XNOR2_X1 U498 ( .A(n576), .B(n494), .ZN(n582) );
  XNOR2_X1 U499 ( .A(n577), .B(n495), .ZN(n494) );
  XNOR2_X1 U500 ( .A(n423), .B(n575), .ZN(n576) );
  NAND2_X1 U501 ( .A1(n459), .A2(n458), .ZN(n457) );
  XNOR2_X1 U502 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U503 ( .A1(n407), .A2(n369), .ZN(n402) );
  NAND2_X1 U504 ( .A1(n621), .A2(n374), .ZN(n398) );
  XNOR2_X1 U505 ( .A(n759), .B(n493), .ZN(n762) );
  XNOR2_X1 U506 ( .A(n761), .B(n760), .ZN(n493) );
  XNOR2_X1 U507 ( .A(n505), .B(n504), .ZN(G75) );
  XNOR2_X1 U508 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n504) );
  NAND2_X1 U509 ( .A1(n370), .A2(n365), .ZN(n505) );
  XNOR2_X1 U510 ( .A(n398), .B(G110), .ZN(G12) );
  NOR2_X1 U511 ( .A1(n744), .A2(G953), .ZN(n365) );
  XOR2_X1 U512 ( .A(n547), .B(n546), .Z(n366) );
  AND2_X1 U513 ( .A1(n403), .A2(n387), .ZN(n367) );
  AND2_X1 U514 ( .A1(n449), .A2(n630), .ZN(n368) );
  NOR2_X1 U515 ( .A1(n602), .A2(n537), .ZN(n369) );
  XOR2_X1 U516 ( .A(KEYINPUT84), .B(n743), .Z(n370) );
  XOR2_X1 U517 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n371) );
  AND2_X1 U518 ( .A1(n610), .A2(KEYINPUT44), .ZN(n372) );
  XNOR2_X1 U519 ( .A(n588), .B(n587), .ZN(n373) );
  AND2_X1 U520 ( .A1(n619), .A2(n630), .ZN(n374) );
  AND2_X1 U521 ( .A1(n647), .A2(n619), .ZN(n375) );
  XOR2_X1 U522 ( .A(n657), .B(KEYINPUT40), .Z(n376) );
  XNOR2_X1 U523 ( .A(KEYINPUT28), .B(KEYINPUT109), .ZN(n377) );
  OR2_X1 U524 ( .A1(n554), .A2(n553), .ZN(n378) );
  XOR2_X1 U525 ( .A(n681), .B(KEYINPUT62), .Z(n379) );
  XNOR2_X1 U526 ( .A(KEYINPUT86), .B(KEYINPUT45), .ZN(n380) );
  XOR2_X1 U527 ( .A(n753), .B(n752), .Z(n381) );
  INV_X1 U528 ( .A(KEYINPUT75), .ZN(n419) );
  INV_X1 U529 ( .A(KEYINPUT48), .ZN(n437) );
  NOR2_X1 U530 ( .A1(G952), .A2(n784), .ZN(n768) );
  INV_X1 U531 ( .A(n768), .ZN(n531) );
  NAND2_X1 U532 ( .A1(n707), .A2(KEYINPUT39), .ZN(n471) );
  BUF_X1 U533 ( .A(n641), .Z(n382) );
  NAND2_X1 U534 ( .A1(n528), .A2(n531), .ZN(n527) );
  NAND2_X1 U535 ( .A1(n532), .A2(n531), .ZN(n530) );
  AND2_X1 U536 ( .A1(n514), .A2(n515), .ZN(n383) );
  AND2_X1 U537 ( .A1(n514), .A2(n515), .ZN(n384) );
  AND2_X2 U538 ( .A1(n514), .A2(n515), .ZN(n764) );
  NAND2_X1 U539 ( .A1(n413), .A2(KEYINPUT75), .ZN(n412) );
  BUF_X1 U540 ( .A(n635), .Z(n385) );
  NOR2_X1 U541 ( .A1(n656), .A2(n464), .ZN(n458) );
  AND2_X1 U542 ( .A1(n782), .A2(n387), .ZN(n741) );
  NAND2_X1 U543 ( .A1(n387), .A2(n784), .ZN(n772) );
  NAND2_X1 U544 ( .A1(n409), .A2(n387), .ZN(n404) );
  XNOR2_X2 U545 ( .A(n420), .B(n380), .ZN(n387) );
  INV_X1 U546 ( .A(n388), .ZN(n438) );
  NAND2_X1 U547 ( .A1(n665), .A2(n664), .ZN(n388) );
  NAND2_X1 U548 ( .A1(n388), .A2(n437), .ZN(n436) );
  XNOR2_X1 U549 ( .A(n389), .B(n581), .ZN(n544) );
  NAND2_X1 U550 ( .A1(n390), .A2(n496), .ZN(n489) );
  AND2_X1 U551 ( .A1(n390), .A2(n445), .ZN(n618) );
  XNOR2_X2 U552 ( .A(n516), .B(KEYINPUT0), .ZN(n390) );
  NAND2_X1 U553 ( .A1(n391), .A2(KEYINPUT39), .ZN(n472) );
  NAND2_X1 U554 ( .A1(n649), .A2(n648), .ZN(n391) );
  INV_X1 U555 ( .A(n391), .ZN(n470) );
  AND2_X1 U556 ( .A1(n470), .A2(n488), .ZN(n650) );
  NAND2_X1 U557 ( .A1(n791), .A2(n398), .ZN(n609) );
  AND2_X1 U558 ( .A1(n399), .A2(n375), .ZN(n684) );
  NAND2_X1 U559 ( .A1(n400), .A2(n465), .ZN(n455) );
  NAND2_X1 U560 ( .A1(n401), .A2(n456), .ZN(n400) );
  NAND2_X1 U561 ( .A1(n416), .A2(n412), .ZN(n411) );
  INV_X1 U562 ( .A(KEYINPUT46), .ZN(n465) );
  NAND2_X1 U563 ( .A1(n444), .A2(n439), .ZN(n540) );
  NOR2_X1 U564 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U565 ( .A(n529), .B(n381), .ZN(n528) );
  XNOR2_X1 U566 ( .A(n533), .B(n379), .ZN(n532) );
  NAND2_X1 U567 ( .A1(n427), .A2(n419), .ZN(n418) );
  XNOR2_X2 U568 ( .A(n406), .B(n405), .ZN(n730) );
  NAND2_X1 U569 ( .A1(n429), .A2(n427), .ZN(n782) );
  INV_X1 U570 ( .A(n427), .ZN(n413) );
  INV_X1 U571 ( .A(n429), .ZN(n415) );
  INV_X1 U572 ( .A(n418), .ZN(n417) );
  NAND2_X1 U573 ( .A1(n521), .A2(n524), .ZN(n420) );
  INV_X1 U574 ( .A(n717), .ZN(n421) );
  NAND2_X1 U575 ( .A1(n434), .A2(n436), .ZN(n428) );
  NOR2_X1 U576 ( .A1(n433), .A2(n432), .ZN(n431) );
  NAND2_X1 U577 ( .A1(n435), .A2(n437), .ZN(n434) );
  NAND2_X1 U578 ( .A1(n658), .A2(n486), .ZN(n435) );
  INV_X1 U579 ( .A(n699), .ZN(n442) );
  INV_X1 U580 ( .A(n684), .ZN(n443) );
  INV_X1 U581 ( .A(n682), .ZN(n444) );
  INV_X1 U582 ( .A(n727), .ZN(n445) );
  INV_X1 U583 ( .A(n558), .ZN(n557) );
  NAND2_X1 U584 ( .A1(n368), .A2(n724), .ZN(n503) );
  XNOR2_X2 U585 ( .A(n447), .B(G131), .ZN(n578) );
  OR2_X2 U586 ( .A1(n681), .A2(G902), .ZN(n467) );
  NOR2_X1 U587 ( .A1(n646), .A2(n450), .ZN(n449) );
  INV_X1 U588 ( .A(n721), .ZN(n450) );
  XNOR2_X1 U589 ( .A(n451), .B(n474), .ZN(n599) );
  XNOR2_X2 U590 ( .A(n476), .B(KEYINPUT70), .ZN(n451) );
  NAND2_X1 U591 ( .A1(n460), .A2(n457), .ZN(n795) );
  NAND2_X1 U592 ( .A1(n455), .A2(n452), .ZN(n486) );
  NAND2_X1 U593 ( .A1(n453), .A2(n460), .ZN(n452) );
  NAND2_X1 U594 ( .A1(n457), .A2(KEYINPUT46), .ZN(n454) );
  INV_X1 U595 ( .A(n793), .ZN(n456) );
  INV_X1 U596 ( .A(n730), .ZN(n459) );
  INV_X1 U597 ( .A(n461), .ZN(n460) );
  NAND2_X1 U598 ( .A1(n463), .A2(n462), .ZN(n461) );
  NAND2_X1 U599 ( .A1(n730), .A2(n464), .ZN(n463) );
  NOR2_X2 U600 ( .A1(n655), .A2(n707), .ZN(n715) );
  XNOR2_X2 U601 ( .A(n488), .B(KEYINPUT38), .ZN(n707) );
  NAND2_X1 U602 ( .A1(n745), .A2(n678), .ZN(n466) );
  NAND2_X1 U603 ( .A1(n643), .A2(n711), .ZN(n644) );
  XNOR2_X2 U604 ( .A(n467), .B(G472), .ZN(n643) );
  NOR2_X1 U605 ( .A1(n707), .A2(KEYINPUT39), .ZN(n469) );
  NAND2_X1 U606 ( .A1(n673), .A2(n696), .ZN(n473) );
  XNOR2_X2 U607 ( .A(G119), .B(KEYINPUT3), .ZN(n476) );
  XNOR2_X1 U608 ( .A(n477), .B(n512), .ZN(n511) );
  XNOR2_X2 U609 ( .A(G143), .B(G128), .ZN(n477) );
  XNOR2_X1 U610 ( .A(n536), .B(n593), .ZN(n535) );
  XNOR2_X1 U611 ( .A(n485), .B(n484), .ZN(n611) );
  NAND2_X1 U612 ( .A1(n609), .A2(KEYINPUT44), .ZN(n485) );
  XNOR2_X1 U613 ( .A(n609), .B(KEYINPUT89), .ZN(n608) );
  NAND2_X1 U614 ( .A1(n608), .A2(n538), .ZN(n523) );
  XNOR2_X1 U615 ( .A(n523), .B(n522), .ZN(n521) );
  NOR2_X1 U616 ( .A1(n372), .A2(n540), .ZN(n525) );
  XNOR2_X1 U617 ( .A(n635), .B(n552), .ZN(n641) );
  XNOR2_X1 U618 ( .A(n564), .B(n562), .ZN(n497) );
  XNOR2_X1 U619 ( .A(n561), .B(n364), .ZN(n562) );
  XNOR2_X1 U620 ( .A(n535), .B(n780), .ZN(n763) );
  XNOR2_X1 U621 ( .A(n497), .B(n563), .ZN(n755) );
  NOR2_X1 U622 ( .A1(n610), .A2(KEYINPUT44), .ZN(n538) );
  NOR2_X2 U623 ( .A1(n748), .A2(n768), .ZN(n751) );
  NAND2_X1 U624 ( .A1(n672), .A2(n711), .ZN(n635) );
  XNOR2_X1 U625 ( .A(n498), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U626 ( .A1(n758), .A2(n768), .ZN(n498) );
  NAND2_X1 U627 ( .A1(n606), .A2(n651), .ZN(n499) );
  NOR2_X2 U628 ( .A1(n641), .A2(n517), .ZN(n516) );
  NAND2_X1 U629 ( .A1(n502), .A2(n501), .ZN(n500) );
  INV_X1 U630 ( .A(n640), .ZN(n501) );
  NAND2_X1 U631 ( .A1(n764), .A2(G475), .ZN(n757) );
  INV_X1 U632 ( .A(n367), .ZN(n515) );
  XNOR2_X2 U633 ( .A(n520), .B(G122), .ZN(n564) );
  XNOR2_X2 U634 ( .A(G113), .B(G104), .ZN(n520) );
  XNOR2_X1 U635 ( .A(n605), .B(n604), .ZN(n606) );
  BUF_X2 U636 ( .A(n643), .Z(n724) );
  XNOR2_X2 U637 ( .A(n585), .B(n584), .ZN(n640) );
  XNOR2_X2 U638 ( .A(n640), .B(KEYINPUT1), .ZN(n718) );
  INV_X1 U639 ( .A(n544), .ZN(n526) );
  XNOR2_X1 U640 ( .A(n527), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U641 ( .A1(n383), .A2(G469), .ZN(n529) );
  XNOR2_X1 U642 ( .A(n530), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U643 ( .A1(n384), .A2(G472), .ZN(n533) );
  XNOR2_X1 U644 ( .A(n647), .B(n534), .ZN(n648) );
  INV_X1 U645 ( .A(KEYINPUT107), .ZN(n534) );
  XNOR2_X1 U646 ( .A(n747), .B(n746), .ZN(n748) );
  XNOR2_X1 U647 ( .A(n757), .B(n756), .ZN(n758) );
  XNOR2_X2 U648 ( .A(n642), .B(KEYINPUT81), .ZN(n693) );
  OR2_X2 U649 ( .A1(n656), .A2(n382), .ZN(n642) );
  XOR2_X1 U650 ( .A(n620), .B(KEYINPUT80), .Z(n537) );
  XNOR2_X1 U651 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n539) );
  XNOR2_X1 U652 ( .A(n575), .B(n557), .ZN(n545) );
  XNOR2_X1 U653 ( .A(n574), .B(KEYINPUT102), .ZN(n655) );
  INV_X1 U654 ( .A(n704), .ZN(n674) );
  INV_X1 U655 ( .A(KEYINPUT82), .ZN(n549) );
  INV_X1 U656 ( .A(KEYINPUT90), .ZN(n636) );
  XNOR2_X1 U657 ( .A(n636), .B(KEYINPUT36), .ZN(n637) );
  INV_X1 U658 ( .A(KEYINPUT111), .ZN(n657) );
  XNOR2_X1 U659 ( .A(n573), .B(n572), .ZN(n614) );
  XNOR2_X1 U660 ( .A(n541), .B(KEYINPUT14), .ZN(n623) );
  XOR2_X1 U661 ( .A(KEYINPUT74), .B(n542), .Z(n548) );
  NAND2_X1 U662 ( .A1(n548), .A2(G214), .ZN(n711) );
  INV_X1 U663 ( .A(n545), .ZN(n543) );
  XOR2_X1 U664 ( .A(KEYINPUT66), .B(G101), .Z(n581) );
  NAND2_X1 U665 ( .A1(G224), .A2(n784), .ZN(n546) );
  NAND2_X1 U666 ( .A1(G210), .A2(n548), .ZN(n550) );
  INV_X1 U667 ( .A(KEYINPUT19), .ZN(n552) );
  NAND2_X1 U668 ( .A1(n784), .A2(G952), .ZN(n627) );
  INV_X1 U669 ( .A(n627), .ZN(n554) );
  NOR2_X1 U670 ( .A1(G898), .A2(n624), .ZN(n553) );
  NAND2_X1 U671 ( .A1(n678), .A2(G234), .ZN(n555) );
  XNOR2_X1 U672 ( .A(n555), .B(KEYINPUT20), .ZN(n586) );
  NAND2_X1 U673 ( .A1(G221), .A2(n586), .ZN(n556) );
  XOR2_X1 U674 ( .A(KEYINPUT21), .B(n556), .Z(n721) );
  NAND2_X1 U675 ( .A1(G214), .A2(n597), .ZN(n559) );
  XNOR2_X1 U676 ( .A(n559), .B(n591), .ZN(n563) );
  XNOR2_X1 U677 ( .A(n578), .B(KEYINPUT11), .ZN(n561) );
  XNOR2_X1 U678 ( .A(G143), .B(G140), .ZN(n560) );
  NOR2_X1 U679 ( .A1(G902), .A2(n755), .ZN(n566) );
  XNOR2_X1 U680 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n565) );
  NAND2_X1 U681 ( .A1(G217), .A2(n592), .ZN(n567) );
  XNOR2_X1 U682 ( .A(G134), .B(n569), .ZN(n571) );
  NOR2_X1 U683 ( .A1(n761), .A2(G902), .ZN(n573) );
  XNOR2_X1 U684 ( .A(KEYINPUT100), .B(G478), .ZN(n572) );
  NAND2_X1 U685 ( .A1(n612), .A2(n614), .ZN(n574) );
  INV_X1 U686 ( .A(n655), .ZN(n710) );
  NAND2_X1 U687 ( .A1(G227), .A2(n784), .ZN(n577) );
  XNOR2_X1 U688 ( .A(n601), .B(n582), .ZN(n753) );
  NOR2_X1 U689 ( .A1(n753), .A2(G902), .ZN(n585) );
  XOR2_X1 U690 ( .A(G469), .B(KEYINPUT69), .Z(n583) );
  XNOR2_X1 U691 ( .A(KEYINPUT68), .B(n583), .ZN(n584) );
  XOR2_X1 U692 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n588) );
  NAND2_X1 U693 ( .A1(n586), .A2(G217), .ZN(n587) );
  INV_X1 U694 ( .A(n589), .ZN(n590) );
  NAND2_X1 U695 ( .A1(G221), .A2(n592), .ZN(n593) );
  NOR2_X1 U696 ( .A1(G902), .A2(n763), .ZN(n594) );
  NOR2_X1 U697 ( .A1(n718), .A2(n487), .ZN(n595) );
  XOR2_X1 U698 ( .A(KEYINPUT104), .B(n595), .Z(n602) );
  NAND2_X1 U699 ( .A1(n597), .A2(G210), .ZN(n598) );
  XNOR2_X1 U700 ( .A(n599), .B(n598), .ZN(n600) );
  XOR2_X1 U701 ( .A(n643), .B(KEYINPUT6), .Z(n631) );
  INV_X1 U702 ( .A(n631), .ZN(n620) );
  INV_X1 U703 ( .A(n724), .ZN(n619) );
  INV_X1 U704 ( .A(n718), .ZN(n669) );
  XNOR2_X1 U705 ( .A(KEYINPUT35), .B(KEYINPUT78), .ZN(n607) );
  NOR2_X1 U706 ( .A1(n719), .A2(n718), .ZN(n616) );
  NAND2_X1 U707 ( .A1(n631), .A2(n616), .ZN(n603) );
  NOR2_X1 U708 ( .A1(n614), .A2(n612), .ZN(n651) );
  INV_X1 U709 ( .A(n610), .ZN(n792) );
  INV_X1 U710 ( .A(n612), .ZN(n613) );
  NAND2_X1 U711 ( .A1(n613), .A2(n614), .ZN(n633) );
  INV_X1 U712 ( .A(n633), .ZN(n696) );
  NOR2_X1 U713 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U714 ( .A(KEYINPUT101), .B(n615), .Z(n698) );
  NOR2_X1 U715 ( .A1(n696), .A2(n698), .ZN(n708) );
  NAND2_X1 U716 ( .A1(n616), .A2(n724), .ZN(n727) );
  XNOR2_X1 U717 ( .A(KEYINPUT31), .B(KEYINPUT95), .ZN(n617) );
  XNOR2_X1 U718 ( .A(n618), .B(n617), .ZN(n699) );
  NAND2_X1 U719 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U720 ( .A1(n630), .A2(n622), .ZN(n682) );
  INV_X1 U721 ( .A(n623), .ZN(n737) );
  NOR2_X1 U722 ( .A1(n737), .A2(n624), .ZN(n625) );
  XNOR2_X1 U723 ( .A(n625), .B(KEYINPUT105), .ZN(n626) );
  NOR2_X1 U724 ( .A1(G900), .A2(n626), .ZN(n629) );
  NOR2_X1 U725 ( .A1(n627), .A2(n737), .ZN(n628) );
  NOR2_X1 U726 ( .A1(n629), .A2(n628), .ZN(n646) );
  NAND2_X1 U727 ( .A1(n631), .A2(n368), .ZN(n632) );
  XOR2_X1 U728 ( .A(KEYINPUT112), .B(n666), .Z(n634) );
  NOR2_X1 U729 ( .A1(n385), .A2(n634), .ZN(n638) );
  NOR2_X1 U730 ( .A1(n718), .A2(n639), .ZN(n702) );
  NAND2_X1 U731 ( .A1(n693), .A2(KEYINPUT83), .ZN(n653) );
  XNOR2_X1 U732 ( .A(n644), .B(KEYINPUT30), .ZN(n645) );
  NOR2_X1 U733 ( .A1(n646), .A2(n645), .ZN(n649) );
  XNOR2_X1 U734 ( .A(KEYINPUT108), .B(n650), .ZN(n652) );
  NAND2_X1 U735 ( .A1(n652), .A2(n651), .ZN(n692) );
  NAND2_X1 U736 ( .A1(n653), .A2(n692), .ZN(n654) );
  NOR2_X1 U737 ( .A1(n702), .A2(n654), .ZN(n658) );
  INV_X1 U738 ( .A(n708), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n693), .A2(n662), .ZN(n659) );
  XNOR2_X1 U740 ( .A(n659), .B(KEYINPUT47), .ZN(n661) );
  INV_X1 U741 ( .A(KEYINPUT83), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U743 ( .A1(KEYINPUT47), .A2(n662), .ZN(n663) );
  NAND2_X1 U744 ( .A1(n663), .A2(KEYINPUT83), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n666), .A2(n711), .ZN(n667) );
  XNOR2_X1 U746 ( .A(KEYINPUT106), .B(n667), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n670), .B(KEYINPUT43), .ZN(n671) );
  NOR2_X1 U748 ( .A1(n488), .A2(n671), .ZN(n705) );
  NAND2_X1 U749 ( .A1(n698), .A2(n673), .ZN(n704) );
  NAND2_X1 U750 ( .A1(n782), .A2(KEYINPUT2), .ZN(n676) );
  INV_X1 U751 ( .A(n678), .ZN(n677) );
  XNOR2_X1 U752 ( .A(n678), .B(KEYINPUT85), .ZN(n679) );
  NAND2_X1 U753 ( .A1(n679), .A2(KEYINPUT2), .ZN(n680) );
  XOR2_X1 U754 ( .A(n682), .B(G101), .Z(G3) );
  NAND2_X1 U755 ( .A1(n684), .A2(n696), .ZN(n683) );
  XNOR2_X1 U756 ( .A(n683), .B(G104), .ZN(G6) );
  XOR2_X1 U757 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n686) );
  NAND2_X1 U758 ( .A1(n684), .A2(n698), .ZN(n685) );
  XNOR2_X1 U759 ( .A(n686), .B(n685), .ZN(n688) );
  XOR2_X1 U760 ( .A(G107), .B(KEYINPUT27), .Z(n687) );
  XNOR2_X1 U761 ( .A(n688), .B(n687), .ZN(G9) );
  XOR2_X1 U762 ( .A(KEYINPUT29), .B(KEYINPUT114), .Z(n690) );
  NAND2_X1 U763 ( .A1(n693), .A2(n698), .ZN(n689) );
  XNOR2_X1 U764 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U765 ( .A(G128), .B(n691), .ZN(G30) );
  XNOR2_X1 U766 ( .A(G143), .B(n692), .ZN(G45) );
  XOR2_X1 U767 ( .A(G146), .B(KEYINPUT115), .Z(n695) );
  NAND2_X1 U768 ( .A1(n693), .A2(n696), .ZN(n694) );
  XNOR2_X1 U769 ( .A(n695), .B(n694), .ZN(G48) );
  NAND2_X1 U770 ( .A1(n699), .A2(n696), .ZN(n697) );
  XNOR2_X1 U771 ( .A(n697), .B(G113), .ZN(G15) );
  NAND2_X1 U772 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U773 ( .A(n700), .B(KEYINPUT116), .ZN(n701) );
  XNOR2_X1 U774 ( .A(G116), .B(n701), .ZN(G18) );
  XNOR2_X1 U775 ( .A(G125), .B(n702), .ZN(n703) );
  XNOR2_X1 U776 ( .A(n703), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U777 ( .A(G134), .B(n704), .ZN(G36) );
  XNOR2_X1 U778 ( .A(G140), .B(n705), .ZN(n706) );
  XNOR2_X1 U779 ( .A(n706), .B(KEYINPUT117), .ZN(G42) );
  OR2_X1 U780 ( .A1(n730), .A2(n717), .ZN(n740) );
  NOR2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n713) );
  INV_X1 U783 ( .A(n711), .ZN(n712) );
  NOR2_X1 U784 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n733) );
  NAND2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U788 ( .A(n720), .B(KEYINPUT50), .ZN(n726) );
  NOR2_X1 U789 ( .A1(n721), .A2(n487), .ZN(n722) );
  XOR2_X1 U790 ( .A(KEYINPUT49), .B(n722), .Z(n723) );
  NOR2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U792 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U793 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U794 ( .A(KEYINPUT51), .B(n729), .ZN(n731) );
  NOR2_X1 U795 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U796 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U797 ( .A(n734), .B(KEYINPUT52), .ZN(n735) );
  XNOR2_X1 U798 ( .A(KEYINPUT118), .B(n735), .ZN(n736) );
  NOR2_X1 U799 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U800 ( .A1(n738), .A2(G952), .ZN(n739) );
  NAND2_X1 U801 ( .A1(n740), .A2(n739), .ZN(n744) );
  NOR2_X1 U802 ( .A1(KEYINPUT2), .A2(n741), .ZN(n742) );
  NOR2_X1 U803 ( .A1(n742), .A2(n367), .ZN(n743) );
  NAND2_X1 U804 ( .A1(n764), .A2(G210), .ZN(n747) );
  XNOR2_X1 U805 ( .A(n745), .B(n539), .ZN(n746) );
  XNOR2_X1 U806 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n749) );
  XNOR2_X1 U807 ( .A(n749), .B(KEYINPUT88), .ZN(n750) );
  XNOR2_X1 U808 ( .A(n751), .B(n750), .ZN(G51) );
  XOR2_X1 U809 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n752) );
  XOR2_X1 U810 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n754) );
  XOR2_X1 U811 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n760) );
  NAND2_X1 U812 ( .A1(n383), .A2(G478), .ZN(n759) );
  NOR2_X1 U813 ( .A1(n768), .A2(n762), .ZN(G63) );
  XOR2_X1 U814 ( .A(n763), .B(KEYINPUT125), .Z(n766) );
  NAND2_X1 U815 ( .A1(n384), .A2(G217), .ZN(n765) );
  XNOR2_X1 U816 ( .A(n766), .B(n765), .ZN(n767) );
  NOR2_X1 U817 ( .A1(n768), .A2(n767), .ZN(G66) );
  NAND2_X1 U818 ( .A1(G953), .A2(G224), .ZN(n769) );
  XNOR2_X1 U819 ( .A(KEYINPUT61), .B(n769), .ZN(n770) );
  NAND2_X1 U820 ( .A1(n770), .A2(G898), .ZN(n771) );
  NAND2_X1 U821 ( .A1(n772), .A2(n771), .ZN(n778) );
  XNOR2_X1 U822 ( .A(n773), .B(G101), .ZN(n774) );
  XNOR2_X1 U823 ( .A(n774), .B(G110), .ZN(n776) );
  NOR2_X1 U824 ( .A1(G898), .A2(n784), .ZN(n775) );
  NOR2_X1 U825 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U826 ( .A(n778), .B(n777), .ZN(n779) );
  XNOR2_X1 U827 ( .A(KEYINPUT126), .B(n779), .ZN(G69) );
  XOR2_X1 U828 ( .A(n781), .B(n780), .Z(n786) );
  INV_X1 U829 ( .A(n786), .ZN(n783) );
  XNOR2_X1 U830 ( .A(n783), .B(n782), .ZN(n785) );
  NAND2_X1 U831 ( .A1(n785), .A2(n784), .ZN(n790) );
  XNOR2_X1 U832 ( .A(G227), .B(n786), .ZN(n787) );
  NAND2_X1 U833 ( .A1(n787), .A2(G900), .ZN(n788) );
  NAND2_X1 U834 ( .A1(n788), .A2(G953), .ZN(n789) );
  NAND2_X1 U835 ( .A1(n790), .A2(n789), .ZN(G72) );
  XNOR2_X1 U836 ( .A(n791), .B(G119), .ZN(G21) );
  XNOR2_X1 U837 ( .A(G122), .B(n792), .ZN(G24) );
  XNOR2_X1 U838 ( .A(G131), .B(KEYINPUT127), .ZN(n794) );
  XNOR2_X1 U839 ( .A(n794), .B(n793), .ZN(G33) );
  XOR2_X1 U840 ( .A(G137), .B(n795), .Z(G39) );
endmodule

