//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .A4(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n201));
  AOI22_X1  g015(.A1(new_n201), .A2(G128), .B1(new_n197), .B2(new_n199), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT64), .B1(new_n207), .B2(G137), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n205), .A2(G134), .ZN(new_n209));
  OAI211_X1 g023(.A(G131), .B(new_n206), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n207), .B2(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(G137), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n203), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n197), .A2(new_n199), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G143), .B(G146), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT0), .B(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n225), .B2(new_n216), .ZN(new_n226));
  NOR3_X1   g040(.A1(new_n218), .A2(new_n226), .A3(KEYINPUT30), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT30), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n216), .ZN(new_n229));
  INV_X1    g043(.A(new_n223), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n216), .B(new_n210), .C1(new_n200), .C2(new_n202), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n194), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NOR2_X1   g049(.A1(G237), .A2(G953), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G210), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n237), .B(KEYINPUT27), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT26), .B(G101), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n194), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n241), .A3(new_n232), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n234), .A2(new_n235), .A3(new_n240), .A4(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT31), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n242), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT30), .B1(new_n218), .B2(new_n226), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n231), .A2(new_n228), .A3(new_n232), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n246), .B1(new_n249), .B2(new_n194), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(new_n235), .A3(KEYINPUT31), .A4(new_n240), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n242), .A2(KEYINPUT67), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT67), .B1(new_n242), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n217), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n201), .A2(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n197), .A2(new_n199), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n221), .A2(G128), .A3(new_n201), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n256), .A2(new_n261), .B1(new_n229), .B2(new_n230), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT66), .B1(new_n262), .B2(new_n241), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n264), .B(new_n194), .C1(new_n218), .C2(new_n226), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n246), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n255), .B1(new_n266), .B2(new_n252), .ZN(new_n267));
  INV_X1    g081(.A(new_n240), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n245), .A2(new_n251), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(G472), .A2(G902), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n187), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n245), .A2(new_n251), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n267), .A2(new_n268), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT68), .A3(new_n270), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT69), .B(KEYINPUT32), .Z(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n267), .A2(new_n268), .ZN(new_n279));
  INV_X1    g093(.A(new_n250), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n279), .A2(new_n282), .A3(KEYINPUT29), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n262), .A2(new_n241), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(new_n246), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n255), .B1(new_n252), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n240), .A2(KEYINPUT29), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(G472), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT70), .B1(new_n291), .B2(KEYINPUT32), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n291), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n278), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n291), .A2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n291), .A2(KEYINPUT70), .A3(KEYINPUT32), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n301), .A2(KEYINPUT71), .A3(new_n290), .A4(new_n278), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  INV_X1    g119(.A(G125), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G140), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT74), .A4(KEYINPUT16), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT16), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n305), .B2(KEYINPUT16), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n196), .B(new_n308), .C1(new_n309), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT75), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n308), .B1(new_n309), .B2(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G146), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n306), .A2(G140), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT16), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n305), .A2(new_n307), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n318), .B(new_n310), .C1(new_n319), .C2(new_n317), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT75), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n196), .A4(new_n308), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n313), .A2(new_n315), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n188), .B2(G128), .ZN(new_n325));
  INV_X1    g139(.A(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT23), .A3(G119), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n188), .A2(G128), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n325), .A2(new_n327), .A3(new_n331), .A4(new_n328), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(G110), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n326), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n328), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT24), .B(G110), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n333), .A2(new_n334), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n323), .B(new_n340), .C1(new_n334), .C2(new_n333), .ZN(new_n341));
  OAI22_X1  g155(.A1(new_n337), .A2(new_n339), .B1(new_n329), .B2(G110), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(KEYINPUT76), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n305), .A2(new_n307), .A3(new_n196), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n343), .A2(new_n344), .A3(new_n315), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G137), .ZN(new_n348));
  INV_X1    g162(.A(G953), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n348), .B(new_n350), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n341), .A2(new_n346), .A3(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G217), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(G234), .B2(new_n284), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n353), .A2(new_n284), .A3(new_n354), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT25), .A4(new_n284), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n360), .B1(new_n365), .B2(new_n357), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  OAI21_X1  g181(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  AND2_X1   g185(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n372));
  NOR2_X1   g186(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G101), .ZN(new_n375));
  OAI22_X1  g189(.A1(new_n370), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(G107), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n374), .A2(new_n375), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G104), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n375), .B1(new_n380), .B2(new_n377), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n261), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n261), .B1(new_n378), .B2(new_n382), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n229), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT12), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n225), .A2(new_n216), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n380), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(new_n377), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n378), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n395), .B(G101), .C1(new_n391), .C2(new_n392), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n230), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n391), .A2(new_n392), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n381), .B1(new_n399), .B2(new_n375), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n400), .B2(new_n261), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n378), .A2(new_n382), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n402), .A2(new_n203), .A3(KEYINPUT10), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n388), .B(new_n397), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n349), .A2(G227), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n203), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n383), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT12), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n229), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n387), .A2(new_n404), .A3(new_n408), .A4(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT78), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n411), .B1(new_n410), .B2(new_n229), .ZN(new_n416));
  AOI211_X1 g230(.A(KEYINPUT12), .B(new_n388), .C1(new_n409), .C2(new_n383), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(KEYINPUT78), .A3(new_n404), .A4(new_n408), .ZN(new_n419));
  INV_X1    g233(.A(new_n404), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n400), .A2(new_n398), .A3(new_n261), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n383), .A2(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n388), .B1(new_n423), .B2(new_n397), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n407), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n415), .A2(new_n419), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G469), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n284), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT79), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n426), .A2(KEYINPUT79), .A3(new_n427), .A4(new_n284), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n408), .B1(new_n420), .B2(new_n424), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n418), .A2(new_n404), .A3(new_n407), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G469), .B1(new_n435), .B2(G902), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n369), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n438), .B(KEYINPUT89), .Z(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G122), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n394), .A2(new_n194), .A3(new_n396), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT81), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n394), .A2(new_n445), .A3(new_n194), .A4(new_n396), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n192), .A2(new_n193), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(new_n189), .ZN(new_n449));
  INV_X1    g263(.A(G113), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n189), .A3(new_n191), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n447), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n400), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n441), .B1(new_n444), .B2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n443), .A2(new_n440), .A3(new_n446), .A4(new_n454), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n456), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(KEYINPUT6), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n446), .A2(new_n454), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n440), .B1(new_n460), .B2(new_n443), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n441), .C1(new_n444), .C2(new_n455), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT83), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n458), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n223), .A2(G125), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT84), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n261), .B2(G125), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n203), .A2(KEYINPUT85), .A3(new_n306), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n349), .A2(G224), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n473), .A2(new_n479), .B1(G125), .B2(new_n223), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n479), .B2(new_n473), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n482), .A2(KEYINPUT88), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(KEYINPUT88), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n475), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT5), .ZN(new_n487));
  OAI221_X1 g301(.A(G113), .B1(new_n448), .B2(new_n189), .C1(new_n192), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n489));
  INV_X1    g303(.A(new_n447), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n400), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XOR2_X1   g307(.A(new_n440), .B(KEYINPUT8), .Z(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n453), .B2(new_n402), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n469), .A2(KEYINPUT7), .A3(new_n473), .A4(new_n475), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n486), .A2(new_n498), .A3(new_n457), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n499), .A2(new_n284), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n439), .B1(new_n478), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n465), .B(new_n464), .C1(new_n459), .C2(new_n461), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n476), .B1(new_n502), .B2(new_n458), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n499), .A2(new_n284), .ZN(new_n504));
  INV_X1    g318(.A(new_n439), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G214), .B1(G237), .B2(G902), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT80), .Z(new_n508));
  NOR3_X1   g322(.A1(new_n501), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G478), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n513), .A2(KEYINPUT13), .B1(new_n198), .B2(G128), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n513), .A2(KEYINPUT13), .ZN(new_n515));
  OAI21_X1  g329(.A(G134), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G128), .B(G143), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n516), .A2(new_n518), .ZN(new_n520));
  OR2_X1    g334(.A1(KEYINPUT96), .A2(G122), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT96), .A2(G122), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G116), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n190), .A2(G122), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n379), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n190), .B1(new_n521), .B2(new_n522), .ZN(new_n527));
  INV_X1    g341(.A(new_n525), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n527), .A2(G107), .A3(new_n528), .ZN(new_n529));
  OAI22_X1  g343(.A1(new_n519), .A2(new_n520), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n529), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n525), .B(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g346(.A(G107), .B1(new_n532), .B2(new_n527), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n517), .B(new_n207), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n367), .A2(new_n356), .A3(G953), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n535), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n512), .B1(new_n541), .B2(new_n284), .ZN(new_n542));
  AOI211_X1 g356(.A(G902), .B(new_n511), .C1(new_n539), .C2(new_n540), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(G234), .A2(G237), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(G902), .A3(G953), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT21), .B(G898), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n349), .A2(G952), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n547), .A2(new_n548), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G475), .ZN(new_n552));
  INV_X1    g366(.A(G237), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n349), .A3(G214), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n198), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n236), .A2(G143), .A3(G214), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(KEYINPUT18), .A2(G131), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT90), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT90), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n555), .A2(new_n561), .A3(new_n556), .A4(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n319), .A2(G146), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n557), .A2(new_n559), .B1(new_n564), .B2(new_n345), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n554), .A2(new_n198), .ZN(new_n567));
  AOI21_X1  g381(.A(G143), .B1(new_n236), .B2(G214), .ZN(new_n568));
  OAI21_X1  g382(.A(G131), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n555), .A2(new_n214), .A3(new_n556), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n557), .A2(KEYINPUT17), .A3(G131), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n566), .B1(new_n323), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(G113), .B(G122), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(new_n370), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n566), .B(new_n577), .C1(new_n323), .C2(new_n574), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n284), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n552), .B1(new_n582), .B2(KEYINPUT95), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n579), .B2(new_n580), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT19), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n304), .A2(G125), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n316), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT19), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT91), .B1(new_n592), .B2(new_n196), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT91), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n594), .B(G146), .C1(new_n590), .C2(new_n591), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n314), .A2(G146), .B1(new_n569), .B2(new_n571), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n596), .A2(new_n597), .B1(new_n563), .B2(new_n565), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT92), .B1(new_n598), .B2(new_n577), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT19), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT19), .B1(new_n305), .B2(new_n307), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n196), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n594), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n569), .A2(new_n571), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n592), .A2(KEYINPUT91), .A3(new_n196), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n315), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n566), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n578), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n599), .A2(new_n580), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n552), .A2(new_n284), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT93), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT20), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n610), .B(new_n612), .C1(new_n614), .C2(KEYINPUT20), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n551), .A2(new_n587), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n437), .A2(new_n509), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n303), .A2(new_n366), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  NAND2_X1  g437(.A1(new_n432), .A2(new_n436), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(new_n366), .A3(new_n368), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n501), .A2(new_n506), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n507), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n272), .A2(new_n276), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT98), .B1(new_n269), .B2(G902), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n275), .A2(new_n630), .A3(new_n284), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n631), .A3(G472), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n625), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n550), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n587), .A2(new_n617), .A3(new_n618), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n541), .B(KEYINPUT33), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n637), .A2(new_n510), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n541), .A2(new_n510), .A3(new_n284), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n510), .A2(new_n284), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n634), .A2(new_n635), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NOR2_X1   g462(.A1(new_n542), .A2(new_n543), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n583), .B2(new_n586), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n613), .A2(KEYINPUT20), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n610), .A2(new_n616), .A3(new_n612), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n550), .B(KEYINPUT99), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n634), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT35), .B(G107), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT100), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(G9));
  AND2_X1   g473(.A1(new_n437), .A2(new_n509), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n341), .A2(new_n661), .A3(new_n346), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n341), .B2(new_n346), .ZN(new_n664));
  OAI22_X1  g478(.A1(new_n663), .A2(new_n664), .B1(KEYINPUT36), .B2(new_n352), .ZN(new_n665));
  INV_X1    g479(.A(new_n664), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n662), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n365), .A2(new_n357), .B1(new_n669), .B2(new_n358), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n619), .A2(new_n670), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n671), .A2(new_n632), .A3(new_n628), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n660), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n549), .A2(new_n545), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT103), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT102), .B(G900), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n547), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n610), .A2(new_n616), .A3(new_n612), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n616), .B1(new_n610), .B2(new_n612), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n586), .ZN(new_n685));
  OAI21_X1  g499(.A(G475), .B1(new_n584), .B2(new_n585), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n544), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n680), .B1(new_n651), .B2(new_n652), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT104), .B1(new_n690), .B2(new_n650), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n507), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n501), .A2(new_n506), .A3(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n670), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n437), .A2(new_n692), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n303), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  XOR2_X1   g512(.A(new_n680), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n437), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n700), .B(KEYINPUT40), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n626), .B(KEYINPUT38), .ZN(new_n702));
  NAND2_X1  g516(.A1(G472), .A2(G902), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n280), .A2(new_n268), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n286), .B2(new_n240), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT105), .Z(new_n707));
  NAND3_X1  g521(.A1(new_n301), .A2(new_n278), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n636), .A2(new_n544), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n695), .A2(new_n709), .A3(new_n693), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n701), .A2(new_n702), .A3(new_n708), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND3_X1  g526(.A1(new_n437), .A2(new_n694), .A3(new_n695), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n636), .A2(new_n643), .A3(new_n681), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT106), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n636), .A2(new_n716), .A3(new_n643), .A4(new_n681), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n303), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  AOI21_X1  g535(.A(new_n427), .B1(new_n426), .B2(new_n284), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n430), .B2(new_n431), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n626), .A2(new_n507), .A3(new_n723), .A4(new_n368), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n645), .A2(new_n366), .A3(new_n635), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n303), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT41), .B(G113), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT107), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n728), .B(new_n730), .ZN(G15));
  INV_X1    g545(.A(new_n303), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n724), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n655), .A2(new_n366), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  NAND2_X1  g551(.A1(new_n733), .A2(new_n671), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  INV_X1    g553(.A(G472), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n275), .B2(new_n284), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n287), .A2(new_n268), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n271), .B1(new_n273), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n366), .A3(new_n654), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n723), .A2(new_n368), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n627), .A2(new_n745), .A3(new_n746), .A4(new_n709), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(G122), .Z(G24));
  NAND4_X1  g562(.A1(new_n715), .A2(new_n695), .A3(new_n717), .A4(new_n744), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n724), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n306), .ZN(G27));
  INV_X1    g565(.A(new_n366), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n291), .B(KEYINPUT32), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n290), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n753), .A2(new_n754), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n718), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n478), .A2(new_n439), .A3(new_n500), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n505), .B1(new_n503), .B2(new_n504), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n693), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n624), .A2(new_n762), .A3(new_n368), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n758), .A2(KEYINPUT42), .A3(new_n759), .A4(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n752), .B1(new_n296), .B2(new_n302), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT108), .A3(new_n759), .A4(new_n764), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT42), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n752), .B(new_n763), .C1(new_n296), .C2(new_n302), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT108), .B1(new_n770), .B2(new_n759), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n765), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  NAND3_X1  g587(.A1(new_n766), .A2(new_n692), .A3(new_n764), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  INV_X1    g589(.A(KEYINPUT46), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n435), .A2(KEYINPUT45), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n427), .B1(new_n435), .B2(KEYINPUT45), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n427), .A2(new_n284), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n779), .B(KEYINPUT46), .C1(new_n427), .C2(new_n284), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n432), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n368), .A3(new_n699), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n617), .A2(new_n618), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n587), .A3(new_n643), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT43), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n633), .A3(new_n695), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n785), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n789), .A2(KEYINPUT44), .A3(new_n633), .A4(new_n695), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n794), .A3(new_n762), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n794), .B1(new_n793), .B2(new_n762), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n205), .ZN(G39));
  NAND2_X1  g613(.A1(new_n784), .A2(new_n368), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(KEYINPUT47), .ZN(new_n802));
  XNOR2_X1  g616(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n803), .B1(new_n784), .B2(new_n368), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n762), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n718), .A2(new_n366), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n805), .A2(new_n732), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  INV_X1    g623(.A(new_n671), .ZN(new_n810));
  AOI221_X4 g624(.A(new_n724), .B1(new_n810), .B2(new_n734), .C1(new_n296), .C2(new_n302), .ZN(new_n811));
  AOI211_X1 g625(.A(new_n726), .B(new_n724), .C1(new_n296), .C2(new_n302), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n811), .A2(new_n812), .A3(new_n747), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n625), .A2(new_n633), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n786), .A2(new_n650), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n644), .A2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n509), .A2(new_n816), .A3(new_n654), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n814), .A2(new_n817), .B1(new_n660), .B2(new_n672), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n622), .A2(new_n818), .A3(KEYINPUT112), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT112), .B1(new_n622), .B2(new_n818), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n749), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n764), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n690), .A2(new_n587), .A3(new_n649), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n763), .A2(new_n670), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n303), .A3(KEYINPUT113), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT113), .B1(new_n825), .B2(new_n303), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n774), .B(new_n823), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n822), .A2(new_n725), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n627), .A2(new_n709), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n695), .A2(new_n680), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n437), .A3(new_n708), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n720), .A2(new_n697), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n750), .B1(new_n303), .B2(new_n696), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT52), .A3(new_n720), .A4(new_n834), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n830), .A2(KEYINPUT53), .A3(new_n772), .A4(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n303), .B(new_n725), .C1(new_n671), .C2(new_n735), .ZN(new_n842));
  INV_X1    g656(.A(new_n747), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n728), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n622), .A2(new_n818), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n622), .A2(new_n818), .A3(KEYINPUT112), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n774), .A2(new_n823), .ZN(new_n850));
  INV_X1    g664(.A(new_n828), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n850), .B1(new_n826), .B2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n840), .A3(new_n772), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n841), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n849), .A2(new_n840), .A3(new_n852), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(KEYINPUT114), .A3(KEYINPUT53), .A4(new_n772), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n746), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n693), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n702), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n702), .B2(new_n864), .ZN(new_n867));
  INV_X1    g681(.A(new_n677), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n366), .A2(new_n789), .A3(new_n868), .A4(new_n744), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n871), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  INV_X1    g689(.A(new_n805), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n723), .A2(new_n369), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n869), .A2(new_n762), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n708), .A2(new_n752), .A3(new_n676), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n806), .A2(new_n746), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n636), .A2(new_n643), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(KEYINPUT118), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n744), .A2(new_n695), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n789), .A2(new_n868), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n882), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT118), .B1(new_n883), .B2(new_n884), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n874), .A2(new_n880), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n758), .A2(new_n887), .A3(new_n882), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT48), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n883), .A2(new_n645), .B1(new_n869), .B2(new_n725), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n874), .A2(KEYINPUT117), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n876), .A2(KEYINPUT115), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n877), .B1(new_n805), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n879), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n872), .A2(new_n902), .A3(new_n873), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n897), .A2(new_n901), .A3(new_n903), .A4(new_n891), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n896), .B1(new_n875), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n841), .A2(new_n855), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n862), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n549), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n862), .A2(new_n905), .A3(KEYINPUT119), .A4(new_n908), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(G953), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n752), .A2(new_n508), .A3(new_n369), .ZN(new_n913));
  INV_X1    g727(.A(new_n723), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n787), .B(new_n913), .C1(KEYINPUT49), .C2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n702), .A2(new_n708), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n915), .B(new_n916), .C1(KEYINPUT49), .C2(new_n914), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n910), .A2(new_n912), .A3(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n349), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n857), .A2(G902), .A3(new_n439), .A4(new_n859), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n467), .B(new_n477), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT55), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n920), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n923), .B2(new_n925), .ZN(G51));
  XNOR2_X1  g741(.A(new_n781), .B(KEYINPUT57), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n857), .A2(KEYINPUT54), .A3(new_n859), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT54), .B1(new_n857), .B2(new_n859), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n426), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n857), .A2(G902), .A3(new_n780), .A4(new_n859), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n919), .B1(new_n932), .B2(new_n933), .ZN(G54));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n935));
  NAND2_X1  g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT120), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n857), .A2(G902), .A3(new_n859), .A4(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n610), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n920), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n939), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n935), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n919), .B1(new_n939), .B2(new_n940), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n945), .B(KEYINPUT121), .C1(new_n940), .C2(new_n939), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(G60));
  NOR2_X1   g761(.A1(new_n929), .A2(new_n930), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n640), .B(KEYINPUT59), .Z(new_n949));
  NAND2_X1  g763(.A1(new_n637), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n920), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n862), .A2(new_n908), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n637), .B1(new_n952), .B2(new_n949), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(G63));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT122), .Z(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT60), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n355), .B1(new_n860), .B2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n857), .A2(new_n669), .A3(new_n859), .A4(new_n957), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n959), .A2(new_n920), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n959), .A2(KEYINPUT61), .A3(new_n920), .A4(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G66));
  NOR2_X1   g779(.A1(new_n849), .A2(G953), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT123), .ZN(new_n967));
  INV_X1    g781(.A(G224), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n548), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n973));
  INV_X1    g787(.A(new_n467), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n349), .A2(G898), .ZN(new_n975));
  AOI22_X1  g789(.A1(new_n972), .A2(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n973), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n975), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n977), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n976), .A2(new_n979), .ZN(G69));
  XOR2_X1   g794(.A(new_n249), .B(new_n592), .Z(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(G900), .B2(G953), .ZN(new_n982));
  INV_X1    g796(.A(new_n785), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n758), .A2(new_n983), .A3(new_n832), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT126), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n985), .A2(new_n774), .A3(new_n808), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n796), .A2(new_n797), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n720), .A2(new_n697), .A3(new_n831), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n989), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n798), .A2(new_n991), .A3(KEYINPUT125), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n986), .B(new_n772), .C1(new_n990), .C2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n982), .B1(new_n993), .B2(G953), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n711), .A2(new_n989), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT62), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n816), .A2(new_n762), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n766), .A2(new_n437), .A3(new_n699), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n988), .A2(new_n808), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n981), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n994), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(KEYINPUT127), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n349), .B1(G227), .B2(G900), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n994), .A2(new_n1001), .A3(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1004), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n1008), .ZN(G72));
  OR2_X1    g823(.A1(new_n993), .A2(new_n821), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n703), .B(KEYINPUT63), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n240), .B(new_n280), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1011), .B1(new_n1000), .B2(new_n849), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n280), .A2(new_n240), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n920), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1012), .B1(new_n282), .B2(new_n704), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n841), .B2(new_n855), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1013), .A2(new_n1016), .A3(new_n1018), .ZN(G57));
endmodule


