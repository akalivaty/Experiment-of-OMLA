//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n194), .B2(new_n192), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT71), .B(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(G143), .B2(new_n187), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n191), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n188), .A2(new_n190), .A3(new_n199), .A4(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n198), .B1(new_n205), .B2(new_n197), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G224), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n206), .B(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G110), .B(G122), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G104), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(G107), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n216), .A2(G104), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n213), .A2(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n212), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n223), .A2(new_n212), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G116), .ZN(new_n228));
  INV_X1    g042(.A(G116), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT5), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(G113), .C1(KEYINPUT5), .C2(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n230), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n226), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n214), .A2(new_n217), .A3(new_n219), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n220), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n233), .B(new_n234), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n243), .A3(G101), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n238), .A2(new_n245), .A3(KEYINPUT80), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT80), .B1(new_n238), .B2(new_n245), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n211), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n238), .A2(new_n210), .A3(new_n245), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n245), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n238), .A2(new_n245), .A3(KEYINPUT80), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n210), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT6), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT81), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n256), .B(new_n211), .C1(new_n246), .C2(new_n247), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n209), .B(new_n250), .C1(new_n257), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n208), .A2(KEYINPUT7), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n206), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n226), .B(new_n236), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n210), .B(KEYINPUT8), .Z(new_n266));
  OAI21_X1  g080(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n264), .B(KEYINPUT82), .C1(new_n265), .C2(new_n266), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n249), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n261), .A2(new_n262), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G210), .B1(G237), .B2(G902), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n261), .A2(new_n262), .A3(new_n273), .A4(new_n271), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  XOR2_X1   g091(.A(KEYINPUT9), .B(G234), .Z(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G221), .B1(new_n279), .B2(G902), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n280), .B(KEYINPUT75), .ZN(new_n281));
  INV_X1    g095(.A(G469), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(new_n262), .ZN(new_n283));
  XOR2_X1   g097(.A(G110), .B(G140), .Z(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT76), .ZN(new_n285));
  INV_X1    g099(.A(G227), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(G953), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n285), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n204), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n241), .A2(new_n196), .A3(new_n244), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT11), .ZN(new_n293));
  INV_X1    g107(.A(G134), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(G137), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(G137), .ZN(new_n296));
  INV_X1    g110(.A(G137), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT11), .A3(G134), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G131), .ZN(new_n300));
  INV_X1    g114(.A(G131), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n295), .A2(new_n298), .A3(new_n301), .A4(new_n296), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n200), .A2(KEYINPUT78), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(G128), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n191), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n203), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n226), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT10), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n292), .A2(new_n304), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n304), .B1(new_n292), .B2(new_n314), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n289), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT79), .B1(new_n226), .B2(new_n204), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n223), .A2(new_n212), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n220), .A2(new_n223), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(new_n212), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n205), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n319), .A2(new_n324), .A3(new_n312), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n303), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT12), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT12), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n328), .A3(new_n303), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n327), .A2(new_n315), .A3(new_n288), .A4(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(G902), .B1(new_n318), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n283), .B1(new_n331), .B2(new_n282), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n315), .A3(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n289), .ZN(new_n334));
  INV_X1    g148(.A(new_n317), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n315), .A3(new_n288), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(G469), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n281), .B1(new_n332), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(G214), .B1(G237), .B2(G902), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n277), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G475), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n187), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n343), .B(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G125), .A2(G140), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n197), .B2(G140), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n345), .B1(new_n187), .B2(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(G237), .A2(G953), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G214), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n189), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(G143), .A3(G214), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT18), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n356), .B2(new_n301), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n301), .B1(new_n352), .B2(new_n353), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT18), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n349), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n301), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT17), .ZN(new_n362));
  INV_X1    g176(.A(new_n358), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT16), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n197), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n347), .B2(new_n365), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n187), .ZN(new_n369));
  OAI211_X1 g183(.A(G146), .B(new_n367), .C1(new_n347), .C2(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n358), .A2(KEYINPUT17), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n364), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(G113), .B(G122), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n213), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n360), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n361), .A2(KEYINPUT83), .A3(new_n363), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n354), .A2(G131), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n377), .B1(new_n378), .B2(new_n358), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT19), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n342), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n187), .B(new_n381), .C1(new_n348), .C2(new_n380), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n376), .A2(new_n379), .A3(new_n370), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n374), .B1(new_n360), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n341), .B(new_n262), .C1(new_n375), .C2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT20), .ZN(new_n386));
  INV_X1    g200(.A(G478), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n388));
  OR2_X1    g202(.A1(new_n388), .A2(KEYINPUT15), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(KEYINPUT15), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n387), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G122), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT14), .B1(new_n392), .B2(G116), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n229), .A3(G122), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(G116), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G107), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(G128), .B(G143), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(new_n294), .ZN(new_n402));
  XNOR2_X1  g216(.A(G116), .B(G122), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n216), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n397), .A2(KEYINPUT84), .A3(G107), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n400), .A2(new_n402), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n403), .B(new_n216), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n401), .A2(new_n294), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n189), .A2(KEYINPUT13), .A3(G128), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(G128), .B2(new_n189), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT13), .B1(new_n189), .B2(G128), .ZN(new_n411));
  OAI21_X1  g225(.A(G134), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n278), .A2(G217), .A3(new_n207), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n406), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n406), .B2(new_n413), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n262), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n391), .B1(new_n418), .B2(KEYINPUT86), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(KEYINPUT86), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(new_n391), .ZN(new_n421));
  NAND2_X1  g235(.A1(G234), .A2(G237), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(G952), .A3(new_n207), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G898), .Z(new_n424));
  NAND3_X1  g238(.A1(new_n422), .A2(G902), .A3(G953), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n374), .B1(new_n360), .B2(new_n372), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n262), .B1(new_n375), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G475), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n386), .A2(new_n421), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n385), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n385), .A2(new_n433), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n434), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT87), .A3(new_n426), .A4(new_n421), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n340), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n242), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n297), .A2(G134), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n294), .A2(G137), .ZN(new_n441));
  OAI21_X1  g255(.A(G131), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n204), .A2(new_n302), .A3(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n195), .A2(new_n193), .B1(new_n300), .B2(new_n302), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n445));
  NOR3_X1   g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n302), .A2(new_n442), .A3(KEYINPUT64), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT64), .B1(new_n302), .B2(new_n442), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n204), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT65), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n444), .ZN(new_n452));
  OAI211_X1 g266(.A(KEYINPUT65), .B(new_n204), .C1(new_n447), .C2(new_n448), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n439), .B(new_n446), .C1(new_n454), .C2(new_n445), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n350), .A2(G210), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT26), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n459), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n218), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(G101), .A3(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n443), .A2(new_n444), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n242), .B(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n455), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n454), .A2(new_n445), .ZN(new_n473));
  INV_X1    g287(.A(new_n446), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n242), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n469), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n465), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT67), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT31), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n477), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT31), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT28), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n454), .A2(new_n242), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(new_n469), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n476), .A2(KEYINPUT28), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT69), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n476), .B1(new_n242), .B2(new_n454), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n483), .B1(new_n492), .B2(new_n465), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n471), .B1(new_n455), .B2(new_n470), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n475), .A2(KEYINPUT67), .A3(new_n477), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n481), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(G472), .A2(G902), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT32), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(KEYINPUT32), .A3(new_n499), .ZN(new_n503));
  INV_X1    g317(.A(G472), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT29), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n475), .A2(new_n469), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n465), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n505), .B(new_n507), .C1(new_n492), .C2(new_n465), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n467), .B(new_n468), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n487), .B1(new_n509), .B2(KEYINPUT28), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n465), .A2(new_n505), .ZN(new_n511));
  AOI21_X1  g325(.A(G902), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n504), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n502), .A2(new_n503), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n207), .A2(G221), .A3(G234), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT73), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT22), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(new_n297), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n227), .A2(G128), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT70), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(G119), .B2(new_n201), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT24), .B(G110), .Z(new_n525));
  AOI22_X1  g339(.A1(new_n369), .A2(new_n370), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n201), .A2(G119), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT23), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n522), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G110), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n524), .A2(new_n525), .B1(new_n529), .B2(G110), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(new_n370), .A3(new_n345), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n520), .A2(new_n531), .A3(new_n533), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n262), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G217), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(G234), .B2(new_n262), .ZN(new_n542));
  AND2_X1   g356(.A1(new_n537), .A2(new_n539), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT74), .B1(new_n537), .B2(new_n539), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n540), .B(new_n542), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n535), .A2(new_n536), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n542), .A2(G902), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n438), .A2(new_n515), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G101), .ZN(G3));
  AOI21_X1  g365(.A(new_n504), .B1(new_n498), .B2(new_n262), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n553));
  INV_X1    g367(.A(new_n499), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT68), .B1(new_n496), .B2(KEYINPUT31), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  AOI211_X1 g370(.A(new_n480), .B(new_n556), .C1(new_n494), .C2(new_n495), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n558), .B2(new_n493), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT88), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n553), .A2(new_n560), .A3(new_n549), .A4(new_n338), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n561), .B(KEYINPUT89), .Z(new_n562));
  OR2_X1    g376(.A1(new_n416), .A2(new_n417), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT33), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n565), .A2(G478), .A3(new_n262), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n418), .A2(new_n387), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n436), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n277), .A2(new_n426), .A3(new_n339), .A4(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n562), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(new_n574), .B(KEYINPUT90), .Z(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT34), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(G104), .ZN(G6));
  NAND3_X1  g391(.A1(new_n434), .A2(new_n429), .A3(new_n435), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n421), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n277), .A2(new_n426), .A3(new_n339), .A4(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n562), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(new_n216), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT91), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT35), .ZN(G9));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n520), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT92), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n588), .A2(new_n534), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n534), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n548), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT93), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n591), .A2(new_n545), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n592), .B1(new_n591), .B2(new_n545), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n438), .A2(new_n553), .A3(new_n560), .A4(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT94), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT37), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(G110), .Z(G12));
  AOI21_X1  g414(.A(new_n513), .B1(new_n500), .B2(new_n501), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n595), .B1(new_n601), .B2(new_n503), .ZN(new_n602));
  INV_X1    g416(.A(new_n340), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n604));
  OR3_X1    g418(.A1(new_n425), .A2(new_n604), .A3(G900), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n425), .B2(G900), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n423), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n579), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n579), .A2(new_n610), .A3(new_n607), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n602), .A2(new_n603), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G128), .ZN(G30));
  XNOR2_X1  g428(.A(new_n607), .B(KEYINPUT39), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n338), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(KEYINPUT99), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT40), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n509), .A2(new_n465), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n496), .A2(G472), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(G472), .A2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT97), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n502), .A2(new_n503), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n591), .A2(new_n545), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n277), .B(KEYINPUT38), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n436), .A2(new_n421), .ZN(new_n628));
  INV_X1    g442(.A(new_n339), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n626), .A2(KEYINPUT98), .A3(new_n631), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n618), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT100), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(new_n189), .ZN(G45));
  NAND2_X1  g452(.A1(new_n277), .A2(new_n339), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n578), .A2(new_n569), .A3(new_n607), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  OR3_X1    g455(.A1(new_n639), .A2(new_n641), .A3(KEYINPUT101), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT101), .B1(new_n639), .B2(new_n641), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n602), .A2(new_n338), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G146), .ZN(G48));
  NOR2_X1   g459(.A1(new_n331), .A2(new_n282), .ZN(new_n646));
  AOI211_X1 g460(.A(G469), .B(G902), .C1(new_n318), .C2(new_n330), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n646), .A2(new_n647), .A3(new_n281), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT102), .Z(new_n649));
  NAND4_X1  g463(.A1(new_n649), .A2(new_n515), .A3(new_n549), .A4(new_n573), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT41), .B(G113), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G15));
  NAND4_X1  g466(.A1(new_n649), .A2(new_n515), .A3(new_n549), .A4(new_n581), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G116), .ZN(G18));
  NAND3_X1  g468(.A1(new_n277), .A2(new_n648), .A3(new_n339), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n277), .A2(new_n648), .A3(KEYINPUT103), .A4(new_n339), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n432), .A2(new_n437), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n602), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT104), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G119), .ZN(G21));
  NOR2_X1   g477(.A1(new_n510), .A2(new_n466), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n496), .B2(KEYINPUT31), .ZN(new_n665));
  INV_X1    g479(.A(new_n483), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n554), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n668));
  AOI21_X1  g482(.A(G902), .B1(new_n558), .B2(new_n493), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n668), .B1(new_n669), .B2(new_n504), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n552), .A2(KEYINPUT105), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n426), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n639), .A2(new_n673), .A3(new_n628), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n549), .A3(new_n649), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G122), .ZN(G24));
  NAND4_X1  g490(.A1(new_n672), .A2(new_n625), .A3(new_n640), .A4(new_n659), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G125), .ZN(G27));
  NAND4_X1  g492(.A1(new_n640), .A2(new_n275), .A3(new_n339), .A4(new_n276), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n336), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n335), .A2(KEYINPUT106), .A3(new_n315), .A4(new_n288), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n334), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n332), .B1(new_n282), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n281), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n515), .A2(new_n549), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n515), .A2(KEYINPUT107), .A3(new_n549), .A4(new_n687), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n559), .A2(KEYINPUT108), .A3(KEYINPUT32), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n503), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n601), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(KEYINPUT42), .A3(new_n549), .A4(new_n687), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G131), .ZN(G33));
  NAND3_X1  g514(.A1(new_n275), .A2(new_n339), .A3(new_n276), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n609), .A2(new_n702), .A3(new_n611), .ZN(new_n703));
  INV_X1    g517(.A(new_n686), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n703), .A2(new_n515), .A3(new_n549), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G134), .ZN(G36));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n683), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n334), .A2(new_n336), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n708), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n709), .A2(G469), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n707), .B1(new_n713), .B2(new_n283), .ZN(new_n714));
  INV_X1    g528(.A(new_n647), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n712), .B(KEYINPUT46), .C1(new_n282), .C2(new_n262), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n685), .A3(new_n615), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT109), .Z(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n553), .A2(new_n560), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n436), .A2(new_n569), .ZN(new_n722));
  XOR2_X1   g536(.A(new_n722), .B(KEYINPUT43), .Z(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n625), .A3(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n725), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n702), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT110), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n730), .A3(new_n702), .A4(new_n727), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n720), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G137), .ZN(G39));
  NAND2_X1  g547(.A1(new_n717), .A2(new_n685), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT47), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n717), .A2(new_n736), .A3(new_n685), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n738), .A2(new_n515), .A3(new_n549), .A4(new_n679), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n366), .ZN(G42));
  INV_X1    g554(.A(new_n648), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n701), .A3(new_n423), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n624), .A2(new_n549), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n436), .A3(new_n570), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n723), .A2(new_n742), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n625), .A3(new_n672), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n423), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n672), .A2(new_n549), .A3(new_n750), .A4(new_n723), .ZN(new_n751));
  INV_X1    g565(.A(new_n627), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n629), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n751), .A2(new_n741), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT50), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(KEYINPUT50), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n749), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n646), .A2(new_n647), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n735), .A2(new_n737), .B1(new_n281), .B2(new_n761), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n762), .A2(new_n701), .A3(new_n751), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT120), .B(new_n749), .C1(new_n756), .C2(new_n757), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n659), .ZN(new_n767));
  OAI211_X1 g581(.A(G952), .B(new_n207), .C1(new_n751), .C2(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n697), .A2(new_n549), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n746), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(KEYINPUT48), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n770), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(KEYINPUT48), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n766), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n778), .B1(new_n756), .B2(new_n757), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n754), .A2(KEYINPUT50), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n755), .A3(KEYINPUT118), .ZN(new_n781));
  AOI211_X1 g595(.A(new_n748), .B(new_n763), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n777), .B1(new_n782), .B2(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n781), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n749), .A3(new_n764), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(KEYINPUT119), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n776), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n743), .A2(new_n571), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n436), .A2(new_n421), .A3(new_n607), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n602), .A2(new_n338), .A3(new_n702), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n672), .A2(new_n625), .A3(new_n687), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n705), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n580), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n572), .B1(new_n580), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n550), .B(new_n597), .C1(new_n797), .C2(new_n561), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n650), .A2(new_n675), .A3(new_n653), .A4(new_n661), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n800), .A3(new_n699), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n502), .A2(new_n623), .A3(new_n503), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n639), .A2(new_n686), .A3(new_n628), .ZN(new_n804));
  INV_X1    g618(.A(new_n625), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n803), .A2(new_n804), .A3(new_n805), .A4(new_n607), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n677), .A2(new_n644), .A3(new_n613), .A4(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT52), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n799), .A2(new_n800), .A3(new_n699), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n644), .A2(new_n613), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n677), .A4(new_n806), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n807), .A2(KEYINPUT115), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n802), .A2(new_n810), .A3(new_n812), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT53), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n807), .A2(KEYINPUT52), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n807), .B(new_n814), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n822), .B2(new_n816), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n812), .A4(new_n802), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n820), .A2(new_n825), .A3(KEYINPUT54), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(new_n824), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n800), .A2(new_n699), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT53), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n800), .B2(new_n699), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n799), .B(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n823), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n827), .A2(new_n828), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n788), .A2(new_n789), .A3(new_n826), .A4(new_n837), .ZN(new_n838));
  OR2_X1    g652(.A1(G952), .A2(G953), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n549), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n841), .A2(new_n281), .A3(new_n629), .A4(new_n722), .ZN(new_n842));
  XOR2_X1   g656(.A(new_n842), .B(KEYINPUT111), .Z(new_n843));
  XNOR2_X1  g657(.A(new_n761), .B(KEYINPUT49), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n624), .A3(new_n752), .A4(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT112), .Z(new_n846));
  NAND2_X1  g660(.A1(new_n840), .A2(new_n846), .ZN(G75));
  NAND2_X1  g661(.A1(new_n827), .A2(new_n836), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(G210), .A3(G902), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n250), .B1(new_n257), .B2(new_n260), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(new_n209), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT55), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n849), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n853), .B1(new_n849), .B2(new_n850), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n207), .A2(G952), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(G51));
  NAND2_X1  g671(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n837), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n283), .B(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n318), .A2(new_n330), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n848), .A2(G902), .A3(new_n713), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n856), .B1(new_n863), .B2(new_n864), .ZN(G54));
  AND2_X1   g679(.A1(KEYINPUT58), .A2(G475), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n848), .A2(G902), .A3(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(new_n375), .A2(new_n384), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n856), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n848), .A2(G902), .A3(new_n868), .A4(new_n866), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT122), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n870), .A2(new_n875), .A3(new_n871), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(G60));
  NAND2_X1  g691(.A1(new_n826), .A2(new_n837), .ZN(new_n878));
  NAND2_X1  g692(.A1(G478), .A2(G902), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n565), .A2(new_n566), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n856), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n827), .A2(new_n828), .A3(new_n836), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n828), .B1(new_n827), .B2(new_n836), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n882), .B(new_n880), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n859), .A2(KEYINPUT123), .A3(new_n882), .A4(new_n880), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n884), .A2(new_n889), .A3(new_n890), .ZN(G63));
  NAND2_X1  g705(.A1(G217), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT124), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT60), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n827), .B2(new_n836), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(new_n547), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n589), .A3(new_n590), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(new_n871), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n897), .A2(KEYINPUT61), .A3(new_n871), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(G66));
  INV_X1    g717(.A(new_n798), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n800), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT125), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n906), .A2(G953), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n207), .B1(new_n424), .B2(G224), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT126), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(KEYINPUT126), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n851), .B1(G898), .B2(new_n207), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(G69));
  NAND2_X1  g726(.A1(new_n813), .A2(new_n677), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(new_n705), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n639), .A2(new_n628), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n729), .A2(new_n731), .B1(new_n916), .B2(new_n769), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n699), .B(new_n915), .C1(new_n917), .C2(new_n719), .ZN(new_n918));
  INV_X1    g732(.A(new_n739), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n207), .ZN(new_n920));
  OAI22_X1  g734(.A1(new_n918), .A2(new_n920), .B1(new_n286), .B2(new_n207), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n473), .A2(new_n474), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n381), .B1(new_n348), .B2(new_n380), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n618), .A2(new_n634), .A3(new_n635), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n913), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n914), .A2(KEYINPUT62), .A3(new_n636), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n739), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n617), .A2(new_n702), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n571), .A2(new_n579), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n931), .A2(new_n515), .A3(new_n549), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n732), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n924), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n207), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(G900), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n935), .B2(new_n286), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n925), .B(new_n936), .C1(new_n207), .C2(new_n938), .ZN(G72));
  XOR2_X1   g753(.A(new_n621), .B(KEYINPUT63), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n906), .A2(new_n919), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n918), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n475), .A3(new_n469), .A4(new_n465), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n930), .A2(new_n732), .A3(new_n906), .A4(new_n933), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n940), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n466), .A3(new_n506), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n496), .A2(new_n507), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n820), .A2(new_n825), .A3(new_n940), .A4(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n943), .A2(new_n946), .A3(new_n871), .A4(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n465), .B1(new_n944), .B2(new_n940), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n856), .B1(new_n952), .B2(new_n506), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n953), .A2(KEYINPUT127), .A3(new_n943), .A4(new_n948), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(G57));
endmodule


