

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X4 U553 ( .A1(n724), .A2(n723), .ZN(n745) );
  NAND2_X1 U554 ( .A1(n735), .A2(G8), .ZN(n792) );
  INV_X1 U555 ( .A(n722), .ZN(n724) );
  XNOR2_X1 U556 ( .A(n730), .B(KEYINPUT30), .ZN(n732) );
  INV_X1 U557 ( .A(G168), .ZN(n731) );
  XOR2_X1 U558 ( .A(KEYINPUT31), .B(n734), .Z(n518) );
  AND2_X1 U559 ( .A1(n732), .A2(n731), .ZN(n519) );
  INV_X1 U560 ( .A(KEYINPUT28), .ZN(n756) );
  INV_X1 U561 ( .A(KEYINPUT94), .ZN(n764) );
  NOR2_X1 U562 ( .A1(n792), .A2(n791), .ZN(n793) );
  INV_X1 U563 ( .A(n745), .ZN(n735) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  NOR2_X1 U565 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n654) );
  NOR2_X2 U567 ( .A1(n553), .A2(n552), .ZN(G160) );
  NAND2_X1 U568 ( .A1(G89), .A2(n654), .ZN(n520) );
  XOR2_X1 U569 ( .A(KEYINPUT4), .B(n520), .Z(n521) );
  XNOR2_X1 U570 ( .A(n521), .B(KEYINPUT73), .ZN(n523) );
  XOR2_X1 U571 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  INV_X1 U572 ( .A(G651), .ZN(n526) );
  NOR2_X1 U573 ( .A1(n628), .A2(n526), .ZN(n650) );
  NAND2_X1 U574 ( .A1(G76), .A2(n650), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U576 ( .A(n524), .B(KEYINPUT5), .ZN(n533) );
  NOR2_X2 U577 ( .A1(G651), .A2(n628), .ZN(n653) );
  NAND2_X1 U578 ( .A1(n653), .A2(G51), .ZN(n525) );
  XNOR2_X1 U579 ( .A(n525), .B(KEYINPUT74), .ZN(n530) );
  NOR2_X1 U580 ( .A1(G543), .A2(n526), .ZN(n528) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n527) );
  XNOR2_X1 U582 ( .A(n528), .B(n527), .ZN(n657) );
  NAND2_X1 U583 ( .A1(G63), .A2(n657), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U585 ( .A(KEYINPUT6), .B(n531), .Z(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 U588 ( .A(G2104), .ZN(n540) );
  NOR2_X4 U589 ( .A1(G2105), .A2(n540), .ZN(n888) );
  NAND2_X1 U590 ( .A1(n888), .A2(G102), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT17), .B(n535), .Z(n536) );
  XNOR2_X2 U592 ( .A(n536), .B(KEYINPUT66), .ZN(n885) );
  NAND2_X1 U593 ( .A1(G138), .A2(n885), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n539), .B(KEYINPUT65), .ZN(n880) );
  NAND2_X1 U597 ( .A1(G114), .A2(n880), .ZN(n542) );
  AND2_X1 U598 ( .A1(n540), .A2(G2105), .ZN(n881) );
  NAND2_X1 U599 ( .A1(G126), .A2(n881), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U601 ( .A1(n544), .A2(n543), .ZN(G164) );
  XOR2_X1 U602 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U603 ( .A(KEYINPUT23), .ZN(n546) );
  NAND2_X1 U604 ( .A1(G101), .A2(n888), .ZN(n545) );
  XNOR2_X1 U605 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U606 ( .A(n547), .B(KEYINPUT64), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G137), .A2(n885), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G113), .A2(n880), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G125), .A2(n881), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U612 ( .A(G2443), .B(G2446), .Z(n555) );
  XNOR2_X1 U613 ( .A(G2427), .B(G2451), .ZN(n554) );
  XNOR2_X1 U614 ( .A(n555), .B(n554), .ZN(n561) );
  XOR2_X1 U615 ( .A(G2430), .B(G2454), .Z(n557) );
  XNOR2_X1 U616 ( .A(G1341), .B(G1348), .ZN(n556) );
  XNOR2_X1 U617 ( .A(n557), .B(n556), .ZN(n559) );
  XOR2_X1 U618 ( .A(G2435), .B(G2438), .Z(n558) );
  XNOR2_X1 U619 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U620 ( .A(n561), .B(n560), .Z(n562) );
  AND2_X1 U621 ( .A1(G14), .A2(n562), .ZN(G401) );
  AND2_X1 U622 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  INV_X1 U625 ( .A(G120), .ZN(G236) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U628 ( .A(G223), .ZN(n823) );
  NAND2_X1 U629 ( .A1(n823), .A2(G567), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U631 ( .A1(G56), .A2(n657), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n565), .Z(n572) );
  NAND2_X1 U633 ( .A1(n650), .A2(G68), .ZN(n566) );
  XNOR2_X1 U634 ( .A(KEYINPUT71), .B(n566), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n654), .A2(G81), .ZN(n567) );
  XOR2_X1 U636 ( .A(KEYINPUT12), .B(n567), .Z(n568) );
  NOR2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n570), .B(KEYINPUT13), .ZN(n571) );
  NOR2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n653), .A2(G43), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n1003) );
  INV_X1 U642 ( .A(G860), .ZN(n618) );
  OR2_X1 U643 ( .A1(n1003), .A2(n618), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G77), .A2(n650), .ZN(n576) );
  NAND2_X1 U645 ( .A1(G90), .A2(n654), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U647 ( .A(KEYINPUT9), .B(n577), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n653), .A2(G52), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G64), .A2(n657), .ZN(n578) );
  AND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(G301) );
  NAND2_X1 U652 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U653 ( .A1(n657), .A2(G66), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G79), .A2(n650), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G92), .A2(n654), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n653), .A2(G54), .ZN(n584) );
  XOR2_X1 U658 ( .A(KEYINPUT72), .B(n584), .Z(n585) );
  NOR2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U661 ( .A(KEYINPUT15), .B(n589), .Z(n991) );
  INV_X1 U662 ( .A(G868), .ZN(n674) );
  NAND2_X1 U663 ( .A1(n991), .A2(n674), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U665 ( .A1(G53), .A2(n653), .ZN(n593) );
  NAND2_X1 U666 ( .A1(G65), .A2(n657), .ZN(n592) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G78), .A2(n650), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G91), .A2(n654), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n995) );
  XOR2_X1 U672 ( .A(n995), .B(KEYINPUT70), .Z(G299) );
  NOR2_X1 U673 ( .A1(G299), .A2(G868), .ZN(n599) );
  NOR2_X1 U674 ( .A1(G286), .A2(n674), .ZN(n598) );
  NOR2_X1 U675 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n618), .A2(G559), .ZN(n600) );
  INV_X1 U677 ( .A(n991), .ZN(n616) );
  NAND2_X1 U678 ( .A1(n600), .A2(n616), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n601), .B(KEYINPUT75), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT16), .B(n602), .Z(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n1003), .ZN(n605) );
  NAND2_X1 U682 ( .A1(G868), .A2(n616), .ZN(n603) );
  NOR2_X1 U683 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U684 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G111), .A2(n880), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n888), .A2(G99), .ZN(n607) );
  NAND2_X1 U687 ( .A1(G135), .A2(n885), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n881), .A2(G123), .ZN(n608) );
  XOR2_X1 U690 ( .A(KEYINPUT18), .B(n608), .Z(n609) );
  NOR2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U693 ( .A(n613), .B(KEYINPUT76), .ZN(n964) );
  XOR2_X1 U694 ( .A(n964), .B(G2096), .Z(n615) );
  XNOR2_X1 U695 ( .A(G2100), .B(KEYINPUT77), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U697 ( .A1(G559), .A2(n616), .ZN(n617) );
  XOR2_X1 U698 ( .A(n1003), .B(n617), .Z(n670) );
  NAND2_X1 U699 ( .A1(n618), .A2(n670), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G80), .A2(n650), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n619), .B(KEYINPUT78), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G67), .A2(n657), .ZN(n621) );
  NAND2_X1 U703 ( .A1(G93), .A2(n654), .ZN(n620) );
  NAND2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U705 ( .A1(G55), .A2(n653), .ZN(n622) );
  XNOR2_X1 U706 ( .A(KEYINPUT79), .B(n622), .ZN(n623) );
  NOR2_X1 U707 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n673) );
  XNOR2_X1 U709 ( .A(n627), .B(n673), .ZN(G145) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G49), .A2(n653), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G87), .A2(n628), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n657), .A2(n631), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U716 ( .A(n634), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U717 ( .A1(n653), .A2(G47), .ZN(n635) );
  XNOR2_X1 U718 ( .A(n635), .B(KEYINPUT68), .ZN(n637) );
  NAND2_X1 U719 ( .A1(G60), .A2(n657), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U721 ( .A(KEYINPUT69), .B(n638), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G72), .A2(n650), .ZN(n640) );
  NAND2_X1 U723 ( .A1(G85), .A2(n654), .ZN(n639) );
  AND2_X1 U724 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U726 ( .A1(G50), .A2(n653), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G62), .A2(n657), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U729 ( .A(KEYINPUT83), .B(n645), .ZN(n649) );
  NAND2_X1 U730 ( .A1(G75), .A2(n650), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G88), .A2(n654), .ZN(n646) );
  AND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(G303) );
  INV_X1 U734 ( .A(G303), .ZN(G166) );
  NAND2_X1 U735 ( .A1(n650), .A2(G73), .ZN(n652) );
  XNOR2_X1 U736 ( .A(KEYINPUT2), .B(KEYINPUT82), .ZN(n651) );
  XNOR2_X1 U737 ( .A(n652), .B(n651), .ZN(n662) );
  NAND2_X1 U738 ( .A1(G48), .A2(n653), .ZN(n656) );
  NAND2_X1 U739 ( .A1(G86), .A2(n654), .ZN(n655) );
  NAND2_X1 U740 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U741 ( .A1(G61), .A2(n657), .ZN(n658) );
  XNOR2_X1 U742 ( .A(KEYINPUT81), .B(n658), .ZN(n659) );
  NOR2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U744 ( .A1(n662), .A2(n661), .ZN(G305) );
  XOR2_X1 U745 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n664) );
  XNOR2_X1 U746 ( .A(G288), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U747 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U748 ( .A(G299), .B(n665), .ZN(n667) );
  XNOR2_X1 U749 ( .A(G290), .B(G166), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U751 ( .A(n668), .B(G305), .Z(n669) );
  XNOR2_X1 U752 ( .A(n673), .B(n669), .ZN(n896) );
  XNOR2_X1 U753 ( .A(n670), .B(n896), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n671), .A2(G868), .ZN(n672) );
  XNOR2_X1 U755 ( .A(n672), .B(KEYINPUT86), .ZN(n676) );
  NAND2_X1 U756 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U757 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2084), .A2(G2078), .ZN(n677) );
  XNOR2_X1 U759 ( .A(n677), .B(KEYINPUT20), .ZN(n678) );
  XNOR2_X1 U760 ( .A(n678), .B(KEYINPUT87), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n679), .A2(G2090), .ZN(n680) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U763 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U765 ( .A1(G69), .A2(G57), .ZN(n682) );
  NOR2_X1 U766 ( .A1(G236), .A2(n682), .ZN(n683) );
  XNOR2_X1 U767 ( .A(KEYINPUT88), .B(n683), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n684), .A2(G108), .ZN(n829) );
  NAND2_X1 U769 ( .A1(G567), .A2(n829), .ZN(n689) );
  NOR2_X1 U770 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U772 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U773 ( .A1(G96), .A2(n687), .ZN(n828) );
  NAND2_X1 U774 ( .A1(G2106), .A2(n828), .ZN(n688) );
  NAND2_X1 U775 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U776 ( .A(KEYINPUT89), .B(n690), .ZN(G319) );
  INV_X1 U777 ( .A(G319), .ZN(n692) );
  NAND2_X1 U778 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n825) );
  NAND2_X1 U780 ( .A1(n825), .A2(G36), .ZN(G176) );
  XNOR2_X1 U781 ( .A(G1986), .B(KEYINPUT90), .ZN(n693) );
  XNOR2_X1 U782 ( .A(n693), .B(G290), .ZN(n1009) );
  NOR2_X2 U783 ( .A1(G164), .A2(G1384), .ZN(n722) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n723) );
  NOR2_X1 U785 ( .A1(n722), .A2(n723), .ZN(n818) );
  NAND2_X1 U786 ( .A1(n1009), .A2(n818), .ZN(n807) );
  XOR2_X1 U787 ( .A(G2067), .B(KEYINPUT37), .Z(n815) );
  NAND2_X1 U788 ( .A1(G116), .A2(n880), .ZN(n695) );
  NAND2_X1 U789 ( .A1(G128), .A2(n881), .ZN(n694) );
  NAND2_X1 U790 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U791 ( .A(n696), .B(KEYINPUT35), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n888), .A2(G104), .ZN(n698) );
  NAND2_X1 U793 ( .A1(G140), .A2(n885), .ZN(n697) );
  NAND2_X1 U794 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U795 ( .A(KEYINPUT34), .B(n699), .Z(n700) );
  NAND2_X1 U796 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U797 ( .A(n702), .B(KEYINPUT36), .ZN(n892) );
  NAND2_X1 U798 ( .A1(n815), .A2(n892), .ZN(n703) );
  XNOR2_X1 U799 ( .A(n703), .B(KEYINPUT91), .ZN(n982) );
  NAND2_X1 U800 ( .A1(n818), .A2(n982), .ZN(n813) );
  NAND2_X1 U801 ( .A1(n888), .A2(G95), .ZN(n705) );
  NAND2_X1 U802 ( .A1(G131), .A2(n885), .ZN(n704) );
  NAND2_X1 U803 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U804 ( .A1(G107), .A2(n880), .ZN(n707) );
  NAND2_X1 U805 ( .A1(G119), .A2(n881), .ZN(n706) );
  NAND2_X1 U806 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X1 U807 ( .A1(n709), .A2(n708), .ZN(n858) );
  AND2_X1 U808 ( .A1(n858), .A2(G1991), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n880), .A2(G117), .ZN(n711) );
  NAND2_X1 U810 ( .A1(G141), .A2(n885), .ZN(n710) );
  NAND2_X1 U811 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n888), .A2(G105), .ZN(n712) );
  XOR2_X1 U813 ( .A(KEYINPUT38), .B(n712), .Z(n713) );
  NOR2_X1 U814 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n881), .A2(G129), .ZN(n715) );
  NAND2_X1 U816 ( .A1(n716), .A2(n715), .ZN(n876) );
  AND2_X1 U817 ( .A1(G1996), .A2(n876), .ZN(n717) );
  NOR2_X1 U818 ( .A1(n718), .A2(n717), .ZN(n972) );
  INV_X1 U819 ( .A(n818), .ZN(n719) );
  NOR2_X1 U820 ( .A1(n972), .A2(n719), .ZN(n810) );
  INV_X1 U821 ( .A(n810), .ZN(n720) );
  NAND2_X1 U822 ( .A1(n813), .A2(n720), .ZN(n805) );
  NOR2_X1 U823 ( .A1(G1981), .A2(G305), .ZN(n721) );
  XNOR2_X1 U824 ( .A(KEYINPUT24), .B(n721), .ZN(n725) );
  INV_X1 U825 ( .A(n792), .ZN(n795) );
  NAND2_X1 U826 ( .A1(n725), .A2(n795), .ZN(n787) );
  XOR2_X1 U827 ( .A(G2078), .B(KEYINPUT25), .Z(n914) );
  INV_X1 U828 ( .A(n745), .ZN(n767) );
  NOR2_X1 U829 ( .A1(n914), .A2(n767), .ZN(n727) );
  NOR2_X1 U830 ( .A1(n745), .A2(G1961), .ZN(n726) );
  NOR2_X1 U831 ( .A1(n727), .A2(n726), .ZN(n761) );
  AND2_X1 U832 ( .A1(G301), .A2(n761), .ZN(n733) );
  NOR2_X1 U833 ( .A1(G1966), .A2(n792), .ZN(n778) );
  NOR2_X1 U834 ( .A1(G2084), .A2(n767), .ZN(n775) );
  NOR2_X1 U835 ( .A1(n778), .A2(n775), .ZN(n728) );
  NAND2_X1 U836 ( .A1(G8), .A2(n728), .ZN(n729) );
  XNOR2_X1 U837 ( .A(KEYINPUT95), .B(n729), .ZN(n730) );
  NOR2_X1 U838 ( .A1(n733), .A2(n519), .ZN(n734) );
  NAND2_X1 U839 ( .A1(G1956), .A2(n735), .ZN(n736) );
  XNOR2_X1 U840 ( .A(n736), .B(KEYINPUT93), .ZN(n740) );
  XOR2_X1 U841 ( .A(KEYINPUT92), .B(KEYINPUT27), .Z(n738) );
  AND2_X1 U842 ( .A1(n745), .A2(G2072), .ZN(n737) );
  XNOR2_X1 U843 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U844 ( .A1(n740), .A2(n739), .ZN(n755) );
  NAND2_X1 U845 ( .A1(n995), .A2(n755), .ZN(n754) );
  AND2_X1 U846 ( .A1(n745), .A2(G1996), .ZN(n741) );
  XOR2_X1 U847 ( .A(n741), .B(KEYINPUT26), .Z(n743) );
  NAND2_X1 U848 ( .A1(n767), .A2(G1341), .ZN(n742) );
  NAND2_X1 U849 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U850 ( .A1(n1003), .A2(n744), .ZN(n749) );
  NAND2_X1 U851 ( .A1(G1348), .A2(n767), .ZN(n747) );
  NAND2_X1 U852 ( .A1(G2067), .A2(n745), .ZN(n746) );
  NAND2_X1 U853 ( .A1(n747), .A2(n746), .ZN(n750) );
  NOR2_X1 U854 ( .A1(n991), .A2(n750), .ZN(n748) );
  OR2_X1 U855 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U856 ( .A1(n991), .A2(n750), .ZN(n751) );
  NAND2_X1 U857 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U858 ( .A1(n754), .A2(n753), .ZN(n759) );
  NOR2_X1 U859 ( .A1(n995), .A2(n755), .ZN(n757) );
  XNOR2_X1 U860 ( .A(n757), .B(n756), .ZN(n758) );
  NAND2_X1 U861 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U862 ( .A(n760), .B(KEYINPUT29), .ZN(n763) );
  NOR2_X1 U863 ( .A1(G301), .A2(n761), .ZN(n762) );
  NOR2_X1 U864 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U865 ( .A(n765), .B(n764), .ZN(n766) );
  NAND2_X1 U866 ( .A1(n518), .A2(n766), .ZN(n776) );
  NAND2_X1 U867 ( .A1(n776), .A2(G286), .ZN(n772) );
  NOR2_X1 U868 ( .A1(G1971), .A2(n792), .ZN(n769) );
  NOR2_X1 U869 ( .A1(G2090), .A2(n767), .ZN(n768) );
  NOR2_X1 U870 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U871 ( .A1(n770), .A2(G303), .ZN(n771) );
  NAND2_X1 U872 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U873 ( .A1(n773), .A2(G8), .ZN(n774) );
  XNOR2_X1 U874 ( .A(n774), .B(KEYINPUT32), .ZN(n782) );
  NAND2_X1 U875 ( .A1(G8), .A2(n775), .ZN(n780) );
  INV_X1 U876 ( .A(n776), .ZN(n777) );
  NOR2_X1 U877 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n789) );
  NOR2_X1 U880 ( .A1(G2090), .A2(G303), .ZN(n783) );
  NAND2_X1 U881 ( .A1(G8), .A2(n783), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n789), .A2(n784), .ZN(n785) );
  NAND2_X1 U883 ( .A1(n792), .A2(n785), .ZN(n786) );
  NAND2_X1 U884 ( .A1(n787), .A2(n786), .ZN(n803) );
  XNOR2_X1 U885 ( .A(G1981), .B(G305), .ZN(n1012) );
  NOR2_X1 U886 ( .A1(G1976), .A2(G288), .ZN(n992) );
  INV_X1 U887 ( .A(G1971), .ZN(n947) );
  NAND2_X1 U888 ( .A1(G166), .A2(n947), .ZN(n788) );
  NAND2_X1 U889 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U890 ( .A1(n992), .A2(n790), .ZN(n791) );
  NAND2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n997) );
  NAND2_X1 U892 ( .A1(n793), .A2(n997), .ZN(n794) );
  INV_X1 U893 ( .A(KEYINPUT33), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n794), .A2(n797), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n795), .A2(n992), .ZN(n796) );
  NOR2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U897 ( .A(n798), .B(KEYINPUT96), .Z(n799) );
  NAND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U899 ( .A1(n1012), .A2(n801), .ZN(n802) );
  NOR2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n821) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n876), .ZN(n974) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n858), .ZN(n962) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n962), .A2(n808), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U907 ( .A1(n974), .A2(n811), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n815), .A2(n892), .ZN(n816) );
  XNOR2_X1 U911 ( .A(n816), .B(KEYINPUT97), .ZN(n979) );
  NAND2_X1 U912 ( .A1(n817), .A2(n979), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G1), .A2(G3), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n827), .B(KEYINPUT98), .ZN(G188) );
  XNOR2_X1 U922 ( .A(G69), .B(KEYINPUT99), .ZN(G235) );
  XNOR2_X1 U923 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G57), .ZN(G237) );
  NOR2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n830), .B(KEYINPUT100), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XOR2_X1 U930 ( .A(G2096), .B(G2100), .Z(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(KEYINPUT43), .B(G2090), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2072), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2084), .B(G2078), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(G227) );
  XOR2_X1 U939 ( .A(KEYINPUT102), .B(G1976), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1956), .B(G1981), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G1971), .B(G1961), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1966), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U948 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT101), .B(G2474), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U951 ( .A1(G100), .A2(n888), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G112), .A2(n880), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n857) );
  NAND2_X1 U954 ( .A1(n881), .A2(G124), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U956 ( .A1(G136), .A2(n885), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U958 ( .A(KEYINPUT103), .B(n855), .Z(n856) );
  NOR2_X1 U959 ( .A1(n857), .A2(n856), .ZN(G162) );
  XOR2_X1 U960 ( .A(G160), .B(n858), .Z(n865) );
  XOR2_X1 U961 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n860) );
  XNOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U964 ( .A(n861), .B(KEYINPUT109), .Z(n863) );
  XNOR2_X1 U965 ( .A(G162), .B(KEYINPUT48), .ZN(n862) );
  XNOR2_X1 U966 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n875) );
  NAND2_X1 U968 ( .A1(G118), .A2(n880), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G130), .A2(n881), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n888), .A2(G106), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G142), .A2(n885), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n870), .Z(n871) );
  XNOR2_X1 U975 ( .A(KEYINPUT104), .B(n871), .ZN(n872) );
  NOR2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U977 ( .A(n875), .B(n874), .Z(n878) );
  XOR2_X1 U978 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U980 ( .A(n879), .B(n964), .Z(n894) );
  NAND2_X1 U981 ( .A1(G115), .A2(n880), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G127), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n884), .B(KEYINPUT47), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G139), .A2(n885), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G103), .A2(n888), .ZN(n889) );
  XNOR2_X1 U988 ( .A(KEYINPUT105), .B(n889), .ZN(n890) );
  NOR2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n965) );
  XNOR2_X1 U990 ( .A(n892), .B(n965), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(G395) );
  INV_X1 U993 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U994 ( .A(G286), .B(n1003), .ZN(n897) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U996 ( .A(n991), .B(G171), .Z(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U998 ( .A1(G37), .A2(n900), .ZN(n901) );
  XNOR2_X1 U999 ( .A(KEYINPUT110), .B(n901), .ZN(G397) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(n902), .B(KEYINPUT49), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(G401), .A2(n903), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n904), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(KEYINPUT111), .B(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(KEYINPUT112), .B(n908), .Z(G308) );
  INV_X1 U1008 ( .A(G308), .ZN(G225) );
  INV_X1 U1009 ( .A(KEYINPUT55), .ZN(n984) );
  XNOR2_X1 U1010 ( .A(KEYINPUT115), .B(G2090), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(n909), .B(G35), .ZN(n928) );
  XNOR2_X1 U1012 ( .A(G2084), .B(G34), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(n910), .B(KEYINPUT54), .ZN(n926) );
  XOR2_X1 U1014 ( .A(G1991), .B(G25), .Z(n911) );
  NAND2_X1 U1015 ( .A1(n911), .A2(G28), .ZN(n912) );
  XNOR2_X1 U1016 ( .A(n912), .B(KEYINPUT116), .ZN(n923) );
  INV_X1 U1017 ( .A(G1996), .ZN(n913) );
  XNOR2_X1 U1018 ( .A(G32), .B(n913), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n914), .B(G27), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(G2067), .B(G26), .ZN(n916) );
  XNOR2_X1 U1021 ( .A(G2072), .B(G33), .ZN(n915) );
  NOR2_X1 U1022 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1023 ( .A(KEYINPUT117), .B(n917), .ZN(n918) );
  NOR2_X1 U1024 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1027 ( .A(n924), .B(KEYINPUT53), .ZN(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(n984), .B(n929), .ZN(n931) );
  INV_X1 U1031 ( .A(G29), .ZN(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1033 ( .A1(G11), .A2(n932), .ZN(n960) );
  XOR2_X1 U1034 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n957) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G21), .ZN(n934) );
  XNOR2_X1 U1036 ( .A(G5), .B(G1961), .ZN(n933) );
  NOR2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n955) );
  XOR2_X1 U1038 ( .A(G1341), .B(G19), .Z(n938) );
  XNOR2_X1 U1039 ( .A(G1956), .B(G20), .ZN(n936) );
  XNOR2_X1 U1040 ( .A(G1981), .B(G6), .ZN(n935) );
  NOR2_X1 U1041 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1042 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1043 ( .A(KEYINPUT124), .B(n939), .ZN(n942) );
  XOR2_X1 U1044 ( .A(KEYINPUT59), .B(G1348), .Z(n940) );
  XNOR2_X1 U1045 ( .A(G4), .B(n940), .ZN(n941) );
  NOR2_X1 U1046 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1047 ( .A(n943), .B(KEYINPUT125), .ZN(n944) );
  XNOR2_X1 U1048 ( .A(n944), .B(KEYINPUT60), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(G1986), .B(G24), .ZN(n946) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n945) );
  NOR2_X1 U1051 ( .A1(n946), .A2(n945), .ZN(n950) );
  XNOR2_X1 U1052 ( .A(G22), .B(KEYINPUT126), .ZN(n948) );
  XNOR2_X1 U1053 ( .A(n948), .B(n947), .ZN(n949) );
  NAND2_X1 U1054 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1055 ( .A(KEYINPUT58), .B(n951), .ZN(n952) );
  NOR2_X1 U1056 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1058 ( .A(n957), .B(n956), .ZN(n958) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n958), .ZN(n959) );
  NOR2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n988) );
  XOR2_X1 U1061 ( .A(G160), .B(G2084), .Z(n961) );
  NOR2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n970) );
  XOR2_X1 U1064 ( .A(G2072), .B(n965), .Z(n967) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n966) );
  NOR2_X1 U1066 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1067 ( .A(KEYINPUT50), .B(n968), .Z(n969) );
  NOR2_X1 U1068 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n978) );
  XOR2_X1 U1070 ( .A(G2090), .B(G162), .Z(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT51), .B(n975), .ZN(n976) );
  XNOR2_X1 U1073 ( .A(KEYINPUT114), .B(n976), .ZN(n977) );
  NOR2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n986), .A2(G29), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(G16), .B(KEYINPUT118), .Z(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT56), .B(n989), .ZN(n1018) );
  XOR2_X1 U1083 ( .A(G1348), .B(KEYINPUT119), .Z(n990) );
  XNOR2_X1 U1084 ( .A(n991), .B(n990), .ZN(n994) );
  XOR2_X1 U1085 ( .A(n992), .B(KEYINPUT121), .Z(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n1007) );
  XNOR2_X1 U1087 ( .A(G166), .B(G1971), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(n995), .B(G1956), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(n996), .B(KEYINPUT120), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G1961), .B(G301), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(G1341), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(KEYINPUT122), .B(n1010), .Z(n1015) );
  XOR2_X1 U1099 ( .A(G1966), .B(G168), .Z(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT57), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT123), .B(n1016), .Z(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

