

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(G2105), .A2(n527), .ZN(n996) );
  NOR2_X2 U555 ( .A1(n531), .A2(n530), .ZN(G160) );
  OR2_X1 U556 ( .A1(n968), .A2(n610), .ZN(n520) );
  OR2_X1 U557 ( .A1(n965), .A2(n620), .ZN(n521) );
  NOR2_X1 U558 ( .A1(n711), .A2(n682), .ZN(n522) );
  OR2_X1 U559 ( .A1(n630), .A2(KEYINPUT27), .ZN(n631) );
  XNOR2_X1 U560 ( .A(KEYINPUT30), .B(KEYINPUT96), .ZN(n648) );
  XNOR2_X1 U561 ( .A(n649), .B(n648), .ZN(n650) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n654) );
  INV_X1 U563 ( .A(KEYINPUT97), .ZN(n658) );
  AND2_X1 U564 ( .A1(G160), .A2(G40), .ZN(n589) );
  XNOR2_X1 U565 ( .A(n590), .B(KEYINPUT64), .ZN(n606) );
  NOR2_X1 U566 ( .A1(G164), .A2(G1384), .ZN(n691) );
  NOR2_X1 U567 ( .A1(G651), .A2(n572), .ZN(n804) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n800) );
  XOR2_X1 U569 ( .A(KEYINPUT17), .B(n523), .Z(n995) );
  INV_X1 U570 ( .A(KEYINPUT40), .ZN(n757) );
  XOR2_X1 U571 ( .A(KEYINPUT70), .B(n605), .Z(n968) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NAND2_X1 U573 ( .A1(G137), .A2(n995), .ZN(n525) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n992) );
  NAND2_X1 U575 ( .A1(G113), .A2(n992), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n531) );
  XNOR2_X1 U577 ( .A(G2104), .B(KEYINPUT65), .ZN(n527) );
  NAND2_X1 U578 ( .A1(G101), .A2(n996), .ZN(n526) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n526), .Z(n529) );
  AND2_X1 U580 ( .A1(n527), .A2(G2105), .ZN(n991) );
  NAND2_X1 U581 ( .A1(n991), .A2(G125), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G138), .A2(n995), .ZN(n533) );
  NAND2_X1 U584 ( .A1(G126), .A2(n991), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n539) );
  NAND2_X1 U586 ( .A1(G102), .A2(n996), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT84), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G114), .A2(n992), .ZN(n535) );
  XOR2_X1 U589 ( .A(KEYINPUT83), .B(n535), .Z(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n539), .A2(n538), .ZN(G164) );
  XOR2_X1 U592 ( .A(G543), .B(KEYINPUT0), .Z(n572) );
  NAND2_X1 U593 ( .A1(G52), .A2(n804), .ZN(n542) );
  INV_X1 U594 ( .A(G651), .ZN(n544) );
  NOR2_X1 U595 ( .A1(G543), .A2(n544), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n540), .Z(n805) );
  NAND2_X1 U597 ( .A1(G64), .A2(n805), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n542), .A2(n541), .ZN(n549) );
  NAND2_X1 U599 ( .A1(n800), .A2(G90), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT67), .B(n543), .Z(n546) );
  NOR2_X1 U601 ( .A1(n572), .A2(n544), .ZN(n801) );
  NAND2_X1 U602 ( .A1(n801), .A2(G77), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U605 ( .A1(n549), .A2(n548), .ZN(G171) );
  INV_X1 U606 ( .A(G171), .ZN(G301) );
  NAND2_X1 U607 ( .A1(n800), .A2(G89), .ZN(n550) );
  XNOR2_X1 U608 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G76), .A2(n801), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U611 ( .A(n553), .B(KEYINPUT5), .ZN(n559) );
  XNOR2_X1 U612 ( .A(KEYINPUT71), .B(KEYINPUT6), .ZN(n557) );
  NAND2_X1 U613 ( .A1(G51), .A2(n804), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G63), .A2(n805), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U618 ( .A(KEYINPUT7), .B(n560), .ZN(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(n561) );
  XNOR2_X1 U620 ( .A(KEYINPUT72), .B(n561), .ZN(G286) );
  NAND2_X1 U621 ( .A1(n800), .A2(G88), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G75), .A2(n801), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT79), .B(n562), .Z(n563) );
  NAND2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U625 ( .A1(G50), .A2(n804), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G62), .A2(n805), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U628 ( .A1(n568), .A2(n567), .ZN(G166) );
  XNOR2_X1 U629 ( .A(G166), .B(KEYINPUT85), .ZN(G303) );
  NAND2_X1 U630 ( .A1(G49), .A2(n804), .ZN(n570) );
  NAND2_X1 U631 ( .A1(G74), .A2(G651), .ZN(n569) );
  NAND2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n805), .A2(n571), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n572), .A2(G87), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(G288) );
  NAND2_X1 U636 ( .A1(G48), .A2(n804), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G86), .A2(n800), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n801), .A2(G73), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT2), .B(n577), .Z(n578) );
  NOR2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n805), .A2(G61), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(G305) );
  NAND2_X1 U644 ( .A1(G47), .A2(n804), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G60), .A2(n805), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT66), .B(n584), .Z(n588) );
  NAND2_X1 U648 ( .A1(G85), .A2(n800), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G72), .A2(n801), .ZN(n585) );
  AND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(G290) );
  XOR2_X1 U652 ( .A(G1961), .B(KEYINPUT91), .Z(n905) );
  NAND2_X1 U653 ( .A1(n589), .A2(n691), .ZN(n590) );
  BUF_X2 U654 ( .A(n606), .Z(n660) );
  INV_X1 U655 ( .A(n660), .ZN(n633) );
  NOR2_X1 U656 ( .A1(n905), .A2(n633), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n591), .B(KEYINPUT92), .ZN(n593) );
  XOR2_X1 U658 ( .A(G2078), .B(KEYINPUT25), .Z(n881) );
  NOR2_X1 U659 ( .A1(n660), .A2(n881), .ZN(n592) );
  NOR2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U661 ( .A(KEYINPUT93), .B(n594), .Z(n651) );
  NOR2_X1 U662 ( .A1(n651), .A2(G301), .ZN(n645) );
  NAND2_X1 U663 ( .A1(G81), .A2(n800), .ZN(n595) );
  XOR2_X1 U664 ( .A(KEYINPUT69), .B(n595), .Z(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT12), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G68), .A2(n801), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U668 ( .A(n599), .B(KEYINPUT13), .ZN(n601) );
  NAND2_X1 U669 ( .A1(G43), .A2(n804), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U671 ( .A1(n805), .A2(G56), .ZN(n602) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n602), .Z(n603) );
  NOR2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n605) );
  INV_X1 U674 ( .A(n606), .ZN(n629) );
  NAND2_X1 U675 ( .A1(n629), .A2(G1996), .ZN(n607) );
  XNOR2_X1 U676 ( .A(n607), .B(KEYINPUT26), .ZN(n609) );
  NAND2_X1 U677 ( .A1(n660), .A2(G1341), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n609), .A2(n608), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G54), .A2(n804), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G66), .A2(n805), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U682 ( .A1(G92), .A2(n800), .ZN(n614) );
  NAND2_X1 U683 ( .A1(G79), .A2(n801), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U686 ( .A(n617), .B(KEYINPUT15), .ZN(n965) );
  NAND2_X1 U687 ( .A1(G2067), .A2(n633), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n660), .A2(G1348), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n520), .A2(n521), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n965), .A2(n620), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n637) );
  NAND2_X1 U693 ( .A1(G53), .A2(n804), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G65), .A2(n805), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U696 ( .A1(G91), .A2(n800), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G78), .A2(n801), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n851) );
  NAND2_X1 U700 ( .A1(G2072), .A2(n629), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n630), .A2(KEYINPUT27), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n635) );
  INV_X1 U703 ( .A(G1956), .ZN(n897) );
  NOR2_X1 U704 ( .A1(n633), .A2(n897), .ZN(n634) );
  NOR2_X1 U705 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U706 ( .A1(n851), .A2(n638), .ZN(n636) );
  NAND2_X1 U707 ( .A1(n637), .A2(n636), .ZN(n641) );
  NOR2_X1 U708 ( .A1(n638), .A2(n851), .ZN(n639) );
  XOR2_X1 U709 ( .A(n639), .B(KEYINPUT28), .Z(n640) );
  NAND2_X1 U710 ( .A1(n641), .A2(n640), .ZN(n643) );
  XNOR2_X1 U711 ( .A(KEYINPUT29), .B(KEYINPUT94), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(n644) );
  NOR2_X1 U713 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U714 ( .A(n646), .B(KEYINPUT95), .ZN(n657) );
  NAND2_X1 U715 ( .A1(n660), .A2(G8), .ZN(n711) );
  NOR2_X1 U716 ( .A1(G1966), .A2(n711), .ZN(n671) );
  NOR2_X1 U717 ( .A1(n660), .A2(G2084), .ZN(n668) );
  NOR2_X1 U718 ( .A1(n671), .A2(n668), .ZN(n647) );
  NAND2_X1 U719 ( .A1(G8), .A2(n647), .ZN(n649) );
  NOR2_X1 U720 ( .A1(G168), .A2(n650), .ZN(n653) );
  AND2_X1 U721 ( .A1(G301), .A2(n651), .ZN(n652) );
  NOR2_X1 U722 ( .A1(n653), .A2(n652), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n669) );
  NAND2_X1 U725 ( .A1(n669), .A2(G286), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n659), .B(n658), .ZN(n665) );
  NOR2_X1 U727 ( .A1(n660), .A2(G2090), .ZN(n662) );
  NOR2_X1 U728 ( .A1(G1971), .A2(n711), .ZN(n661) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U730 ( .A1(G303), .A2(n663), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n666), .A2(G8), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(KEYINPUT32), .ZN(n675) );
  NAND2_X1 U734 ( .A1(G8), .A2(n668), .ZN(n673) );
  INV_X1 U735 ( .A(n669), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n706) );
  NOR2_X1 U739 ( .A1(G288), .A2(G1976), .ZN(n676) );
  XNOR2_X1 U740 ( .A(n676), .B(KEYINPUT98), .ZN(n683) );
  NOR2_X1 U741 ( .A1(G1971), .A2(G303), .ZN(n677) );
  OR2_X1 U742 ( .A1(n683), .A2(n677), .ZN(n859) );
  XNOR2_X1 U743 ( .A(n859), .B(KEYINPUT99), .ZN(n678) );
  NAND2_X1 U744 ( .A1(n706), .A2(n678), .ZN(n680) );
  INV_X1 U745 ( .A(KEYINPUT100), .ZN(n682) );
  NAND2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n857) );
  AND2_X1 U747 ( .A1(n522), .A2(n857), .ZN(n679) );
  AND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U749 ( .A1(KEYINPUT33), .A2(n681), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n682), .A2(n683), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n683), .A2(KEYINPUT33), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n684), .A2(KEYINPUT100), .ZN(n685) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U754 ( .A1(n711), .A2(n687), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n703) );
  XOR2_X1 U756 ( .A(G1981), .B(G305), .Z(n863) );
  NAND2_X1 U757 ( .A1(G160), .A2(G40), .ZN(n690) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n751) );
  NAND2_X1 U759 ( .A1(G140), .A2(n995), .ZN(n693) );
  NAND2_X1 U760 ( .A1(G104), .A2(n996), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n695) );
  XOR2_X1 U762 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n694) );
  XNOR2_X1 U763 ( .A(n695), .B(n694), .ZN(n700) );
  NAND2_X1 U764 ( .A1(G128), .A2(n991), .ZN(n697) );
  NAND2_X1 U765 ( .A1(G116), .A2(n992), .ZN(n696) );
  NAND2_X1 U766 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U767 ( .A(KEYINPUT35), .B(n698), .Z(n699) );
  NOR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(KEYINPUT36), .B(n701), .ZN(n1016) );
  XNOR2_X1 U770 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  NOR2_X1 U771 ( .A1(n1016), .A2(n742), .ZN(n921) );
  NAND2_X1 U772 ( .A1(n751), .A2(n921), .ZN(n739) );
  AND2_X1 U773 ( .A1(n863), .A2(n739), .ZN(n702) );
  NAND2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n747) );
  NOR2_X1 U775 ( .A1(G2090), .A2(G303), .ZN(n704) );
  NAND2_X1 U776 ( .A1(G8), .A2(n704), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n706), .A2(n705), .ZN(n708) );
  AND2_X1 U778 ( .A1(n711), .A2(n739), .ZN(n707) );
  AND2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n714) );
  NOR2_X1 U780 ( .A1(G1981), .A2(G305), .ZN(n709) );
  XOR2_X1 U781 ( .A(n709), .B(KEYINPUT24), .Z(n710) );
  NOR2_X1 U782 ( .A1(n711), .A2(n710), .ZN(n712) );
  AND2_X1 U783 ( .A1(n739), .A2(n712), .ZN(n713) );
  NOR2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n745) );
  NAND2_X1 U785 ( .A1(G107), .A2(n992), .ZN(n716) );
  NAND2_X1 U786 ( .A1(G95), .A2(n996), .ZN(n715) );
  NAND2_X1 U787 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U788 ( .A1(G131), .A2(n995), .ZN(n718) );
  NAND2_X1 U789 ( .A1(G119), .A2(n991), .ZN(n717) );
  NAND2_X1 U790 ( .A1(n718), .A2(n717), .ZN(n719) );
  OR2_X1 U791 ( .A1(n720), .A2(n719), .ZN(n1010) );
  NAND2_X1 U792 ( .A1(G1991), .A2(n1010), .ZN(n731) );
  XOR2_X1 U793 ( .A(KEYINPUT38), .B(KEYINPUT89), .Z(n722) );
  NAND2_X1 U794 ( .A1(G105), .A2(n996), .ZN(n721) );
  XNOR2_X1 U795 ( .A(n722), .B(n721), .ZN(n729) );
  NAND2_X1 U796 ( .A1(G141), .A2(n995), .ZN(n724) );
  NAND2_X1 U797 ( .A1(G129), .A2(n991), .ZN(n723) );
  NAND2_X1 U798 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n992), .A2(G117), .ZN(n725) );
  XOR2_X1 U800 ( .A(KEYINPUT88), .B(n725), .Z(n726) );
  NOR2_X1 U801 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U802 ( .A1(n729), .A2(n728), .ZN(n1004) );
  NAND2_X1 U803 ( .A1(G1996), .A2(n1004), .ZN(n730) );
  NAND2_X1 U804 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U805 ( .A(KEYINPUT90), .B(n732), .Z(n750) );
  INV_X1 U806 ( .A(n750), .ZN(n920) );
  NOR2_X1 U807 ( .A1(G1986), .A2(G290), .ZN(n733) );
  NOR2_X1 U808 ( .A1(G1991), .A2(n1010), .ZN(n922) );
  NOR2_X1 U809 ( .A1(n733), .A2(n922), .ZN(n734) );
  NOR2_X1 U810 ( .A1(n920), .A2(n734), .ZN(n736) );
  NOR2_X1 U811 ( .A1(G1996), .A2(n1004), .ZN(n735) );
  XOR2_X1 U812 ( .A(KEYINPUT101), .B(n735), .Z(n942) );
  NOR2_X1 U813 ( .A1(n736), .A2(n942), .ZN(n737) );
  XNOR2_X1 U814 ( .A(n737), .B(KEYINPUT39), .ZN(n738) );
  XNOR2_X1 U815 ( .A(n738), .B(KEYINPUT102), .ZN(n740) );
  NAND2_X1 U816 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U817 ( .A(KEYINPUT103), .B(n741), .Z(n743) );
  NAND2_X1 U818 ( .A1(n1016), .A2(n742), .ZN(n925) );
  NAND2_X1 U819 ( .A1(n743), .A2(n925), .ZN(n744) );
  NAND2_X1 U820 ( .A1(n744), .A2(n751), .ZN(n748) );
  AND2_X1 U821 ( .A1(n745), .A2(n748), .ZN(n746) );
  NAND2_X1 U822 ( .A1(n747), .A2(n746), .ZN(n756) );
  INV_X1 U823 ( .A(n748), .ZN(n754) );
  XOR2_X1 U824 ( .A(G1986), .B(KEYINPUT86), .Z(n749) );
  XNOR2_X1 U825 ( .A(G290), .B(n749), .ZN(n869) );
  NAND2_X1 U826 ( .A1(n750), .A2(n869), .ZN(n752) );
  NAND2_X1 U827 ( .A1(n752), .A2(n751), .ZN(n753) );
  OR2_X1 U828 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n758) );
  XNOR2_X1 U830 ( .A(n758), .B(n757), .ZN(G329) );
  XOR2_X1 U831 ( .A(G2454), .B(G2446), .Z(n760) );
  XNOR2_X1 U832 ( .A(G2443), .B(KEYINPUT104), .ZN(n759) );
  XNOR2_X1 U833 ( .A(n760), .B(n759), .ZN(n770) );
  XOR2_X1 U834 ( .A(G2451), .B(G2427), .Z(n762) );
  XNOR2_X1 U835 ( .A(G1341), .B(G2435), .ZN(n761) );
  XNOR2_X1 U836 ( .A(n762), .B(n761), .ZN(n766) );
  XOR2_X1 U837 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n764) );
  XNOR2_X1 U838 ( .A(G2430), .B(G2438), .ZN(n763) );
  XNOR2_X1 U839 ( .A(n764), .B(n763), .ZN(n765) );
  XOR2_X1 U840 ( .A(n766), .B(n765), .Z(n768) );
  XNOR2_X1 U841 ( .A(G1348), .B(KEYINPUT105), .ZN(n767) );
  XNOR2_X1 U842 ( .A(n768), .B(n767), .ZN(n769) );
  XNOR2_X1 U843 ( .A(n770), .B(n769), .ZN(n771) );
  AND2_X1 U844 ( .A1(n771), .A2(G14), .ZN(G401) );
  XNOR2_X1 U845 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U847 ( .A(G860), .ZN(n779) );
  OR2_X1 U848 ( .A1(n779), .A2(n968), .ZN(G153) );
  INV_X1 U849 ( .A(G57), .ZN(G237) );
  NAND2_X1 U850 ( .A1(G7), .A2(G661), .ZN(n772) );
  XNOR2_X1 U851 ( .A(n772), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U852 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n774) );
  INV_X1 U853 ( .A(G223), .ZN(n835) );
  NAND2_X1 U854 ( .A1(G567), .A2(n835), .ZN(n773) );
  XNOR2_X1 U855 ( .A(n774), .B(n773), .ZN(G234) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n776) );
  INV_X1 U857 ( .A(G868), .ZN(n817) );
  NAND2_X1 U858 ( .A1(n965), .A2(n817), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n776), .A2(n775), .ZN(G284) );
  INV_X1 U860 ( .A(n851), .ZN(G299) );
  NAND2_X1 U861 ( .A1(G868), .A2(G286), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G299), .A2(n817), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n779), .A2(G559), .ZN(n780) );
  INV_X1 U865 ( .A(n965), .ZN(n797) );
  NAND2_X1 U866 ( .A1(n780), .A2(n797), .ZN(n781) );
  XNOR2_X1 U867 ( .A(n781), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U868 ( .A1(n968), .A2(G868), .ZN(n782) );
  XOR2_X1 U869 ( .A(KEYINPUT73), .B(n782), .Z(n785) );
  NAND2_X1 U870 ( .A1(G868), .A2(n797), .ZN(n783) );
  NOR2_X1 U871 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U873 ( .A(KEYINPUT74), .B(n786), .ZN(G282) );
  XOR2_X1 U874 ( .A(G2100), .B(KEYINPUT76), .Z(n796) );
  NAND2_X1 U875 ( .A1(G111), .A2(n992), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G99), .A2(n996), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U878 ( .A(n789), .B(KEYINPUT75), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G135), .A2(n995), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U881 ( .A1(n991), .A2(G123), .ZN(n792) );
  XOR2_X1 U882 ( .A(KEYINPUT18), .B(n792), .Z(n793) );
  NOR2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n1009) );
  XNOR2_X1 U884 ( .A(G2096), .B(n1009), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(G156) );
  NAND2_X1 U886 ( .A1(G559), .A2(n797), .ZN(n798) );
  XNOR2_X1 U887 ( .A(n798), .B(n968), .ZN(n959) );
  XNOR2_X1 U888 ( .A(KEYINPUT19), .B(G305), .ZN(n799) );
  XNOR2_X1 U889 ( .A(n799), .B(G288), .ZN(n812) );
  NAND2_X1 U890 ( .A1(G93), .A2(n800), .ZN(n803) );
  NAND2_X1 U891 ( .A1(G80), .A2(n801), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n810) );
  NAND2_X1 U893 ( .A1(G55), .A2(n804), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G67), .A2(n805), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U896 ( .A(KEYINPUT77), .B(n808), .Z(n809) );
  NOR2_X1 U897 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U898 ( .A(KEYINPUT78), .B(n811), .Z(n961) );
  XOR2_X1 U899 ( .A(n812), .B(n961), .Z(n814) );
  XNOR2_X1 U900 ( .A(n851), .B(G166), .ZN(n813) );
  XNOR2_X1 U901 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U902 ( .A(n815), .B(G290), .ZN(n967) );
  XNOR2_X1 U903 ( .A(n959), .B(n967), .ZN(n816) );
  NAND2_X1 U904 ( .A1(n816), .A2(G868), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n961), .A2(n817), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n820) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U909 ( .A1(G2090), .A2(n821), .ZN(n822) );
  XNOR2_X1 U910 ( .A(KEYINPUT21), .B(n822), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n823), .A2(G2072), .ZN(G158) );
  NAND2_X1 U912 ( .A1(G69), .A2(G120), .ZN(n824) );
  NOR2_X1 U913 ( .A1(G237), .A2(n824), .ZN(n825) );
  NAND2_X1 U914 ( .A1(G108), .A2(n825), .ZN(n962) );
  NAND2_X1 U915 ( .A1(G567), .A2(n962), .ZN(n826) );
  XNOR2_X1 U916 ( .A(n826), .B(KEYINPUT81), .ZN(n832) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(KEYINPUT80), .Z(n828) );
  NAND2_X1 U918 ( .A1(G132), .A2(G82), .ZN(n827) );
  XNOR2_X1 U919 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n829), .A2(G96), .ZN(n830) );
  OR2_X1 U921 ( .A1(G218), .A2(n830), .ZN(n963) );
  AND2_X1 U922 ( .A1(G2106), .A2(n963), .ZN(n831) );
  NOR2_X1 U923 ( .A1(n832), .A2(n831), .ZN(G319) );
  NAND2_X1 U924 ( .A1(G483), .A2(G661), .ZN(n833) );
  INV_X1 U925 ( .A(G319), .ZN(n1023) );
  NOR2_X1 U926 ( .A1(n833), .A2(n1023), .ZN(n834) );
  XNOR2_X1 U927 ( .A(n834), .B(KEYINPUT82), .ZN(n839) );
  NAND2_X1 U928 ( .A1(G36), .A2(n839), .ZN(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n835), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n836) );
  XOR2_X1 U931 ( .A(KEYINPUT108), .B(n836), .Z(n837) );
  NAND2_X1 U932 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G188) );
  NAND2_X1 U936 ( .A1(G124), .A2(n991), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n840), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U938 ( .A1(G112), .A2(n992), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT113), .B(n841), .Z(n842) );
  NAND2_X1 U940 ( .A1(n843), .A2(n842), .ZN(n848) );
  NAND2_X1 U941 ( .A1(n995), .A2(G136), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n844), .B(KEYINPUT112), .ZN(n846) );
  NAND2_X1 U943 ( .A1(G100), .A2(n996), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n847) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(G162) );
  XNOR2_X1 U946 ( .A(KEYINPUT56), .B(G16), .ZN(n872) );
  XOR2_X1 U947 ( .A(n968), .B(G1341), .Z(n850) );
  XNOR2_X1 U948 ( .A(G171), .B(G1961), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n850), .A2(n849), .ZN(n855) );
  XOR2_X1 U950 ( .A(n965), .B(G1348), .Z(n853) );
  XNOR2_X1 U951 ( .A(n851), .B(G1956), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(n862) );
  NAND2_X1 U954 ( .A1(G1971), .A2(G303), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U957 ( .A(KEYINPUT123), .B(n860), .Z(n861) );
  NAND2_X1 U958 ( .A1(n862), .A2(n861), .ZN(n868) );
  XNOR2_X1 U959 ( .A(G1966), .B(G168), .ZN(n864) );
  NAND2_X1 U960 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U961 ( .A(KEYINPUT57), .B(n865), .Z(n866) );
  XNOR2_X1 U962 ( .A(KEYINPUT122), .B(n866), .ZN(n867) );
  NOR2_X1 U963 ( .A1(n868), .A2(n867), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n870), .A2(n869), .ZN(n871) );
  NAND2_X1 U965 ( .A1(n872), .A2(n871), .ZN(n957) );
  XNOR2_X1 U966 ( .A(G1996), .B(G32), .ZN(n874) );
  XNOR2_X1 U967 ( .A(G1991), .B(G25), .ZN(n873) );
  NOR2_X1 U968 ( .A1(n874), .A2(n873), .ZN(n880) );
  XOR2_X1 U969 ( .A(G2072), .B(G33), .Z(n875) );
  NAND2_X1 U970 ( .A1(n875), .A2(G28), .ZN(n878) );
  XOR2_X1 U971 ( .A(KEYINPUT121), .B(G2067), .Z(n876) );
  XNOR2_X1 U972 ( .A(G26), .B(n876), .ZN(n877) );
  NOR2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U974 ( .A1(n880), .A2(n879), .ZN(n883) );
  XNOR2_X1 U975 ( .A(G27), .B(n881), .ZN(n882) );
  NOR2_X1 U976 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U977 ( .A(KEYINPUT53), .B(n884), .Z(n887) );
  XOR2_X1 U978 ( .A(G34), .B(KEYINPUT54), .Z(n885) );
  XNOR2_X1 U979 ( .A(G2084), .B(n885), .ZN(n886) );
  NAND2_X1 U980 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U981 ( .A(G35), .B(G2090), .ZN(n888) );
  NOR2_X1 U982 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U983 ( .A(KEYINPUT55), .B(n890), .ZN(n892) );
  INV_X1 U984 ( .A(G29), .ZN(n891) );
  NAND2_X1 U985 ( .A1(n892), .A2(n891), .ZN(n893) );
  NAND2_X1 U986 ( .A1(n893), .A2(G11), .ZN(n955) );
  XNOR2_X1 U987 ( .A(G1341), .B(G19), .ZN(n895) );
  XNOR2_X1 U988 ( .A(G1981), .B(G6), .ZN(n894) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U990 ( .A(KEYINPUT124), .B(n896), .ZN(n899) );
  XNOR2_X1 U991 ( .A(n897), .B(G20), .ZN(n898) );
  NAND2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n903) );
  XNOR2_X1 U993 ( .A(KEYINPUT59), .B(G4), .ZN(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(KEYINPUT125), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n901), .B(G1348), .ZN(n902) );
  NOR2_X1 U996 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U997 ( .A(KEYINPUT60), .B(n904), .ZN(n909) );
  XNOR2_X1 U998 ( .A(G1966), .B(G21), .ZN(n907) );
  XNOR2_X1 U999 ( .A(n905), .B(G5), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(n907), .A2(n906), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(n909), .A2(n908), .ZN(n916) );
  XNOR2_X1 U1002 ( .A(G1971), .B(G22), .ZN(n911) );
  XNOR2_X1 U1003 ( .A(G23), .B(G1976), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(n911), .A2(n910), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G1986), .B(G24), .Z(n912) );
  NAND2_X1 U1006 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(KEYINPUT58), .B(n914), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1009 ( .A(KEYINPUT61), .B(n917), .Z(n918) );
  NOR2_X1 U1010 ( .A1(G16), .A2(n918), .ZN(n919) );
  XOR2_X1 U1011 ( .A(KEYINPUT126), .B(n919), .Z(n953) );
  NOR2_X1 U1012 ( .A1(n921), .A2(n920), .ZN(n930) );
  NOR2_X1 U1013 ( .A1(n922), .A2(n1009), .ZN(n923) );
  XOR2_X1 U1014 ( .A(KEYINPUT119), .B(n923), .Z(n924) );
  NAND2_X1 U1015 ( .A1(n925), .A2(n924), .ZN(n928) );
  XOR2_X1 U1016 ( .A(G2084), .B(G160), .Z(n926) );
  XNOR2_X1 U1017 ( .A(KEYINPUT118), .B(n926), .ZN(n927) );
  NOR2_X1 U1018 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1019 ( .A1(n930), .A2(n929), .ZN(n947) );
  NAND2_X1 U1020 ( .A1(G139), .A2(n995), .ZN(n932) );
  NAND2_X1 U1021 ( .A1(G103), .A2(n996), .ZN(n931) );
  NAND2_X1 U1022 ( .A1(n932), .A2(n931), .ZN(n937) );
  NAND2_X1 U1023 ( .A1(G127), .A2(n991), .ZN(n934) );
  NAND2_X1 U1024 ( .A1(G115), .A2(n992), .ZN(n933) );
  NAND2_X1 U1025 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1026 ( .A(KEYINPUT47), .B(n935), .Z(n936) );
  NOR2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n1015) );
  XOR2_X1 U1028 ( .A(G2072), .B(n1015), .Z(n939) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n940), .ZN(n945) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n941) );
  NOR2_X1 U1033 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n943), .Z(n944) );
  NAND2_X1 U1035 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1036 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1037 ( .A(KEYINPUT52), .B(n948), .Z(n949) );
  NOR2_X1 U1038 ( .A1(KEYINPUT55), .A2(n949), .ZN(n950) );
  XOR2_X1 U1039 ( .A(KEYINPUT120), .B(n950), .Z(n951) );
  NAND2_X1 U1040 ( .A1(G29), .A2(n951), .ZN(n952) );
  NAND2_X1 U1041 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1042 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1043 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1044 ( .A(KEYINPUT62), .B(n958), .Z(G311) );
  XNOR2_X1 U1045 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  NOR2_X1 U1046 ( .A1(n959), .A2(G860), .ZN(n960) );
  XOR2_X1 U1047 ( .A(n961), .B(n960), .Z(G145) );
  INV_X1 U1048 ( .A(G132), .ZN(G219) );
  INV_X1 U1049 ( .A(G120), .ZN(G236) );
  INV_X1 U1050 ( .A(G96), .ZN(G221) );
  INV_X1 U1051 ( .A(G82), .ZN(G220) );
  INV_X1 U1052 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1053 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(KEYINPUT109), .B(n964), .ZN(G261) );
  INV_X1 U1055 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U1056 ( .A(G171), .B(n965), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n966), .B(G286), .ZN(n970) );
  XNOR2_X1 U1058 ( .A(n968), .B(n967), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(n970), .B(n969), .ZN(n971) );
  NOR2_X1 U1060 ( .A1(G37), .A2(n971), .ZN(G397) );
  XOR2_X1 U1061 ( .A(KEYINPUT111), .B(G2678), .Z(n973) );
  XNOR2_X1 U1062 ( .A(G2072), .B(G2090), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1064 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n975) );
  XNOR2_X1 U1065 ( .A(G2067), .B(KEYINPUT42), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n975), .B(n974), .ZN(n976) );
  XOR2_X1 U1067 ( .A(n977), .B(n976), .Z(n979) );
  XNOR2_X1 U1068 ( .A(G2100), .B(G2096), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(n979), .B(n978), .ZN(n981) );
  XOR2_X1 U1070 ( .A(G2078), .B(G2084), .Z(n980) );
  XNOR2_X1 U1071 ( .A(n981), .B(n980), .ZN(G227) );
  XOR2_X1 U1072 ( .A(G1981), .B(G1971), .Z(n983) );
  XNOR2_X1 U1073 ( .A(G1996), .B(G1966), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n983), .B(n982), .ZN(n984) );
  XOR2_X1 U1075 ( .A(n984), .B(KEYINPUT41), .Z(n986) );
  XNOR2_X1 U1076 ( .A(G1991), .B(G1976), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(n986), .B(n985), .ZN(n990) );
  XOR2_X1 U1078 ( .A(G2474), .B(G1956), .Z(n988) );
  XNOR2_X1 U1079 ( .A(G1986), .B(G1961), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n988), .B(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n990), .B(n989), .ZN(G229) );
  NAND2_X1 U1082 ( .A1(G130), .A2(n991), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(G118), .A2(n992), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n1001) );
  NAND2_X1 U1085 ( .A1(G142), .A2(n995), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(G106), .A2(n996), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT45), .B(n999), .Z(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1014) );
  XOR2_X1 U1090 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1003), .B(n1002), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(n1004), .B(G162), .ZN(n1006) );
  XNOR2_X1 U1094 ( .A(G164), .B(G160), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1008), .B(n1007), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(n1010), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(n1012), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1014), .B(n1013), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(n1016), .B(n1015), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NOR2_X1 U1102 ( .A1(G37), .A2(n1019), .ZN(G395) );
  NOR2_X1 U1103 ( .A1(G227), .A2(G229), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(KEYINPUT117), .B(n1020), .Z(n1021) );
  XNOR2_X1 U1105 ( .A(n1021), .B(KEYINPUT49), .ZN(n1022) );
  NOR2_X1 U1106 ( .A1(G397), .A2(n1022), .ZN(n1027) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(G401), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT116), .B(n1024), .Z(n1025) );
  NOR2_X1 U1109 ( .A1(G395), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(G225) );
  INV_X1 U1111 ( .A(G225), .ZN(G308) );
  INV_X1 U1112 ( .A(G108), .ZN(G238) );
endmodule

