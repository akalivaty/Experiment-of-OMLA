//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n533, new_n535, new_n536, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n579, new_n580, new_n583,
    new_n585, new_n586, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G221), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT67), .Z(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT68), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n464), .A2(new_n472), .ZN(G160));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n461), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n467), .A2(G136), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  NAND2_X1  g056(.A1(new_n470), .A2(G102), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n465), .A2(new_n466), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n483), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n484), .B2(new_n474), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n474), .C1(new_n459), .C2(new_n460), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n483), .A2(KEYINPUT4), .A3(G138), .A4(new_n474), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n485), .A2(new_n490), .ZN(G164));
  INV_X1    g066(.A(G543), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(KEYINPUT69), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT5), .A3(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(KEYINPUT6), .B(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G88), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  XNOR2_X1  g079(.A(new_n503), .B(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(G303));
  INV_X1    g084(.A(G303), .ZN(G166));
  XNOR2_X1  g085(.A(new_n501), .B(KEYINPUT71), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G51), .ZN(new_n512));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT72), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT7), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n498), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n516));
  INV_X1    g091(.A(new_n497), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n512), .A2(new_n515), .A3(new_n518), .ZN(G168));
  NAND2_X1  g094(.A1(new_n511), .A2(G52), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n497), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n521), .A2(new_n507), .ZN(new_n522));
  INV_X1    g097(.A(new_n499), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G90), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(G301));
  INV_X1    g100(.A(G301), .ZN(G171));
  NAND2_X1  g101(.A1(new_n511), .A2(G43), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n497), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n507), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n523), .A2(G81), .ZN(new_n530));
  AND3_X1   g105(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G860), .ZN(G153));
  AND3_X1   g107(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G36), .ZN(G176));
  NAND2_X1  g109(.A1(G1), .A2(G3), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT8), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n533), .A2(new_n536), .ZN(G188));
  AOI22_X1  g112(.A1(new_n497), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G91), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n538), .A2(new_n507), .B1(new_n539), .B2(new_n499), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT6), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G651), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n542), .A2(new_n544), .A3(G53), .A4(G543), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT9), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(G299));
  INV_X1    g125(.A(G168), .ZN(G286));
  OAI21_X1  g126(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n552));
  AND3_X1   g127(.A1(new_n542), .A2(new_n544), .A3(G543), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n552), .A2(KEYINPUT74), .B1(G49), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n523), .A2(G87), .ZN(new_n555));
  OAI211_X1 g130(.A(new_n554), .B(new_n555), .C1(KEYINPUT74), .C2(new_n552), .ZN(G288));
  NAND2_X1  g131(.A1(new_n553), .A2(G48), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n497), .A2(G86), .A3(new_n498), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n497), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n557), .B(new_n558), .C1(new_n559), .C2(new_n507), .ZN(G305));
  XOR2_X1   g135(.A(KEYINPUT75), .B(G85), .Z(new_n561));
  NAND2_X1  g136(.A1(new_n523), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n553), .B(KEYINPUT71), .ZN(new_n564));
  INV_X1    g139(.A(G47), .ZN(new_n565));
  OAI221_X1 g140(.A(new_n562), .B1(new_n507), .B2(new_n563), .C1(new_n564), .C2(new_n565), .ZN(G290));
  NAND2_X1  g141(.A1(G301), .A2(G868), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n523), .A2(G92), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n497), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT76), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n511), .A2(G54), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n567), .B1(new_n576), .B2(G868), .ZN(G284));
  OAI21_X1  g152(.A(new_n567), .B1(new_n576), .B2(G868), .ZN(G321));
  INV_X1    g153(.A(G868), .ZN(new_n579));
  NAND2_X1  g154(.A1(G299), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n580), .B1(new_n579), .B2(G168), .ZN(G297));
  OAI21_X1  g156(.A(new_n580), .B1(new_n579), .B2(G168), .ZN(G280));
  INV_X1    g157(.A(G559), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n576), .B1(new_n583), .B2(G860), .ZN(G148));
  NAND2_X1  g159(.A1(new_n576), .A2(new_n583), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G868), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(G868), .B2(new_n531), .ZN(G323));
  XNOR2_X1  g162(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g163(.A1(new_n483), .A2(new_n470), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT12), .Z(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT13), .Z(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(G2100), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n474), .A2(G111), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n469), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI221_X1 g170(.A(new_n595), .B1(new_n594), .B2(new_n593), .C1(G99), .C2(G2105), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n475), .A2(G123), .B1(G135), .B2(new_n467), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g173(.A(KEYINPUT78), .B(G2096), .Z(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n600), .ZN(G156));
  XNOR2_X1  g176(.A(KEYINPUT15), .B(G2435), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(G2438), .ZN(new_n603));
  XOR2_X1   g178(.A(G2427), .B(G2430), .Z(new_n604));
  XNOR2_X1  g179(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT79), .B(KEYINPUT14), .Z(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(G2443), .B(G2446), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n610));
  XNOR2_X1  g185(.A(G1341), .B(G1348), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n609), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(G2451), .B(G2454), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G14), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT81), .ZN(G401));
  XOR2_X1   g192(.A(G2084), .B(G2090), .Z(new_n618));
  XNOR2_X1  g193(.A(G2067), .B(G2678), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n620), .A2(KEYINPUT17), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n618), .A2(new_n619), .ZN(new_n622));
  AOI21_X1  g197(.A(KEYINPUT18), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2072), .B(G2078), .Z(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n620), .B2(KEYINPUT18), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G2096), .B(G2100), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(G227));
  XNOR2_X1  g203(.A(G1971), .B(G1976), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT19), .ZN(new_n630));
  XOR2_X1   g205(.A(G1956), .B(G2474), .Z(new_n631));
  XOR2_X1   g206(.A(G1961), .B(G1966), .Z(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n630), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n631), .A2(new_n632), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n634), .A2(KEYINPUT20), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n638), .A2(new_n630), .A3(new_n633), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n637), .B(new_n639), .C1(KEYINPUT20), .C2(new_n634), .ZN(new_n640));
  XOR2_X1   g215(.A(G1991), .B(G1996), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n640), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1981), .B(G1986), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(G229));
  NOR2_X1   g222(.A1(G29), .A2(G33), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n470), .A2(G103), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT25), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n467), .A2(G139), .ZN(new_n651));
  AOI22_X1  g226(.A1(new_n483), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n650), .B(new_n651), .C1(new_n474), .C2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n648), .B1(new_n654), .B2(G29), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(G2072), .Z(new_n656));
  INV_X1    g231(.A(G16), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G4), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n576), .B2(new_n657), .ZN(new_n659));
  INV_X1    g234(.A(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  AOI22_X1  g236(.A1(new_n475), .A2(G129), .B1(G141), .B2(new_n467), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n470), .A2(G105), .ZN(new_n663));
  NAND3_X1  g238(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT26), .Z(new_n665));
  NAND3_X1  g240(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  MUX2_X1   g241(.A(G32), .B(new_n666), .S(G29), .Z(new_n667));
  XOR2_X1   g242(.A(KEYINPUT27), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(G27), .ZN(new_n670));
  OAI21_X1  g245(.A(KEYINPUT92), .B1(new_n670), .B2(G29), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n670), .A2(KEYINPUT92), .A3(G29), .ZN(new_n672));
  INV_X1    g247(.A(G29), .ZN(new_n673));
  OAI211_X1 g248(.A(new_n671), .B(new_n672), .C1(G164), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G2078), .ZN(new_n675));
  INV_X1    g250(.A(G28), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(KEYINPUT30), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(KEYINPUT30), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n678), .A3(new_n673), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n598), .B2(new_n673), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n669), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n656), .A2(new_n661), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n657), .A2(G20), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT94), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT23), .ZN(new_n685));
  INV_X1    g260(.A(G299), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n657), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT95), .Z(new_n688));
  AOI21_X1  g263(.A(new_n682), .B1(G1956), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G11), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n673), .A2(G35), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G162), .B2(new_n673), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2090), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G16), .A2(G19), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n531), .B2(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G1341), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(G168), .A2(G16), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G16), .B2(G21), .ZN(new_n701));
  INV_X1    g276(.A(G1966), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT88), .B(G34), .Z(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT24), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT24), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n673), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G160), .B2(new_n673), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  INV_X1    g284(.A(G2084), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT90), .B1(G5), .B2(G16), .ZN(new_n712));
  OR3_X1    g287(.A1(KEYINPUT90), .A2(G5), .A3(G16), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n712), .B(new_n713), .C1(G301), .C2(new_n657), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT91), .B(G1961), .Z(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n703), .A2(new_n711), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n701), .A2(new_n702), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n719), .B1(G1341), .B2(new_n697), .C1(new_n710), .C2(new_n709), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT28), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n673), .A2(G26), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n475), .A2(G128), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n467), .A2(G140), .ZN(new_n724));
  NOR2_X1   g299(.A1(G104), .A2(G2105), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(new_n474), .B2(G116), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n721), .B(new_n722), .C1(new_n727), .C2(G29), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n721), .B2(new_n722), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT86), .B(G2067), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NOR4_X1   g306(.A1(new_n699), .A2(new_n718), .A3(new_n720), .A4(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n688), .A2(G1956), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n689), .A2(new_n690), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT96), .Z(new_n735));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n736));
  MUX2_X1   g311(.A(G24), .B(G290), .S(G16), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1986), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n657), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n657), .ZN(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n657), .A2(G6), .ZN(new_n743));
  INV_X1    g318(.A(G305), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n657), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT83), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT32), .B(G1981), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(KEYINPUT84), .B1(G16), .B2(G23), .ZN(new_n749));
  OR3_X1    g324(.A1(KEYINPUT84), .A2(G16), .A3(G23), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n749), .B(new_n750), .C1(G288), .C2(new_n657), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT33), .B(G1976), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n742), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n736), .B(new_n738), .C1(new_n754), .C2(KEYINPUT34), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n673), .A2(G25), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n475), .A2(G119), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n467), .A2(G131), .ZN(new_n758));
  OR2_X1    g333(.A1(G95), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n673), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT35), .B(G1991), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n763), .B(new_n765), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n755), .B(new_n766), .C1(KEYINPUT34), .C2(new_n754), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT36), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n735), .A2(new_n768), .ZN(G150));
  INV_X1    g344(.A(G150), .ZN(G311));
  NAND2_X1  g345(.A1(new_n523), .A2(G93), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n497), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n772));
  INV_X1    g347(.A(G55), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n771), .B1(new_n507), .B2(new_n772), .C1(new_n564), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G860), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT37), .Z(new_n776));
  NOR2_X1   g351(.A1(new_n575), .A2(new_n583), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT39), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n531), .B(new_n774), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(G860), .ZN(G145));
  NAND2_X1  g358(.A1(new_n475), .A2(G130), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT99), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(G106), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G118), .C2(new_n474), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n467), .A2(G142), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(new_n761), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n793), .A2(new_n590), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n590), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(G114), .A2(G2104), .ZN(new_n798));
  INV_X1    g373(.A(G126), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n461), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n800), .A2(G2105), .B1(G102), .B2(new_n470), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT98), .ZN(new_n802));
  AOI21_X1  g377(.A(KEYINPUT98), .B1(new_n488), .B2(new_n489), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(new_n727), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(new_n666), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(new_n653), .ZN(new_n807));
  INV_X1    g382(.A(new_n654), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n797), .A2(new_n810), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n795), .A2(new_n796), .B1(new_n807), .B2(new_n809), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n598), .B(G160), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(new_n480), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n811), .A2(new_n812), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT103), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(KEYINPUT103), .ZN(new_n820));
  AOI21_X1  g395(.A(G37), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT101), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n811), .A2(new_n822), .A3(new_n812), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n823), .B(new_n814), .C1(new_n822), .C2(new_n812), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g401(.A(G303), .B(G290), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(G288), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(G288), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(new_n744), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n744), .B1(new_n828), .B2(new_n829), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT42), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT105), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n827), .B(G288), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G305), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n830), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT105), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT42), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n841));
  NAND3_X1  g416(.A1(new_n836), .A2(new_n830), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT107), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g419(.A1(new_n836), .A2(KEYINPUT107), .A3(new_n830), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n575), .B(G299), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT41), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n781), .B(new_n585), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(new_n847), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n848), .B2(new_n849), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n854), .B2(new_n851), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n840), .A2(new_n846), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n840), .B2(new_n846), .ZN(new_n857));
  OAI21_X1  g432(.A(G868), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n774), .A2(new_n579), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(G295));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n858), .A2(new_n861), .A3(new_n859), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n861), .B1(new_n858), .B2(new_n859), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(G331));
  NOR2_X1   g439(.A1(new_n781), .A2(G171), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n774), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(G301), .ZN(new_n868));
  OAI21_X1  g443(.A(G286), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n781), .A2(G171), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(G301), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(G168), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n847), .A3(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n869), .A2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n874), .B2(new_n848), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(new_n837), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT109), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n878), .A3(new_n837), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n875), .B2(new_n837), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n876), .B(new_n877), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT43), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n875), .A2(new_n837), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(KEYINPUT109), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n885), .B2(new_n879), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n887), .A3(new_n876), .ZN(new_n888));
  XNOR2_X1  g463(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n883), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT44), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n883), .B2(new_n888), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(G397));
  INV_X1    g469(.A(G8), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT111), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT4), .B1(new_n467), .B2(G138), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n486), .A2(new_n487), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT98), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n485), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n896), .B1(new_n902), .B2(G1384), .ZN(new_n903));
  INV_X1    g478(.A(G1384), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n804), .A2(KEYINPUT111), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(G160), .A2(G40), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n895), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT49), .ZN(new_n910));
  XNOR2_X1  g485(.A(G305), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT113), .B1(new_n559), .B2(new_n507), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(G1981), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(G1981), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n744), .A2(new_n910), .ZN(new_n915));
  NOR2_X1   g490(.A1(G305), .A2(KEYINPUT49), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT114), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n918), .A2(new_n909), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n918), .B2(new_n909), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n922), .A2(G1976), .A3(G288), .ZN(new_n923));
  NOR2_X1   g498(.A1(G305), .A2(G1981), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n909), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n804), .A2(KEYINPUT45), .A3(new_n904), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n904), .B1(new_n485), .B2(new_n490), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n908), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n741), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n902), .A2(new_n896), .A3(G1384), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT111), .B1(new_n804), .B2(new_n904), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT112), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n907), .B1(new_n927), .B2(KEYINPUT50), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n906), .A2(new_n938), .A3(new_n932), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n931), .B1(new_n940), .B2(G2090), .ZN(new_n941));
  NAND2_X1  g516(.A1(G303), .A2(G8), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(G8), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n908), .B1(new_n933), .B2(new_n934), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G8), .ZN(new_n947));
  INV_X1    g522(.A(G1976), .ZN(new_n948));
  NOR2_X1   g523(.A1(G288), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT52), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT52), .B1(G288), .B2(new_n948), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n909), .B(new_n951), .C1(new_n948), .C2(G288), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n950), .B(new_n952), .C1(new_n920), .C2(new_n921), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n925), .B1(new_n945), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(KEYINPUT115), .B(G2084), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n936), .A2(new_n937), .A3(new_n939), .A4(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n927), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT45), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n908), .B(new_n958), .C1(new_n906), .C2(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n702), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(G8), .A3(G168), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT116), .ZN(new_n963));
  INV_X1    g538(.A(new_n953), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n903), .A2(KEYINPUT50), .A3(new_n905), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n957), .A2(new_n932), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n966), .A3(new_n908), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n931), .B1(new_n967), .B2(G2090), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G8), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n943), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n964), .A2(new_n970), .A3(new_n945), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n963), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT63), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n941), .A2(new_n976), .A3(G8), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n941), .B2(G8), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n943), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n964), .A2(new_n945), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n963), .A2(new_n979), .A3(KEYINPUT63), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n954), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(G168), .A2(new_n895), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n956), .B2(new_n960), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n961), .A2(G8), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n984), .ZN(new_n988));
  OAI211_X1 g563(.A(KEYINPUT51), .B(G8), .C1(new_n961), .C2(G286), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT62), .B(new_n985), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  OR3_X1    g566(.A1(new_n959), .A2(new_n991), .A3(G2078), .ZN(new_n992));
  INV_X1    g567(.A(G1961), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n940), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n930), .B2(G2078), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G171), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n998), .A2(new_n970), .A3(new_n945), .A4(new_n964), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT127), .B1(new_n990), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n971), .A2(new_n997), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n988), .A2(new_n989), .ZN(new_n1003));
  INV_X1    g578(.A(new_n985), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1001), .B(new_n1002), .C1(new_n1005), .C2(KEYINPUT62), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT121), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n938), .B1(new_n906), .B2(new_n932), .ZN(new_n1010));
  AOI211_X1 g585(.A(KEYINPUT112), .B(KEYINPUT50), .C1(new_n903), .C2(new_n905), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1348), .B1(new_n1012), .B2(new_n937), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT120), .B1(new_n906), .B2(new_n908), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n1015), .B(new_n907), .C1(new_n903), .C2(new_n905), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1014), .A2(new_n1016), .A3(G2067), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1009), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1017), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n940), .A2(new_n660), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1020), .A3(KEYINPUT121), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1956), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n967), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n930), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n547), .B1(new_n540), .B2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g605(.A(KEYINPUT118), .B1(new_n499), .B2(new_n539), .C1(new_n538), .C2(new_n507), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1028), .B(KEYINPUT57), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n540), .A2(new_n1029), .ZN(new_n1033));
  INV_X1    g608(.A(new_n547), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT119), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1032), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n541), .B(KEYINPUT57), .C1(new_n548), .C2(new_n549), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1024), .A2(new_n1027), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n576), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n967), .A2(new_n1023), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1028), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1035), .A2(KEYINPUT119), .A3(new_n1036), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n1044), .A2(new_n1047), .A3(new_n1039), .A4(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1022), .A2(new_n1042), .B1(new_n1043), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT61), .ZN(new_n1052));
  AND3_X1   g627(.A1(new_n1024), .A2(new_n1027), .A3(new_n1040), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1040), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT61), .B(new_n1041), .C1(new_n1050), .C2(new_n1043), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n1057));
  XOR2_X1   g632(.A(KEYINPUT58), .B(G1341), .Z(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n930), .A2(G1996), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1057), .B1(new_n1062), .B2(new_n531), .ZN(new_n1063));
  AOI211_X1 g638(.A(KEYINPUT59), .B(new_n866), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1055), .B(new_n1056), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT123), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1058), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n946), .A2(new_n1015), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n906), .A2(KEYINPUT120), .A3(new_n908), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n531), .B1(new_n1070), .B2(new_n1060), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT59), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1062), .A2(new_n1057), .A3(new_n531), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1056), .A4(new_n1055), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1066), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT60), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1018), .A2(new_n1078), .A3(new_n1021), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n575), .B1(new_n1022), .B2(KEYINPUT60), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n1078), .B(new_n576), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1051), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n804), .A2(new_n904), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n472), .B1(new_n1085), .B2(new_n928), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n463), .B(KEYINPUT124), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G2105), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(G2078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(G2078), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n991), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1088), .A2(G40), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1086), .A2(new_n926), .A3(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n1094), .B(KEYINPUT126), .Z(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n995), .A3(new_n994), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1084), .B1(new_n998), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(G171), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(KEYINPUT54), .C1(G171), .C2(new_n996), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1098), .A2(new_n1005), .A3(new_n1100), .A4(new_n972), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n982), .B(new_n1008), .C1(new_n1083), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1996), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n666), .B(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G2067), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n727), .B(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n765), .B2(new_n762), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n765), .B2(new_n762), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(G1986), .B2(G290), .ZN(new_n1110));
  OR2_X1    g685(.A1(G290), .A2(G1986), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1085), .A2(new_n928), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(new_n907), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1102), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1114), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1117), .A2(new_n1111), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT48), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1114), .B2(new_n1109), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT46), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1117), .B2(G1996), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1106), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1114), .B1(new_n666), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1114), .A2(KEYINPUT46), .A3(new_n1103), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT47), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n762), .A2(new_n765), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1107), .A2(new_n1128), .B1(G2067), .B2(new_n727), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1120), .B(new_n1127), .C1(new_n1114), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1116), .A2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g706(.A(new_n456), .ZN(new_n1133));
  NOR2_X1   g707(.A1(G227), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g708(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g709(.A(new_n1135), .B1(new_n821), .B2(new_n824), .ZN(new_n1136));
  NAND2_X1  g710(.A1(new_n883), .A2(new_n888), .ZN(new_n1137));
  AOI21_X1  g711(.A(G229), .B1(G14), .B2(new_n615), .ZN(new_n1138));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(G225));
  INV_X1    g713(.A(G225), .ZN(G308));
endmodule


