//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1244, new_n1245, new_n1246, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(G244), .Z(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G87), .A2(G250), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  OAI211_X1 g0047(.A(new_n247), .B(new_n217), .C1(G1), .C2(new_n208), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n208), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G150), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n208), .A2(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n252), .A2(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(G20), .B2(new_n204), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n247), .A2(new_n217), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n250), .B1(G50), .B2(new_n251), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT9), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G222), .ZN(new_n264));
  INV_X1    g0064(.A(G223), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n262), .B(new_n264), .C1(new_n265), .C2(new_n263), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n266), .B(new_n269), .C1(G77), .C2(new_n262), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT65), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(new_n217), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n267), .A2(KEYINPUT65), .A3(G1), .A4(G13), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n273), .A2(new_n275), .A3(G274), .A4(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G226), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n273), .A2(new_n276), .A3(new_n274), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n270), .B(new_n277), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G190), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(G200), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n261), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT10), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT10), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n261), .A2(new_n287), .A3(new_n283), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n281), .A2(G179), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n281), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n260), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G238), .A2(G1698), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n262), .B(new_n295), .C1(new_n234), .C2(G1698), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n296), .B(new_n269), .C1(G107), .C2(new_n262), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n277), .C1(new_n220), .C2(new_n280), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n298), .A2(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n291), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT15), .B(G87), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n253), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n302), .A2(new_n303), .B1(G20), .B2(G77), .ZN(new_n304));
  INV_X1    g0104(.A(new_n252), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n259), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n251), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n221), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n221), .B2(new_n248), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n299), .A2(new_n300), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n298), .A2(G200), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n312), .C1(new_n282), .C2(new_n298), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n203), .A2(G20), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n319), .B1(new_n253), .B2(new_n221), .C1(new_n201), .C2(new_n256), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n247), .A2(new_n217), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT11), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT12), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n249), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G13), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n325), .A2(new_n328), .A3(G1), .ZN(new_n329));
  INV_X1    g0129(.A(new_n319), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n329), .A2(new_n330), .B1(new_n325), .B2(new_n251), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n322), .B2(new_n323), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(G226), .A2(G1698), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n234), .B2(G1698), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n262), .B1(G33), .B2(G97), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n337), .A2(new_n268), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n273), .A2(G238), .A3(new_n276), .A4(new_n274), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n277), .A4(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n277), .B(new_n340), .C1(new_n337), .C2(new_n268), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT67), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT14), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(G169), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(G179), .A3(new_n343), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n344), .B2(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n334), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n334), .B1(G200), .B2(new_n344), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n282), .B2(new_n344), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n305), .A2(new_n248), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT69), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n252), .A2(new_n251), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n355), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT68), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G58), .A2(G68), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n208), .B1(new_n214), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n306), .A2(G159), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n361), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(G58), .A2(G68), .ZN(new_n367));
  NOR2_X1   g0167(.A1(G58), .A2(G68), .ZN(new_n368));
  OAI21_X1  g0168(.A(G20), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT68), .A3(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT7), .B1(new_n374), .B2(new_n208), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR4_X1   g0176(.A1(new_n372), .A2(new_n373), .A3(new_n376), .A4(G20), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n259), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n371), .A2(new_n378), .A3(KEYINPUT16), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n360), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n265), .A2(new_n263), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n278), .A2(G1698), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(new_n372), .C2(new_n373), .ZN(new_n386));
  INV_X1    g0186(.A(G87), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n255), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(KEYINPUT70), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT70), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n386), .A2(new_n392), .A3(new_n389), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n391), .A2(new_n269), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G179), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n273), .A2(G232), .A3(new_n276), .A4(new_n274), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n277), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n277), .A2(new_n396), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n268), .B1(new_n390), .B2(KEYINPUT70), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n393), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(G169), .B2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n383), .A2(KEYINPUT18), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT18), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n369), .A2(KEYINPUT68), .A3(new_n364), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT68), .B1(new_n369), .B2(new_n364), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OR2_X1    g0207(.A1(KEYINPUT3), .A2(G33), .ZN(new_n408));
  NAND2_X1  g0208(.A1(KEYINPUT3), .A2(G33), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n208), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n376), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n408), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n409), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n203), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n380), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(new_n321), .A3(new_n382), .ZN(new_n415));
  INV_X1    g0215(.A(new_n360), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n418));
  AOI21_X1  g0218(.A(G169), .B1(new_n394), .B2(new_n397), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n404), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n403), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G223), .A2(G1698), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n278), .B2(G1698), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n388), .B1(new_n424), .B2(new_n262), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n269), .B1(new_n425), .B2(new_n392), .ZN(new_n426));
  INV_X1    g0226(.A(new_n393), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n397), .B(new_n282), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G200), .B2(new_n401), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n429), .A2(new_n416), .A3(new_n415), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT17), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n383), .A2(new_n432), .A3(new_n429), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n422), .A2(new_n434), .ZN(new_n435));
  NOR4_X1   g0235(.A1(new_n294), .A2(new_n318), .A3(new_n354), .A4(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT76), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  INV_X1    g0240(.A(G41), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT5), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G41), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n440), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n445), .A2(G274), .A3(new_n273), .A4(new_n276), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n440), .A2(new_n442), .A3(new_n444), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n447), .A2(new_n273), .A3(G270), .A4(new_n276), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n263), .A2(G257), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G264), .A2(G1698), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n451), .C1(new_n372), .C2(new_n373), .ZN(new_n452));
  INV_X1    g0252(.A(G303), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n408), .A2(new_n453), .A3(new_n409), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n269), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT73), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n452), .A2(new_n454), .A3(new_n269), .A4(KEYINPUT73), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n449), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G169), .ZN(new_n461));
  INV_X1    g0261(.A(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n309), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n207), .A2(G33), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n259), .A2(new_n251), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n465), .B2(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n208), .C1(G33), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n462), .A2(G20), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT74), .B1(new_n321), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(KEYINPUT20), .B(new_n469), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n438), .B1(new_n461), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n477), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n291), .B1(new_n449), .B2(new_n459), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(KEYINPUT76), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT21), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n460), .A2(G200), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n477), .C1(new_n282), .C2(new_n460), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT75), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n457), .A2(new_n458), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n446), .A2(new_n448), .ZN(new_n488));
  OAI211_X1 g0288(.A(KEYINPUT21), .B(G169), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n449), .A2(new_n459), .A3(G179), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n486), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  AOI211_X1 g0292(.A(KEYINPUT75), .B(new_n477), .C1(new_n489), .C2(new_n490), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n483), .B(new_n485), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n302), .A2(new_n251), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n465), .A2(new_n387), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n208), .B(G68), .C1(new_n372), .C2(new_n373), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT72), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT72), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n262), .A2(new_n499), .A3(new_n208), .A4(G68), .ZN(new_n500));
  OR2_X1    g0300(.A1(KEYINPUT71), .A2(KEYINPUT19), .ZN(new_n501));
  NAND2_X1  g0301(.A1(KEYINPUT71), .A2(KEYINPUT19), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(new_n253), .C2(new_n468), .ZN(new_n503));
  XNOR2_X1  g0303(.A(KEYINPUT71), .B(KEYINPUT19), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n387), .A2(new_n468), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n208), .B1(new_n255), .B2(new_n468), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n498), .A2(new_n500), .A3(new_n503), .A4(new_n508), .ZN(new_n509));
  AOI211_X1 g0309(.A(new_n495), .B(new_n496), .C1(new_n509), .C2(new_n321), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n439), .A2(G1), .A3(G274), .ZN(new_n511));
  INV_X1    g0311(.A(G250), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n439), .B2(G1), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n273), .A2(new_n511), .A3(new_n276), .A4(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G238), .A2(G1698), .ZN(new_n515));
  INV_X1    g0315(.A(G244), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(G1698), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(new_n262), .B1(G33), .B2(G116), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n282), .B(new_n514), .C1(new_n518), .C2(new_n268), .ZN(new_n519));
  AND4_X1   g0319(.A1(new_n273), .A2(new_n511), .A3(new_n276), .A4(new_n513), .ZN(new_n520));
  OR2_X1    g0320(.A1(G238), .A2(G1698), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n516), .A2(G1698), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n521), .B(new_n522), .C1(new_n372), .C2(new_n373), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G116), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n268), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n519), .B1(new_n526), .B2(G200), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n509), .A2(new_n321), .ZN(new_n528));
  INV_X1    g0328(.A(new_n495), .ZN(new_n529));
  INV_X1    g0329(.A(new_n465), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n302), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(G179), .B(new_n514), .C1(new_n518), .C2(new_n268), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n526), .B2(new_n291), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n510), .A2(new_n527), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  AND3_X1   g0335(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI22_X1  g0339(.A1(new_n539), .A2(new_n208), .B1(new_n221), .B2(new_n256), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n505), .B1(new_n411), .B2(new_n412), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n321), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n251), .A2(G97), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n465), .B2(new_n468), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT4), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n374), .B2(new_n516), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(G1698), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n262), .A2(G244), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n467), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n262), .A2(G250), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n263), .B1(new_n553), .B2(KEYINPUT4), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n269), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n447), .A2(new_n273), .A3(G257), .A4(new_n276), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n446), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n395), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n446), .A2(new_n556), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n512), .B1(new_n408), .B2(new_n409), .ZN(new_n560));
  OAI21_X1  g0360(.A(G1698), .B1(new_n560), .B2(new_n548), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n561), .A2(new_n467), .A3(new_n549), .A4(new_n551), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n559), .B1(new_n562), .B2(new_n269), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n547), .B(new_n558), .C1(G169), .C2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(G107), .B1(new_n375), .B2(new_n377), .ZN(new_n565));
  AND2_X1   g0365(.A1(G97), .A2(G107), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G97), .A2(G107), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n538), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(G20), .B1(G77), .B2(new_n306), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n545), .B1(new_n572), .B2(new_n321), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n555), .A2(G190), .A3(new_n557), .ZN(new_n574));
  INV_X1    g0374(.A(G200), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(new_n563), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n535), .A2(new_n564), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT25), .ZN(new_n578));
  AOI211_X1 g0378(.A(G107), .B(new_n251), .C1(KEYINPUT78), .C2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(KEYINPUT78), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n530), .A2(G107), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n208), .B2(G107), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n505), .A2(KEYINPUT23), .A3(G20), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n303), .A2(G116), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT22), .ZN(new_n590));
  AOI21_X1  g0390(.A(G20), .B1(new_n408), .B2(new_n409), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(G87), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n208), .B(G87), .C1(new_n372), .C2(new_n373), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n589), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI211_X1 g0397(.A(KEYINPUT77), .B(new_n589), .C1(new_n592), .C2(new_n594), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(KEYINPUT24), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n591), .A2(new_n590), .A3(G87), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT77), .B1(new_n602), .B2(new_n589), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT24), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n259), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n585), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G250), .B(new_n263), .C1(new_n372), .C2(new_n373), .ZN(new_n607));
  AND2_X1   g0407(.A1(G257), .A2(G1698), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n372), .B2(new_n373), .ZN(new_n609));
  NAND2_X1  g0409(.A1(G33), .A2(G294), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT79), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT79), .A4(new_n610), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n268), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n447), .A2(new_n273), .A3(G264), .A4(new_n276), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n446), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n575), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n615), .A2(G190), .A3(new_n617), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT80), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n262), .A2(new_n608), .B1(G33), .B2(G294), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT79), .B1(new_n622), .B2(new_n607), .ZN(new_n623));
  INV_X1    g0423(.A(new_n614), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n269), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n617), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n627), .A2(KEYINPUT80), .A3(G190), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n606), .B1(new_n621), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n577), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n581), .A2(new_n582), .B1(new_n530), .B2(G107), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n598), .A2(KEYINPUT24), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n603), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n595), .A2(new_n596), .A3(new_n604), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n321), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(G169), .B1(new_n625), .B2(new_n626), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n615), .A2(G179), .A3(new_n617), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NOR4_X1   g0441(.A1(new_n437), .A2(new_n494), .A3(new_n630), .A4(new_n641), .ZN(G372));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n510), .A2(new_n527), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n532), .A2(new_n534), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n643), .B1(new_n646), .B2(new_n564), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n555), .A2(new_n395), .A3(new_n557), .ZN(new_n648));
  AOI21_X1  g0448(.A(G169), .B1(new_n555), .B2(new_n557), .ZN(new_n649));
  NOR3_X1   g0449(.A1(new_n648), .A2(new_n649), .A3(new_n573), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n650), .A2(KEYINPUT26), .A3(new_n535), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n647), .A2(new_n651), .B1(new_n532), .B2(new_n534), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n491), .A2(new_n479), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n483), .A2(new_n653), .A3(new_n640), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n654), .B2(new_n630), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n436), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g0456(.A(new_n656), .B(KEYINPUT81), .Z(new_n657));
  INV_X1    g0457(.A(new_n293), .ZN(new_n658));
  INV_X1    g0458(.A(new_n351), .ZN(new_n659));
  INV_X1    g0459(.A(new_n314), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n353), .B2(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n432), .A2(new_n429), .A3(new_n416), .A4(new_n415), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n432), .B1(new_n383), .B2(new_n429), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n422), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n658), .B1(new_n665), .B2(new_n289), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n657), .A2(new_n666), .ZN(G369));
  AND2_X1   g0467(.A1(new_n483), .A2(new_n653), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  XOR2_X1   g0470(.A(new_n670), .B(KEYINPUT82), .Z(new_n671));
  INV_X1    g0471(.A(G213), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n669), .B2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(KEYINPUT83), .B(G343), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n479), .ZN(new_n679));
  OR3_X1    g0479(.A1(new_n668), .A2(KEYINPUT84), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n494), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n679), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT84), .B1(new_n668), .B2(new_n679), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT85), .Z(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n636), .B1(new_n639), .B2(new_n678), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n629), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n640), .A2(new_n677), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n483), .B1(new_n492), .B2(new_n493), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n693), .A2(new_n677), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n694), .A2(new_n688), .B1(new_n641), .B2(new_n677), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n211), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G41), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G1), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n506), .A2(G116), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n700), .A2(new_n701), .B1(new_n215), .B2(new_n699), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n646), .A2(new_n564), .A3(new_n643), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT26), .B1(new_n650), .B2(new_n535), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n645), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n577), .A2(new_n629), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n483), .B(new_n640), .C1(new_n492), .C2(new_n493), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n706), .A2(KEYINPUT87), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT87), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n652), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n678), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT88), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT29), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n706), .A2(KEYINPUT87), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n707), .A2(new_n708), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n677), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT88), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n655), .A2(new_n677), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n488), .B1(new_n457), .B2(new_n458), .ZN(new_n724));
  INV_X1    g0524(.A(new_n616), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n533), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n724), .A2(new_n563), .A3(new_n625), .A4(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n615), .A2(new_n725), .A3(new_n533), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n724), .A4(new_n563), .ZN(new_n731));
  INV_X1    g0531(.A(new_n563), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n526), .A2(G179), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n460), .A3(new_n627), .A4(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n678), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n678), .B1(new_n636), .B2(new_n639), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n577), .A2(new_n741), .A3(new_n629), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n681), .A2(KEYINPUT86), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT86), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n577), .A2(new_n741), .A3(new_n629), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n494), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n740), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G330), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n723), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n703), .B1(new_n751), .B2(G1), .ZN(G364));
  NOR2_X1   g0552(.A1(new_n328), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n700), .B1(G45), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n685), .B2(G330), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G330), .B2(new_n685), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n217), .B1(G20), .B2(new_n291), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n208), .A2(G179), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(G190), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT92), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n374), .B1(new_n765), .B2(G87), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT93), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT93), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n282), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n208), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n468), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n208), .A2(new_n395), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n772), .B1(new_n201), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n759), .A2(new_n282), .A3(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G107), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n773), .A2(G190), .A3(new_n575), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G190), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n780), .A2(G58), .B1(new_n783), .B2(G77), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n773), .A2(new_n282), .A3(G200), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n203), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT32), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n759), .A2(new_n781), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(KEYINPUT32), .A3(G159), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n786), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n767), .A2(new_n768), .A3(new_n778), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n774), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G326), .A2(new_n795), .B1(new_n777), .B2(G283), .ZN(new_n796));
  INV_X1    g0596(.A(G294), .ZN(new_n797));
  XOR2_X1   g0597(.A(KEYINPUT33), .B(G317), .Z(new_n798));
  OAI221_X1 g0598(.A(new_n796), .B1(new_n797), .B2(new_n770), .C1(new_n785), .C2(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n780), .A2(G322), .B1(new_n791), .B2(G329), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n800), .B(new_n374), .C1(new_n801), .C2(new_n782), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n764), .B(KEYINPUT94), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n805), .B2(new_n453), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n758), .B1(new_n794), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n754), .B(KEYINPUT89), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n211), .A2(new_n374), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(new_n439), .B2(new_n216), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n242), .B2(new_n439), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n697), .A2(new_n374), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n813), .A2(G355), .B1(new_n462), .B2(new_n697), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n815), .A2(KEYINPUT90), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G13), .A2(G33), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  XOR2_X1   g0619(.A(new_n819), .B(KEYINPUT91), .Z(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n757), .B(new_n821), .C1(new_n815), .C2(KEYINPUT90), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n807), .B(new_n809), .C1(new_n816), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT95), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n685), .B2(new_n820), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n756), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(G396));
  OAI21_X1  g0627(.A(new_n316), .B1(new_n312), .B2(new_n677), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n314), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n314), .A2(new_n678), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n720), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n832), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n655), .A2(new_n677), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n754), .B1(new_n750), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n750), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n757), .A2(new_n817), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n809), .B1(new_n221), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n374), .B1(new_n788), .B2(new_n801), .C1(new_n779), .C2(new_n797), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n772), .B1(new_n453), .B2(new_n774), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n841), .B(new_n842), .C1(G87), .C2(new_n777), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n785), .A2(new_n844), .B1(new_n782), .B2(new_n462), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT96), .Z(new_n846));
  OAI211_X1 g0646(.A(new_n843), .B(new_n846), .C1(new_n805), .C2(new_n505), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n805), .A2(new_n201), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n780), .A2(G143), .B1(new_n783), .B2(G159), .ZN(new_n849));
  INV_X1    g0649(.A(G137), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n850), .B2(new_n774), .C1(new_n254), .C2(new_n785), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  OR2_X1    g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI221_X1 g0655(.A(new_n262), .B1(new_n788), .B2(new_n855), .C1(new_n203), .C2(new_n776), .ZN(new_n856));
  INV_X1    g0656(.A(new_n770), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(G58), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n847), .B1(new_n848), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n757), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n840), .B(new_n861), .C1(new_n834), .C2(new_n818), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n838), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  OR2_X1    g0664(.A1(new_n570), .A2(KEYINPUT35), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n570), .A2(KEYINPUT35), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n865), .A2(new_n866), .A3(G116), .A4(new_n218), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT97), .B(KEYINPUT36), .Z(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n216), .A2(G77), .A3(new_n362), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n201), .A2(G68), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n207), .B(G13), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n678), .A2(new_n334), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n351), .A2(new_n353), .A3(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n334), .B(new_n678), .C1(new_n349), .C2(new_n350), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n834), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n743), .A2(new_n746), .ZN(new_n879));
  INV_X1    g0679(.A(new_n740), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n383), .A2(new_n674), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(new_n422), .B2(new_n434), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT98), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(KEYINPUT37), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n430), .A2(new_n888), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n402), .A2(new_n674), .B1(new_n415), .B2(new_n416), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n383), .A2(new_n429), .B1(new_n886), .B2(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(new_n887), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n417), .B1(new_n420), .B2(new_n675), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n882), .B1(new_n885), .B2(new_n896), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n889), .A2(new_n887), .A3(new_n890), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n893), .B1(new_n892), .B2(new_n894), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT18), .B1(new_n383), .B2(new_n402), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n417), .A2(new_n420), .A3(new_n404), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n883), .B1(new_n664), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n900), .A2(new_n904), .A3(KEYINPUT38), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n897), .A2(new_n905), .A3(KEYINPUT99), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT99), .B1(new_n897), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n881), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n897), .B2(new_n905), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n881), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n437), .A2(new_n747), .ZN(new_n914));
  OAI21_X1  g0714(.A(G330), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT100), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n914), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n916), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n897), .A2(new_n905), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT39), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n897), .A2(new_n905), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n659), .A2(new_n677), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT99), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n885), .A2(new_n896), .A3(new_n882), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT38), .B1(new_n900), .B2(new_n904), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n897), .A2(new_n905), .A3(KEYINPUT99), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n877), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n835), .B2(new_n831), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n903), .A2(new_n674), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n928), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n714), .A2(new_n719), .A3(new_n436), .A4(new_n722), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n666), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n920), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT101), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n207), .B2(new_n753), .C1(new_n942), .C2(new_n920), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n943), .A2(KEYINPUT101), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n873), .B1(new_n945), .B2(new_n946), .ZN(G367));
  NAND2_X1  g0747(.A1(new_n650), .A2(new_n678), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT103), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n564), .B(new_n576), .C1(new_n573), .C2(new_n677), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n692), .A2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n564), .B1(new_n952), .B2(new_n640), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n688), .A3(new_n694), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n955), .A2(new_n677), .B1(KEYINPUT42), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(KEYINPUT42), .B2(new_n956), .ZN(new_n958));
  OR3_X1    g0758(.A1(new_n677), .A2(new_n645), .A3(new_n510), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT102), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n535), .B1(new_n510), .B2(new_n677), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(KEYINPUT102), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n958), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n968));
  OR3_X1    g0768(.A1(new_n954), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n954), .B1(new_n967), .B2(new_n968), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n698), .B(KEYINPUT41), .Z(new_n971));
  MUX2_X1   g0771(.A(new_n690), .B(new_n688), .S(new_n694), .Z(new_n972));
  XOR2_X1   g0772(.A(new_n686), .B(new_n972), .Z(new_n973));
  OR3_X1    g0773(.A1(new_n695), .A2(KEYINPUT44), .A3(new_n951), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT44), .B1(new_n695), .B2(new_n951), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n695), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT45), .B1(new_n695), .B2(new_n951), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n691), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n691), .A2(new_n978), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n973), .A2(new_n979), .A3(new_n751), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n971), .B1(new_n981), .B2(new_n751), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n753), .A2(G45), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(G1), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n969), .B(new_n970), .C1(new_n982), .C2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n262), .B1(new_n788), .B2(new_n850), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n776), .A2(new_n221), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G143), .B2(new_n795), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n789), .B2(new_n785), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n986), .B(new_n989), .C1(G50), .C2(new_n783), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n202), .B2(new_n764), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n770), .A2(new_n203), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(G150), .B2(new_n780), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT109), .Z(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT46), .B1(new_n765), .B2(G116), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT107), .Z(new_n996));
  NAND3_X1  g0796(.A1(new_n804), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  INV_X1    g0797(.A(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n374), .B1(new_n788), .B2(new_n998), .C1(new_n468), .C2(new_n776), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(KEYINPUT108), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n857), .A2(G107), .B1(new_n783), .B2(G283), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(KEYINPUT105), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT106), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n779), .A2(new_n453), .B1(new_n774), .B2(new_n801), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n1001), .A2(KEYINPUT105), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT108), .B2(new_n999), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n785), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1004), .A2(new_n1003), .B1(G294), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n997), .A2(new_n1002), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n991), .A2(new_n994), .B1(new_n996), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT47), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n758), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n821), .A2(new_n757), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n238), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1014), .B1(new_n211), .B2(new_n301), .C1(new_n1015), .C2(new_n810), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n808), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT104), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1013), .B(new_n1018), .C1(new_n820), .C2(new_n963), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n985), .A2(new_n1019), .ZN(G387));
  OAI22_X1  g0820(.A1(new_n782), .A2(new_n203), .B1(new_n788), .B2(new_n254), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n374), .B(new_n1021), .C1(G50), .C2(new_n780), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n765), .A2(G77), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n305), .A2(new_n1007), .B1(new_n777), .B2(G97), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n770), .A2(new_n301), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G159), .B2(new_n795), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n262), .B1(new_n791), .B2(G326), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n764), .A2(new_n797), .B1(new_n844), .B2(new_n770), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n780), .A2(G317), .B1(new_n783), .B2(G303), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n795), .A2(G322), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(new_n801), .C2(new_n785), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT48), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1029), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT49), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1028), .B1(new_n462), .B2(new_n776), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1027), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n757), .ZN(new_n1040));
  AOI211_X1 g0840(.A(G45), .B(new_n701), .C1(G68), .C2(G77), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n252), .A2(G50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n810), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n235), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1044), .B1(new_n1045), .B2(new_n439), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n813), .A2(new_n701), .B1(new_n505), .B2(new_n697), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT110), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n809), .B1(new_n1049), .B2(new_n1014), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1040), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n690), .B2(new_n821), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n973), .B2(new_n984), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n973), .A2(new_n751), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n698), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n973), .A2(new_n751), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1053), .B1(new_n1055), .B2(new_n1056), .ZN(G393));
  NAND3_X1  g0857(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n245), .A2(new_n810), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1014), .B1(new_n468), .B2(new_n211), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n808), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n779), .A2(new_n789), .B1(new_n774), .B2(new_n254), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n765), .A2(G68), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n770), .A2(new_n221), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G87), .B2(new_n777), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n791), .A2(G143), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n374), .B1(new_n783), .B2(new_n305), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1007), .A2(G50), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n765), .A2(G283), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n374), .B1(new_n782), .B2(new_n797), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(G322), .B2(new_n791), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1007), .A2(G303), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n857), .A2(G116), .B1(new_n777), .B2(G107), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n779), .A2(new_n801), .B1(new_n774), .B2(new_n998), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT52), .Z(new_n1080));
  OAI22_X1  g0880(.A1(new_n1066), .A2(new_n1072), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1061), .B1(new_n1081), .B2(new_n757), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n951), .B2(new_n820), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1058), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT112), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n979), .A2(new_n980), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1054), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n698), .A3(new_n981), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(G390));
  INV_X1    g0890(.A(new_n839), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n808), .B1(new_n305), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(G125), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n262), .B1(new_n788), .B2(new_n1093), .C1(new_n779), .C2(new_n855), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT54), .B(G143), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n785), .A2(new_n850), .B1(new_n782), .B2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT114), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n776), .A2(new_n201), .ZN(new_n1098));
  INV_X1    g0898(.A(G128), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n770), .A2(new_n789), .B1(new_n774), .B2(new_n1099), .ZN(new_n1100));
  OR4_X1    g0900(.A1(new_n1094), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n765), .A2(G150), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT53), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n805), .A2(new_n387), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n774), .A2(new_n844), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1105), .B(new_n1067), .C1(G107), .C2(new_n1007), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n374), .B1(new_n782), .B2(new_n468), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G116), .B2(new_n780), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n776), .A2(new_n203), .B1(new_n788), .B2(new_n797), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT115), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1101), .A2(new_n1103), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1092), .B1(new_n1112), .B2(new_n757), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n925), .B2(new_n818), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n921), .A2(new_n926), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n830), .B1(new_n712), .B2(new_n829), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1116), .B1(new_n1117), .B2(new_n935), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n922), .B(new_n924), .C1(new_n936), .C2(new_n927), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n747), .A2(new_n748), .A3(new_n832), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT113), .B1(new_n1120), .B2(new_n877), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT86), .B1(new_n681), .B2(new_n742), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n494), .A2(new_n745), .A3(new_n744), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n880), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(G330), .A3(new_n834), .A4(new_n877), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT113), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1118), .B(new_n1119), .C1(new_n1121), .C2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n835), .A2(new_n831), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n927), .B1(new_n1130), .B2(new_n877), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n925), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n717), .A2(new_n677), .A3(new_n829), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n831), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1115), .B1(new_n1134), .B2(new_n877), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1129), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1128), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n984), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1114), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1124), .A2(G330), .A3(new_n834), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1134), .B1(new_n935), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n935), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1125), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1130), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n750), .A2(new_n437), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n941), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n699), .B1(new_n1149), .B2(new_n1137), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1146), .A2(new_n1148), .A3(new_n1128), .A4(new_n1136), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1139), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(G378));
  INV_X1    g0953(.A(new_n939), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT40), .B1(new_n934), .B2(new_n881), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n912), .A2(G330), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n289), .B2(new_n293), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n289), .A2(new_n293), .A3(new_n1158), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1160), .A2(new_n260), .A3(new_n675), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n260), .A2(new_n675), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1161), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n1159), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1155), .A2(new_n1156), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1166), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n748), .B1(new_n881), .B2(new_n911), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n910), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1154), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1166), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n910), .A2(new_n1169), .A3(new_n1168), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n939), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1171), .A2(KEYINPUT119), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .A4(new_n939), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1120), .A2(KEYINPUT113), .A3(new_n877), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1180), .A2(new_n1141), .B1(new_n1144), .B2(new_n1130), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1148), .B1(new_n1137), .B2(new_n1181), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1175), .A2(KEYINPUT57), .A3(new_n1177), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT120), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT57), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n1151), .B2(new_n1148), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT120), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1177), .A4(new_n1175), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1182), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n699), .B1(new_n1190), .B2(new_n1185), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1184), .A2(new_n1188), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1168), .A2(new_n817), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n374), .A2(new_n441), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1194), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n785), .A2(new_n468), .B1(new_n776), .B2(new_n202), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n992), .B(new_n1196), .C1(G116), .C2(new_n795), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1194), .B1(G283), .B2(new_n791), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n780), .A2(G107), .B1(new_n783), .B2(new_n302), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1197), .A2(new_n1023), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1195), .B1(new_n1201), .B2(KEYINPUT58), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n795), .A2(G125), .B1(new_n783), .B2(G137), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G150), .A2(new_n857), .B1(new_n1007), .B2(G132), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n764), .A2(new_n1095), .B1(new_n1099), .B2(new_n779), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1205), .A2(KEYINPUT116), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(KEYINPUT116), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1203), .B(new_n1204), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT117), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(G124), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(G124), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n791), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G33), .A2(G41), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n789), .C2(new_n776), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1208), .B2(KEYINPUT59), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1209), .A2(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1202), .B(new_n1217), .C1(KEYINPUT58), .C2(new_n1201), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1218), .A2(new_n758), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT118), .Z(new_n1220));
  OAI21_X1  g1020(.A(new_n754), .B1(G50), .B2(new_n1091), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1189), .A2(new_n984), .B1(new_n1193), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1192), .A2(new_n1223), .ZN(G375));
  OAI21_X1  g1024(.A(new_n1181), .B1(new_n941), .B2(new_n1147), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n971), .B(KEYINPUT121), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1225), .A2(new_n1149), .A3(new_n1226), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n804), .A2(G97), .B1(G303), .B2(new_n791), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT122), .Z(new_n1229));
  OAI221_X1 g1029(.A(new_n374), .B1(new_n782), .B2(new_n505), .C1(new_n844), .C2(new_n779), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n785), .A2(new_n462), .B1(new_n774), .B2(new_n797), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n987), .A4(new_n1025), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n804), .A2(G159), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n770), .A2(new_n201), .B1(new_n774), .B2(new_n855), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n785), .A2(new_n1095), .B1(new_n776), .B2(new_n202), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n262), .B1(new_n779), .B2(new_n850), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n782), .A2(new_n254), .B1(new_n788), .B2(new_n1099), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1229), .A2(new_n1232), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n808), .B1(G68), .B2(new_n1091), .C1(new_n1239), .C2(new_n758), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(new_n935), .B2(new_n817), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1146), .B2(new_n984), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1227), .A2(new_n1242), .ZN(G381));
  NAND4_X1  g1043(.A1(new_n985), .A2(new_n1086), .A3(new_n1019), .A4(new_n1089), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n826), .B(new_n1053), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1245));
  OR3_X1    g1045(.A1(new_n1245), .A2(G384), .A3(G381), .ZN(new_n1246));
  OR4_X1    g1046(.A1(G378), .A2(new_n1244), .A3(new_n1246), .A4(G375), .ZN(G407));
  NOR2_X1   g1047(.A1(new_n676), .A2(new_n672), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1152), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G375), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT123), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1250), .B(new_n1251), .ZN(G409));
  NAND2_X1  g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT125), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1245), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1244), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n985), .A2(new_n1019), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(G390), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1255), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1254), .B1(new_n1253), .B2(new_n1245), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1259), .B(new_n1244), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(KEYINPUT126), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1258), .A2(new_n1262), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT60), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n698), .B(new_n1149), .C1(new_n1225), .C2(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1225), .A2(new_n1269), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1242), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1272), .A2(new_n863), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n863), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1248), .A2(G2897), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1275), .B(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1175), .A2(new_n984), .A3(new_n1177), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1222), .A2(new_n1193), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1226), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1278), .B(new_n1279), .C1(new_n1190), .C2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1152), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1192), .A2(G378), .A3(new_n1223), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(KEYINPUT124), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT124), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1192), .A2(new_n1286), .A3(G378), .A4(new_n1223), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1283), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1277), .B1(new_n1288), .B2(new_n1248), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1288), .A2(new_n1248), .A3(new_n1275), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT62), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1268), .B(new_n1289), .C1(new_n1290), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1282), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1248), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1275), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1267), .B1(new_n1292), .B2(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1289), .A2(new_n1268), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT63), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1290), .A2(KEYINPUT63), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1300), .A2(new_n1302), .A3(new_n1303), .A4(new_n1263), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(G405));
  NAND2_X1  g1105(.A1(G375), .A2(new_n1152), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1275), .B1(new_n1293), .B2(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1293), .A2(new_n1275), .A3(new_n1306), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1267), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1307), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(G402));
endmodule


