//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  XNOR2_X1  g001(.A(G143), .B(G146), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n191), .A3(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n192), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(KEYINPUT0), .A2(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n189), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n190), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n203), .A2(G134), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT11), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n210), .B1(new_n205), .B2(G137), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n213));
  AOI211_X1 g027(.A(G131), .B(new_n207), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n211), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n204), .A2(new_n206), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n202), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NOR3_X1   g035(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n223));
  INV_X1    g037(.A(G113), .ZN(new_n224));
  OAI22_X1  g038(.A1(new_n221), .A2(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(G116), .B(G119), .Z(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G116), .B(G119), .ZN(new_n228));
  OAI221_X1 g042(.A(new_n228), .B1(new_n223), .B2(new_n224), .C1(new_n221), .C2(new_n222), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n233));
  AOI211_X1 g047(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n203), .C2(G134), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n217), .B(new_n215), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n208), .A2(new_n206), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n194), .A2(new_n196), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n193), .A2(G143), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  OAI21_X1  g057(.A(G128), .B1(new_n192), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G128), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(new_n240), .B2(KEYINPUT1), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT66), .B1(new_n197), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n246), .A2(KEYINPUT1), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n188), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n238), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n187), .B1(new_n232), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n217), .B1(new_n233), .B2(new_n234), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n235), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n230), .B1(new_n256), .B2(new_n202), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n242), .B1(new_n241), .B2(new_n244), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n197), .A2(KEYINPUT66), .A3(new_n247), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n251), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n238), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n257), .A2(new_n262), .A3(KEYINPUT68), .ZN(new_n263));
  NOR2_X1   g077(.A1(G237), .A2(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G210), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT27), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n253), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n253), .A2(new_n263), .A3(KEYINPUT69), .A4(new_n268), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT30), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n262), .B2(new_n219), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n201), .B1(new_n255), .B2(new_n235), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n252), .A2(KEYINPUT30), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n230), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT31), .B1(new_n271), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n230), .B1(new_n252), .B2(new_n275), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n253), .A2(new_n263), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT28), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT28), .B1(new_n257), .B2(new_n262), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n268), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n269), .A2(new_n270), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n272), .A4(new_n277), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(new_n287), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n262), .A2(new_n273), .A3(new_n219), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT30), .B1(new_n252), .B2(new_n275), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n231), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n253), .A2(new_n263), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n286), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT70), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n282), .A2(new_n268), .A3(new_n284), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n305), .B(new_n286), .C1(new_n299), .C2(new_n300), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT71), .B(G902), .Z(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI211_X1 g123(.A(new_n286), .B(new_n283), .C1(new_n281), .C2(KEYINPUT28), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n295), .A2(new_n296), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT25), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT77), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT77), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n320), .A2(new_n321), .A3(G146), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n317), .A2(new_n319), .A3(new_n323), .A4(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(new_n316), .A3(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(new_n328), .B2(KEYINPUT16), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n322), .B1(new_n330), .B2(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n246), .A2(G119), .ZN(new_n332));
  INV_X1    g146(.A(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G128), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .A4(KEYINPUT23), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT72), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(KEYINPUT23), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n338), .A2(new_n339), .A3(G119), .A4(new_n246), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT74), .B(G110), .Z(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n332), .A2(new_n334), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT76), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n343), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT75), .B1(new_n341), .B2(new_n342), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n331), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G137), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G953), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(G221), .A3(G234), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n355), .B(new_n357), .Z(new_n358));
  OAI21_X1  g172(.A(new_n193), .B1(new_n327), .B2(new_n329), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n317), .A2(new_n319), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT73), .B1(new_n360), .B2(new_n325), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(G146), .A3(new_n324), .A4(new_n326), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n344), .A2(new_n345), .ZN(new_n364));
  INV_X1    g178(.A(new_n341), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n365), .B2(G110), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n352), .A2(new_n358), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n358), .B1(new_n352), .B2(new_n367), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n315), .B(new_n308), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(new_n308), .B2(G234), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n352), .A2(new_n367), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n355), .B(new_n357), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n352), .A2(new_n358), .A3(new_n367), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n315), .B1(new_n378), .B2(new_n308), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT79), .B1(new_n373), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n308), .B1(new_n368), .B2(new_n369), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT25), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n370), .A4(new_n372), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT80), .B1(new_n376), .B2(new_n377), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n372), .A2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n380), .B(new_n384), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n320), .A2(new_n321), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT19), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n397), .B2(new_n360), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n193), .ZN(new_n400));
  INV_X1    g214(.A(G237), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n356), .A3(G214), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G143), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n264), .B(G214), .C1(new_n403), .C2(G143), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT92), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n215), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n406), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT92), .B1(new_n410), .B2(G131), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(G131), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n413), .A3(new_n362), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n407), .A2(new_n215), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n360), .A2(G146), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n396), .B2(G146), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n407), .B1(new_n419), .B2(new_n215), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n395), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT17), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n409), .B(new_n425), .C1(new_n411), .C2(new_n412), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n415), .A2(KEYINPUT17), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n363), .A2(KEYINPUT93), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT93), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n359), .A2(new_n362), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n424), .B1(new_n428), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT94), .B1(new_n433), .B2(new_n395), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n359), .A2(new_n362), .A3(new_n430), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n430), .B1(new_n359), .B2(new_n362), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n426), .B(new_n427), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(KEYINPUT94), .A3(new_n395), .A4(new_n421), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n423), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n395), .A3(new_n421), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n422), .B1(new_n446), .B2(new_n438), .ZN(new_n447));
  INV_X1    g261(.A(new_n442), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT20), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n395), .B1(new_n437), .B2(new_n421), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n446), .B2(new_n438), .ZN(new_n452));
  OAI21_X1  g266(.A(G475), .B1(new_n452), .B2(G902), .ZN(new_n453));
  NAND2_X1  g267(.A1(G234), .A2(G237), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n454), .A2(G952), .A3(new_n356), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n309), .A2(G953), .A3(new_n454), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT98), .Z(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(G898), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT99), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G478), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT97), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n191), .A2(G128), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n246), .A2(G143), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n464), .A2(new_n465), .A3(new_n205), .ZN(new_n466));
  INV_X1    g280(.A(G116), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G122), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n467), .A2(G122), .ZN(new_n470));
  OR3_X1    g284(.A1(new_n469), .A2(G107), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(G107), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT95), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n464), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n476), .B(new_n465), .C1(new_n475), .C2(new_n464), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n464), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g292(.A(G134), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G107), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n468), .B1(new_n470), .B2(KEYINPUT14), .ZN(new_n482));
  OR2_X1    g296(.A1(new_n482), .A2(KEYINPUT96), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n468), .A2(KEYINPUT14), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n484), .B1(new_n482), .B2(KEYINPUT96), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n205), .B1(new_n464), .B2(new_n465), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n471), .B1(new_n466), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n480), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT9), .B(G234), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n490), .A2(new_n371), .A3(G953), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n480), .B(new_n491), .C1(new_n486), .C2(new_n488), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n463), .B1(new_n495), .B2(new_n308), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT97), .B(new_n309), .C1(new_n493), .C2(new_n494), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n462), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n495), .A2(new_n308), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(KEYINPUT15), .B2(new_n461), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n460), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n450), .A2(new_n453), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G214), .B1(G237), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT3), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n481), .A3(G104), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n394), .A2(G107), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT4), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(G101), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT82), .B(G101), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n514), .A2(new_n508), .A3(new_n509), .A4(new_n506), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(KEYINPUT4), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n230), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n467), .A2(G119), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT5), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n224), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n226), .B2(new_n519), .ZN(new_n521));
  INV_X1    g335(.A(new_n509), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n394), .A2(G107), .ZN(new_n523));
  OAI21_X1  g337(.A(G101), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n229), .A2(new_n521), .A3(new_n515), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(G110), .B(G122), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n517), .A2(new_n527), .A3(new_n525), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n529), .A2(KEYINPUT6), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n202), .A2(G125), .ZN(new_n532));
  INV_X1    g346(.A(new_n251), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n245), .B2(new_n248), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n532), .B1(new_n534), .B2(G125), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT87), .ZN(new_n536));
  INV_X1    g350(.A(G224), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n536), .B1(new_n537), .B2(G953), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n356), .A2(KEYINPUT87), .A3(G224), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT86), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n532), .B(new_n541), .C1(new_n534), .C2(G125), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n526), .A2(new_n546), .A3(new_n528), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n531), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n532), .B(new_n553), .C1(new_n534), .C2(G125), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT90), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n527), .B(KEYINPUT8), .ZN(new_n556));
  AND4_X1   g370(.A1(new_n229), .A2(new_n521), .A3(new_n515), .A4(new_n524), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n229), .A2(new_n521), .B1(new_n515), .B2(new_n524), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT89), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n229), .A2(new_n521), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n515), .A2(new_n524), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(new_n525), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n556), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n517), .A2(new_n525), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n560), .A2(new_n566), .B1(new_n527), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n535), .A2(KEYINPUT7), .A3(new_n552), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n555), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n531), .A2(new_n545), .A3(KEYINPUT88), .A4(new_n547), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n550), .A2(new_n551), .A3(new_n570), .A4(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G210), .B1(G237), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n559), .A2(KEYINPUT89), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n565), .B1(new_n564), .B2(new_n556), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n530), .B(new_n569), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n579), .B2(new_n555), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n580), .A2(new_n573), .A3(new_n571), .A4(new_n550), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n505), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G221), .B1(new_n490), .B2(G902), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XOR2_X1   g398(.A(KEYINPUT85), .B(KEYINPUT10), .Z(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n188), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n244), .A3(KEYINPUT84), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT84), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n247), .B2(new_n188), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n188), .A2(KEYINPUT83), .A3(new_n250), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT83), .B1(new_n188), .B2(new_n250), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n588), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n562), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n202), .A2(new_n516), .A3(new_n512), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(KEYINPUT10), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n534), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n214), .A2(new_n218), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n534), .A2(new_n562), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n593), .A2(new_n594), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT12), .B1(new_n605), .B2(new_n256), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT12), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n607), .B(new_n601), .C1(new_n603), .C2(new_n604), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n602), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(G110), .B(G140), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT81), .ZN(new_n611));
  INV_X1    g425(.A(G227), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(G953), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n611), .B(new_n613), .Z(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n599), .A2(new_n595), .A3(new_n596), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n616), .B2(new_n601), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n597), .A2(new_n600), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n256), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n609), .A2(new_n615), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G469), .B1(new_n620), .B2(G902), .ZN(new_n621));
  INV_X1    g435(.A(G469), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n606), .A2(new_n608), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n602), .A2(new_n614), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n614), .B1(new_n619), .B2(new_n602), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n622), .B(new_n308), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n584), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n582), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n314), .A2(new_n392), .A3(new_n503), .A4(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(new_n514), .Z(G3));
  AOI21_X1  g445(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n447), .A2(KEYINPUT20), .A3(new_n448), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n453), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n493), .B2(KEYINPUT100), .ZN(new_n636));
  OR2_X1    g450(.A1(new_n636), .A2(new_n495), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n495), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(G478), .A3(new_n308), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n496), .A2(new_n497), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(G478), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n634), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n575), .A2(new_n581), .ZN(new_n645));
  INV_X1    g459(.A(new_n460), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n504), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G472), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n291), .B2(new_n308), .ZN(new_n650));
  INV_X1    g464(.A(new_n292), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n288), .A2(new_n272), .A3(new_n277), .ZN(new_n652));
  AOI22_X1  g466(.A1(new_n652), .A2(KEYINPUT31), .B1(new_n285), .B2(new_n286), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n653), .B2(new_n290), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n650), .A2(new_n654), .A3(new_n391), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n648), .A2(new_n655), .A3(new_n628), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G6));
  NAND2_X1  g472(.A1(new_n453), .A2(KEYINPUT102), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n498), .A2(new_n500), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n662), .B(G475), .C1(new_n452), .C2(G902), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n450), .A2(new_n659), .A3(new_n661), .A4(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n647), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n655), .A3(new_n628), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT103), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT35), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G107), .ZN(G9));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n375), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT104), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(new_n374), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n374), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n389), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n380), .A2(new_n675), .A3(new_n384), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n650), .A2(new_n654), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n629), .A3(new_n679), .A4(new_n503), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n455), .B1(new_n457), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n664), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n314), .A2(new_n685), .A3(new_n678), .A4(new_n629), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  NAND2_X1  g503(.A1(new_n621), .A2(new_n627), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n583), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n684), .B(KEYINPUT39), .Z(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n645), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n281), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n652), .B1(new_n268), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n649), .B1(new_n701), .B2(new_n551), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n295), .A2(new_n296), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n695), .A2(KEYINPUT40), .ZN(new_n705));
  INV_X1    g519(.A(new_n634), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n706), .A2(new_n660), .A3(new_n505), .A4(new_n676), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n699), .A2(new_n704), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  INV_X1    g523(.A(new_n684), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n634), .A2(new_n643), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n314), .A2(new_n678), .A3(new_n711), .A4(new_n629), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G146), .ZN(G48));
  NOR2_X1   g527(.A1(new_n625), .A2(new_n626), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(new_n309), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n583), .A3(new_n627), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n648), .A2(new_n314), .A3(new_n392), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT108), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n665), .A2(new_n314), .A3(new_n392), .A4(new_n717), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NAND2_X1  g537(.A1(new_n645), .A2(new_n504), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(new_n716), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n314), .A2(new_n725), .A3(new_n678), .A4(new_n503), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  AND3_X1   g541(.A1(new_n582), .A2(new_n634), .A3(new_n661), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n716), .A2(new_n460), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n655), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G122), .ZN(G24));
  NAND4_X1  g545(.A1(new_n725), .A2(new_n711), .A3(new_n679), .A4(new_n676), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  NAND3_X1  g547(.A1(new_n575), .A2(new_n581), .A3(new_n504), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n691), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n314), .A2(new_n392), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT109), .A3(new_n711), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n314), .A2(new_n711), .A3(new_n392), .A4(new_n735), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT110), .B(KEYINPUT42), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n737), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n711), .A2(new_n735), .A3(KEYINPUT42), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n296), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n291), .A2(KEYINPUT111), .A3(KEYINPUT32), .A4(new_n292), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n746), .A2(new_n295), .A3(new_n313), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT112), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n392), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n749), .B1(new_n748), .B2(new_n392), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n744), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n743), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G131), .ZN(G33));
  INV_X1    g569(.A(new_n664), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n757), .A3(new_n710), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT113), .B1(new_n664), .B2(new_n684), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n736), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NAND2_X1  g576(.A1(new_n706), .A2(new_n643), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(KEYINPUT43), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n676), .B1(new_n650), .B2(new_n654), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n734), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  INV_X1    g589(.A(new_n627), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n620), .B(KEYINPUT45), .Z(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n777), .B2(G902), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n776), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(KEYINPUT46), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n583), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n693), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n774), .A2(new_n775), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  XNOR2_X1  g598(.A(new_n781), .B(KEYINPUT47), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n711), .A2(new_n391), .A3(new_n770), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(new_n314), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  INV_X1    g603(.A(new_n704), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n716), .A2(new_n734), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n392), .A3(new_n455), .A4(new_n791), .ZN(new_n792));
  OAI211_X1 g606(.A(G952), .B(new_n356), .C1(new_n792), .C2(new_n644), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n764), .A2(new_n455), .A3(new_n765), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n655), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n724), .A3(new_n716), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT119), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT119), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n794), .A2(new_n791), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n748), .A2(new_n392), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT112), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n750), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT48), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT120), .ZN(new_n807));
  INV_X1    g621(.A(new_n715), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n776), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n584), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n785), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n795), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n770), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n698), .A2(new_n505), .A3(new_n717), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n795), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT50), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n792), .A2(new_n634), .A3(new_n643), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n679), .A2(new_n676), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n817), .B1(new_n800), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n813), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n807), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n738), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n741), .B1(new_n826), .B2(KEYINPUT109), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n827), .A2(new_n740), .B1(new_n803), .B2(new_n744), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n630), .A2(new_n680), .A3(new_n730), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n726), .A2(new_n656), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n450), .A2(new_n659), .A3(new_n660), .A4(new_n663), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n314), .A2(new_n678), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n679), .A2(new_n634), .A3(new_n643), .A4(new_n676), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n691), .A2(new_n734), .A3(new_n684), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n835), .A2(new_n836), .B1(new_n736), .B2(new_n760), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n460), .B(new_n505), .C1(new_n575), .C2(new_n581), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n706), .A3(KEYINPUT115), .A4(new_n661), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n450), .A2(new_n453), .A3(new_n661), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n647), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n839), .A2(new_n842), .A3(new_n628), .A4(new_n655), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n843), .A2(new_n718), .A3(new_n722), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n831), .A2(new_n837), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT116), .B1(new_n828), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n676), .A2(new_n684), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT117), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n628), .A3(new_n704), .A4(new_n728), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n712), .A2(new_n732), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n686), .A2(new_n687), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n686), .A2(new_n687), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n688), .A2(KEYINPUT52), .A3(new_n849), .A4(new_n850), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n843), .A2(new_n718), .A3(new_n722), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n829), .A3(new_n830), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n754), .A2(new_n858), .A3(new_n860), .A4(new_n837), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n846), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n846), .A2(new_n857), .A3(new_n861), .A4(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n864), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n828), .A2(new_n845), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n857), .A2(new_n872), .A3(KEYINPUT53), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n825), .A2(new_n875), .B1(G952), .B2(G953), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n809), .B(KEYINPUT49), .Z(new_n877));
  NOR4_X1   g691(.A1(new_n877), .A2(new_n391), .A3(new_n584), .A4(new_n505), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n706), .A3(new_n643), .A4(new_n698), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n876), .B1(new_n704), .B2(new_n879), .ZN(G75));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n308), .B1(new_n870), .B2(new_n873), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT56), .B1(new_n882), .B2(new_n574), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n531), .A2(new_n547), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n545), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n356), .A2(G952), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n883), .B2(new_n886), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n881), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n883), .A2(new_n886), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(KEYINPUT121), .A3(new_n887), .A4(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(G51));
  NAND3_X1  g709(.A1(new_n882), .A2(G469), .A3(new_n777), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT122), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n870), .A2(new_n873), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n874), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(G469), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT57), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n901), .A2(new_n903), .B1(new_n626), .B2(new_n625), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n889), .B1(new_n897), .B2(new_n904), .ZN(G54));
  AND3_X1   g719(.A1(new_n882), .A2(KEYINPUT58), .A3(G475), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n890), .B1(new_n906), .B2(new_n440), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n440), .B2(new_n906), .ZN(G60));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n639), .B1(new_n875), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n637), .B2(new_n638), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n900), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n890), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT123), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n889), .B1(new_n900), .B2(new_n913), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n910), .B1(new_n869), .B2(new_n874), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n917), .B(new_n918), .C1(new_n919), .C2(new_n639), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n916), .A2(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT60), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n870), .B2(new_n873), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n673), .A2(new_n674), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n889), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n388), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n924), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT124), .B1(new_n924), .B2(new_n925), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(KEYINPUT61), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n928), .B(new_n930), .ZN(G66));
  OAI21_X1  g745(.A(G953), .B1(new_n459), .B2(new_n537), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n860), .B2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n884), .B1(G898), .B2(new_n356), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  NOR2_X1   g749(.A1(new_n356), .A2(G900), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n782), .A2(new_n728), .A3(new_n803), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n788), .A2(new_n761), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n688), .A2(new_n850), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n938), .A2(new_n754), .A3(new_n783), .A4(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n940), .B2(new_n356), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n298), .A2(new_n297), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n399), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n612), .B2(new_n683), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n939), .A2(new_n708), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  AOI211_X1 g763(.A(new_n734), .B(new_n695), .C1(new_n644), .C2(new_n841), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n392), .A3(new_n314), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT125), .Z(new_n952));
  NAND4_X1  g766(.A1(new_n949), .A2(new_n783), .A3(new_n788), .A4(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n943), .B1(new_n953), .B2(new_n356), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n945), .A2(new_n947), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n947), .B1(new_n945), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(G72));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT63), .Z(new_n959));
  INV_X1    g773(.A(new_n860), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n953), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n277), .A2(new_n253), .A3(new_n263), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n268), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n959), .B1(new_n940), .B2(new_n960), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n962), .A2(new_n268), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n889), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n867), .A2(new_n868), .ZN(new_n968));
  INV_X1    g782(.A(new_n959), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n302), .A2(new_n306), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n652), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n967), .B1(new_n968), .B2(new_n971), .ZN(G57));
endmodule


