//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT77), .ZN(new_n193));
  INV_X1    g007(.A(G953), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n194), .A2(G227), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n193), .B(new_n195), .Z(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT83), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT78), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G104), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n203), .A3(G104), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n207), .A2(new_n203), .A3(KEYINPUT79), .A4(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n206), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT4), .B1(new_n214), .B2(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(G101), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT80), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n202), .A2(new_n205), .B1(new_n210), .B2(new_n211), .ZN(new_n218));
  AOI21_X1  g032(.A(G101), .B1(new_n199), .B2(G107), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND4_X1   g034(.A1(new_n217), .A2(new_n206), .A3(new_n212), .A4(new_n219), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n215), .B1(new_n222), .B2(KEYINPUT4), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G143), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n231), .B(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n204), .A2(new_n213), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G101), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n206), .A2(new_n212), .A3(new_n219), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT80), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n218), .A2(new_n217), .A3(new_n219), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  AND4_X1   g057(.A1(new_n243), .A2(new_n226), .A3(new_n228), .A4(G128), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  OAI22_X1  g059(.A1(new_n245), .A2(G128), .B1(new_n243), .B2(new_n228), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI221_X1 g062(.A(KEYINPUT69), .B1(new_n243), .B2(new_n228), .C1(new_n245), .C2(G128), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT10), .ZN(new_n252));
  OAI22_X1  g066(.A1(new_n223), .A2(new_n234), .B1(new_n242), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT10), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n239), .A2(new_n240), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n236), .B1(new_n246), .B2(new_n244), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT81), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n259));
  AOI211_X1 g073(.A(new_n259), .B(new_n256), .C1(new_n239), .C2(new_n240), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n254), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT82), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n220), .B2(new_n221), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n259), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n255), .A2(KEYINPUT81), .A3(new_n257), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT82), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(new_n254), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n253), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G131), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G134), .ZN(new_n274));
  AOI21_X1  g088(.A(G137), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT66), .B1(new_n275), .B2(KEYINPUT11), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT66), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT65), .B(G134), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(G137), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g095(.A1(KEYINPUT67), .A2(G137), .ZN(new_n282));
  NAND2_X1  g096(.A1(KEYINPUT67), .A2(G137), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n282), .A2(KEYINPUT11), .A3(G134), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n272), .A2(new_n274), .A3(G137), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n270), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  AOI211_X1 g102(.A(G131), .B(new_n286), .C1(new_n276), .C2(new_n280), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n198), .B1(new_n269), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n242), .A2(new_n252), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n293));
  INV_X1    g107(.A(new_n215), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n231), .B(new_n233), .Z(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n267), .B1(new_n266), .B2(new_n254), .ZN(new_n298));
  AOI211_X1 g112(.A(KEYINPUT82), .B(KEYINPUT10), .C1(new_n264), .C2(new_n265), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n290), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(KEYINPUT83), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n290), .B(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n197), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(KEYINPUT84), .A3(new_n197), .ZN(new_n306));
  OAI22_X1  g120(.A1(new_n258), .A2(new_n260), .B1(new_n251), .B2(new_n241), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n301), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT12), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(KEYINPUT12), .A3(new_n301), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT84), .B1(new_n304), .B2(new_n197), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n190), .B(new_n191), .C1(new_n305), .C2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n190), .A2(new_n191), .ZN(new_n317));
  INV_X1    g131(.A(new_n304), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(new_n196), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n312), .A2(new_n304), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n303), .A2(new_n319), .B1(new_n196), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n317), .B1(new_n321), .B2(G469), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n189), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT90), .ZN(new_n326));
  NAND2_X1  g140(.A1(KEYINPUT18), .A2(G131), .ZN(new_n327));
  INV_X1    g141(.A(G237), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n194), .A3(G214), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n227), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n328), .A2(new_n194), .A3(G143), .A4(G214), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT87), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT87), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n334), .A3(new_n331), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n327), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G125), .B(G140), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(G146), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n330), .A2(new_n327), .A3(new_n331), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT88), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(KEYINPUT16), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n344), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n225), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(G146), .A3(new_n345), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(KEYINPUT17), .A3(G131), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n332), .A2(G131), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT17), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n330), .A2(new_n270), .A3(new_n331), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G113), .B(G122), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(new_n199), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n342), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n339), .A2(new_n341), .B1(new_n350), .B2(new_n354), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT89), .B1(new_n361), .B2(new_n357), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n361), .A2(new_n357), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n326), .B(new_n191), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n358), .A2(new_n359), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(KEYINPUT89), .A3(new_n357), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT90), .B1(new_n368), .B2(G902), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(new_n369), .A3(G475), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT20), .ZN(new_n371));
  NOR2_X1   g185(.A1(G475), .A2(G902), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n348), .B(KEYINPUT74), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n337), .B(KEYINPUT19), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n225), .A2(new_n374), .B1(new_n351), .B2(new_n353), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n357), .B1(new_n342), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n371), .B(new_n372), .C1(new_n363), .C2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n377), .B1(new_n366), .B2(new_n367), .ZN(new_n379));
  INV_X1    g193(.A(G475), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n191), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT20), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G952), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(G953), .ZN(new_n385));
  NAND2_X1  g199(.A1(G234), .A2(G237), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(G902), .A3(G953), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT21), .B(G898), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G143), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n227), .A2(G128), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n279), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n397), .A2(KEYINPUT92), .A3(new_n279), .A4(new_n398), .ZN(new_n402));
  XNOR2_X1  g216(.A(G116), .B(G122), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(new_n203), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n395), .B(KEYINPUT91), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT13), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n398), .B(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G134), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n401), .A2(new_n402), .A3(new_n404), .A4(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G122), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G116), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n203), .B1(new_n411), .B2(KEYINPUT14), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(new_n399), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n279), .B1(new_n397), .B2(new_n398), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n187), .A2(new_n418), .A3(G953), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n409), .A2(new_n416), .A3(new_n419), .ZN(new_n422));
  AOI21_X1  g236(.A(G902), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(KEYINPUT15), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n425), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n370), .A2(new_n383), .A3(new_n393), .A4(new_n429), .ZN(new_n430));
  MUX2_X1   g244(.A(new_n250), .B(new_n234), .S(G125), .Z(new_n431));
  INV_X1    g245(.A(G224), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(G953), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(G953), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n234), .A2(new_n344), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n250), .A2(G125), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT2), .B(G113), .Z(new_n440));
  XNOR2_X1  g254(.A(G116), .B(G119), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G119), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G116), .ZN(new_n447));
  OAI21_X1  g261(.A(G113), .B1(new_n447), .B2(KEYINPUT5), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n241), .B(new_n443), .C1(new_n445), .C2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n440), .B(new_n441), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n449), .B1(new_n223), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G122), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n449), .B(new_n454), .C1(new_n223), .C2(new_n451), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT6), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT4), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n255), .B2(new_n216), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n450), .B1(new_n460), .B2(new_n215), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n454), .B1(new_n461), .B2(new_n449), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n439), .B(new_n456), .C1(new_n458), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n452), .A2(new_n455), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n464), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n457), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n438), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n434), .A2(KEYINPUT7), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n431), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n454), .B(KEYINPUT8), .ZN(new_n470));
  INV_X1    g284(.A(new_n449), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n445), .A2(new_n448), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n241), .B1(new_n443), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n469), .B(new_n474), .C1(new_n438), .C2(new_n468), .ZN(new_n475));
  INV_X1    g289(.A(new_n457), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n191), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G210), .B1(G237), .B2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT86), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n467), .A2(new_n478), .A3(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT86), .B(new_n480), .C1(new_n466), .C2(new_n477), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n325), .B(new_n430), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n323), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n296), .B1(new_n288), .B2(new_n289), .ZN(new_n489));
  AOI21_X1  g303(.A(G134), .B1(new_n282), .B2(new_n283), .ZN(new_n490));
  OAI21_X1  g304(.A(G131), .B1(new_n490), .B2(new_n275), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT68), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n281), .A2(new_n270), .A3(new_n287), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n251), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT30), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n489), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n489), .B2(new_n495), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n450), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT70), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n450), .B(KEYINPUT71), .Z(new_n502));
  NAND3_X1  g316(.A1(new_n489), .A2(new_n495), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n328), .A2(new_n194), .A3(G210), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT27), .Z(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G101), .ZN(new_n506));
  XOR2_X1   g320(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n508), .B(new_n450), .C1(new_n498), .C2(new_n499), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n501), .A2(new_n503), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT31), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n509), .A2(new_n503), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n513), .A2(KEYINPUT31), .A3(new_n507), .A4(new_n501), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT28), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n503), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT72), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n503), .A2(KEYINPUT72), .A3(new_n515), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n489), .A2(new_n495), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n503), .B1(new_n522), .B2(new_n451), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT28), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n507), .ZN(new_n526));
  AOI22_X1  g340(.A1(new_n512), .A2(new_n514), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G472), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n191), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n488), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n509), .A2(new_n503), .ZN(new_n533));
  INV_X1    g347(.A(new_n499), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n497), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n508), .B1(new_n535), .B2(new_n450), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n526), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n520), .A2(new_n524), .A3(new_n507), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n522), .A2(new_n502), .ZN(new_n541));
  INV_X1    g355(.A(new_n503), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT28), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n526), .A2(new_n539), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n543), .A2(new_n519), .A3(new_n518), .A4(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n545), .A2(new_n191), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n528), .B1(new_n540), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n512), .A2(new_n514), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n525), .A2(new_n526), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n529), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n547), .B1(new_n550), .B2(KEYINPUT32), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT73), .B(new_n488), .C1(new_n527), .C2(new_n529), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n532), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n418), .B1(G234), .B2(new_n191), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n347), .A2(new_n348), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n394), .A2(G119), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT23), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n446), .A2(G128), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n394), .A2(KEYINPUT23), .A3(G119), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n557), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT24), .B(G110), .ZN(new_n564));
  OAI221_X1 g378(.A(new_n555), .B1(new_n556), .B2(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n556), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n564), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n566), .A2(new_n567), .B1(new_n225), .B2(new_n337), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n373), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n194), .A2(G221), .A3(G234), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT75), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n570), .A2(new_n574), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(G902), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT25), .ZN(new_n579));
  OAI211_X1 g393(.A(KEYINPUT25), .B(new_n191), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n554), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n554), .A2(G902), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(KEYINPUT76), .Z(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n575), .B2(new_n576), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n323), .A2(KEYINPUT93), .A3(new_n484), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n487), .A2(new_n553), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  INV_X1    g404(.A(new_n323), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n527), .B2(G902), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n529), .B2(new_n527), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n591), .A2(new_n586), .A3(new_n593), .ZN(new_n594));
  OR3_X1    g408(.A1(new_n423), .A2(KEYINPUT94), .A3(G478), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT94), .B1(new_n423), .B2(G478), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n421), .A2(new_n422), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT33), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n421), .A2(new_n599), .A3(new_n422), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n424), .A2(G902), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n595), .A2(new_n596), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n370), .B2(new_n383), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n479), .B1(new_n467), .B2(new_n478), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n466), .A2(new_n477), .A3(new_n480), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n325), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n594), .A2(new_n393), .A3(new_n604), .A4(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  OAI211_X1 g425(.A(new_n324), .B(new_n393), .C1(new_n605), .C2(new_n606), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n370), .A2(new_n383), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n428), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n594), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NOR2_X1   g432(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n570), .B(new_n619), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n584), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n582), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n593), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n487), .A2(new_n588), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT37), .B(G110), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G12));
  OAI211_X1 g441(.A(new_n622), .B(new_n324), .C1(new_n606), .C2(new_n605), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n389), .A2(G900), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n387), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n614), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n553), .A2(new_n629), .A3(new_n323), .A4(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT95), .B(G128), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G30));
  NAND2_X1  g450(.A1(new_n370), .A2(new_n383), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n324), .A3(new_n428), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n622), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(new_n639), .B(KEYINPUT96), .Z(new_n640));
  NAND2_X1  g454(.A1(new_n482), .A2(new_n483), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT38), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n631), .B(KEYINPUT39), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n323), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n646), .A2(KEYINPUT40), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(KEYINPUT40), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n507), .B1(new_n533), .B2(new_n536), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n541), .A2(new_n542), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n650), .B2(new_n526), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n528), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n550), .B2(KEYINPUT32), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n532), .A2(new_n653), .A3(new_n552), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n644), .A2(new_n647), .A3(new_n648), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n604), .A2(new_n657), .A3(new_n631), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n657), .B1(new_n604), .B2(new_n631), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n553), .A2(new_n629), .A3(new_n323), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  NAND2_X1  g476(.A1(new_n553), .A2(new_n587), .ZN(new_n663));
  INV_X1    g477(.A(new_n603), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n637), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n663), .A2(new_n665), .A3(new_n612), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n316), .A2(KEYINPUT98), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n318), .B1(new_n291), .B2(new_n302), .ZN(new_n668));
  OAI22_X1  g482(.A1(new_n668), .A2(new_n197), .B1(new_n313), .B2(new_n314), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n190), .B1(new_n669), .B2(new_n191), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AOI211_X1 g485(.A(KEYINPUT98), .B(new_n190), .C1(new_n669), .C2(new_n191), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n188), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(KEYINPUT99), .B(new_n188), .C1(new_n671), .C2(new_n672), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n666), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G15));
  XNOR2_X1  g493(.A(new_n667), .B(new_n670), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT99), .B1(new_n680), .B2(new_n188), .ZN(new_n681));
  INV_X1    g495(.A(new_n676), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n553), .A2(new_n587), .A3(new_n615), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NOR2_X1   g500(.A1(new_n628), .A2(new_n430), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n553), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  AOI21_X1  g504(.A(new_n507), .B1(new_n520), .B2(new_n543), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n512), .B2(new_n514), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n692), .A2(new_n529), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(new_n592), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n694), .A2(new_n587), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n607), .A2(new_n638), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n392), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n675), .A2(new_n676), .A3(new_n695), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT100), .B(G122), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G24));
  NAND4_X1  g515(.A1(new_n660), .A2(new_n693), .A3(new_n592), .A4(new_n622), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n675), .A2(new_n608), .A3(new_n676), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  NAND2_X1  g519(.A1(new_n530), .A2(KEYINPUT101), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT101), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n707), .B(new_n488), .C1(new_n527), .C2(new_n529), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n706), .A2(new_n551), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n587), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n641), .A2(new_n325), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n323), .A2(new_n660), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT42), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n323), .A2(new_n711), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n660), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n717), .A3(new_n553), .A4(new_n587), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n270), .ZN(G33));
  NAND4_X1  g534(.A1(new_n715), .A2(new_n553), .A3(new_n587), .A4(new_n633), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n637), .B2(KEYINPUT103), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n637), .A2(new_n603), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n613), .B(new_n664), .C1(new_n727), .C2(KEYINPUT43), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n593), .A3(new_n622), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n593), .A3(KEYINPUT44), .A4(new_n622), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n711), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n732), .A2(new_n733), .A3(new_n736), .A4(new_n711), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT46), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n321), .A2(KEYINPUT45), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n321), .B2(KEYINPUT45), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n303), .A2(new_n319), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n320), .A2(new_n196), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n190), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT102), .A3(new_n741), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n739), .B1(new_n751), .B2(new_n317), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n317), .B1(new_n744), .B2(new_n750), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n316), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n188), .A3(new_n645), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(new_n757), .B(G137), .Z(G39));
  INV_X1    g572(.A(new_n711), .ZN(new_n759));
  OR4_X1    g573(.A1(new_n553), .A2(new_n716), .A3(new_n587), .A4(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n754), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n316), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n188), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n760), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT105), .B(G140), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G42));
  INV_X1    g583(.A(new_n680), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT49), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT49), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n587), .A2(new_n188), .A3(new_n324), .A4(new_n725), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n654), .A2(new_n642), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT106), .Z(new_n776));
  NOR2_X1   g590(.A1(new_n759), .A2(new_n387), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n675), .A2(new_n676), .A3(new_n729), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n694), .A2(new_n622), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n654), .A2(new_n586), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n637), .A2(new_n664), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n683), .A2(new_n777), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n387), .B1(new_n726), .B2(new_n728), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n695), .A2(new_n784), .A3(new_n643), .A4(new_n325), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n681), .A2(new_n785), .A3(new_n682), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(KEYINPUT50), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n681), .A2(new_n785), .A3(new_n682), .A4(new_n788), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n780), .B(new_n783), .C1(new_n787), .C2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n680), .A2(new_n189), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT114), .A4(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n695), .A2(new_n784), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n711), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n765), .A2(new_n766), .A3(new_n794), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n793), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n792), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n799), .A2(new_n797), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n793), .B1(new_n804), .B2(new_n790), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n683), .A2(new_n608), .A3(new_n796), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n683), .A2(new_n777), .A3(new_n781), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n385), .B(new_n806), .C1(new_n807), .C2(new_n665), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n778), .B2(new_n710), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n778), .A2(new_n809), .A3(new_n710), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT48), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n809), .B(KEYINPUT48), .C1(new_n778), .C2(new_n710), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n805), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n622), .A2(new_n632), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n654), .A2(new_n696), .A3(new_n323), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n661), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n704), .A2(new_n634), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n704), .A2(new_n823), .A3(new_n634), .A4(new_n819), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n593), .A2(new_n586), .ZN(new_n827));
  AOI211_X1 g641(.A(new_n325), .B(new_n392), .C1(new_n482), .C2(new_n483), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n428), .B(KEYINPUT109), .Z(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n613), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n827), .A2(new_n323), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n625), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n675), .B(new_n676), .C1(new_n684), .C2(new_n688), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n834), .A2(new_n677), .A3(new_n835), .A4(new_n699), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT108), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n665), .B(KEYINPUT107), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n827), .A2(new_n323), .A3(new_n828), .A4(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n589), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n589), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n713), .A2(new_n718), .A3(new_n721), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT110), .ZN(new_n844));
  NOR4_X1   g658(.A1(new_n623), .A2(new_n637), .A3(new_n632), .A4(new_n829), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n553), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n714), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n715), .A2(KEYINPUT110), .A3(new_n553), .A4(new_n845), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n703), .A2(new_n715), .A3(KEYINPUT111), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT111), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n702), .B2(new_n714), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n847), .A2(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n836), .A2(new_n842), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n826), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n847), .A2(new_n848), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n849), .A2(new_n851), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n713), .A2(new_n718), .A3(new_n721), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n835), .A2(new_n699), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n589), .A2(new_n839), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT108), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n589), .A2(new_n837), .A3(new_n839), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n833), .B1(new_n683), .B2(new_n666), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n860), .A2(new_n861), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n824), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n855), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n826), .A2(new_n854), .A3(KEYINPUT53), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n870), .B1(new_n867), .B2(new_n869), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n803), .A2(new_n816), .A3(new_n872), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n384), .A2(new_n194), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n776), .B1(new_n880), .B2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n194), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n191), .B1(new_n873), .B2(new_n874), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n885), .B2(G210), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n463), .A2(new_n465), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n438), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n467), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  OAI21_X1  g705(.A(new_n884), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n886), .B2(new_n891), .ZN(G51));
  AND2_X1   g707(.A1(new_n885), .A2(new_n751), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n317), .B(KEYINPUT57), .ZN(new_n895));
  AND3_X1   g709(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n875), .B1(new_n873), .B2(new_n874), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n898), .B2(new_n669), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT117), .B1(new_n899), .B2(new_n883), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  INV_X1    g715(.A(new_n669), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n873), .A2(new_n874), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT54), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n876), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n905), .B2(new_n895), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n901), .B(new_n884), .C1(new_n906), .C2(new_n894), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n900), .A2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(new_n379), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n379), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n910), .A2(new_n911), .A3(new_n883), .ZN(G60));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n872), .B2(new_n876), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n884), .B1(new_n915), .B2(new_n601), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n598), .B2(new_n600), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n905), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n905), .A2(KEYINPUT118), .A3(new_n917), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT119), .Z(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT60), .Z(new_n925));
  AOI21_X1  g739(.A(KEYINPUT120), .B1(new_n903), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n927));
  INV_X1    g741(.A(new_n925), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n927), .B(new_n928), .C1(new_n873), .C2(new_n874), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n620), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n869), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT53), .B1(new_n931), .B2(new_n854), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n867), .A2(new_n825), .A3(new_n870), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n925), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n927), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n903), .A2(KEYINPUT120), .A3(new_n925), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n577), .A3(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n930), .A2(new_n937), .A3(new_n884), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n930), .A2(new_n937), .A3(KEYINPUT61), .A4(new_n884), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  OAI21_X1  g756(.A(G953), .B1(new_n391), .B2(new_n432), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n836), .A2(new_n842), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(G953), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n888), .B1(G898), .B2(new_n194), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  AOI21_X1  g761(.A(new_n194), .B1(G227), .B2(G900), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n950));
  INV_X1    g764(.A(new_n374), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n535), .B(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n655), .A2(new_n704), .A3(new_n634), .A4(new_n661), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT121), .ZN(new_n955));
  INV_X1    g769(.A(new_n767), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n711), .B1(new_n838), .B2(new_n831), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n663), .A2(new_n646), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n738), .ZN(new_n959));
  INV_X1    g773(.A(new_n756), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n956), .B(new_n961), .C1(KEYINPUT62), .C2(new_n953), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT122), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n953), .A2(KEYINPUT62), .ZN(new_n964));
  NOR4_X1   g778(.A1(new_n964), .A2(new_n767), .A3(new_n757), .A4(new_n958), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT121), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n954), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n952), .B1(new_n970), .B2(G953), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n949), .A2(KEYINPUT124), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n710), .A2(new_n697), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n859), .B1(new_n960), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n956), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n704), .A2(new_n634), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n661), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n757), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT123), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT123), .B1(new_n977), .B2(new_n757), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n194), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n952), .B1(G900), .B2(G953), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n972), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n950), .B1(new_n971), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(G953), .B1(new_n963), .B2(new_n969), .ZN(new_n988));
  INV_X1    g802(.A(new_n952), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n986), .B(new_n950), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n987), .A2(new_n991), .ZN(G72));
  OR2_X1    g806(.A1(new_n855), .A2(new_n871), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n537), .A2(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  NAND3_X1  g810(.A1(new_n537), .A2(KEYINPUT127), .A3(new_n510), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n963), .A2(new_n969), .A3(new_n944), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n996), .B(KEYINPUT125), .Z(new_n1001));
  AOI21_X1  g815(.A(new_n649), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1001), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n983), .B2(new_n944), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n513), .A2(new_n526), .A3(new_n501), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1003), .B(new_n884), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n981), .A2(new_n982), .ZN(new_n1008));
  INV_X1    g822(.A(new_n975), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1008), .A2(new_n944), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1006), .B1(new_n1010), .B2(new_n1001), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT126), .B1(new_n1011), .B2(new_n883), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n999), .B(new_n1002), .C1(new_n1007), .C2(new_n1012), .ZN(G57));
endmodule


