

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604;

  AND2_X1 U326 ( .A1(n582), .A2(n436), .ZN(n437) );
  INV_X1 U327 ( .A(KEYINPUT103), .ZN(n474) );
  XNOR2_X1 U328 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U329 ( .A(n477), .B(n476), .ZN(n484) );
  INV_X1 U330 ( .A(n451), .ZN(n452) );
  INV_X1 U331 ( .A(KEYINPUT70), .ZN(n327) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U333 ( .A(n328), .B(n327), .ZN(n329) );
  INV_X1 U334 ( .A(KEYINPUT64), .ZN(n333) );
  XNOR2_X1 U335 ( .A(n455), .B(n454), .ZN(n459) );
  XNOR2_X1 U336 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U337 ( .A(n333), .B(KEYINPUT41), .ZN(n334) );
  NOR2_X1 U338 ( .A1(n500), .A2(n530), .ZN(n491) );
  INV_X1 U339 ( .A(KEYINPUT58), .ZN(n464) );
  XNOR2_X1 U340 ( .A(n591), .B(n334), .ZN(n572) );
  XOR2_X1 U341 ( .A(n462), .B(n461), .Z(n571) );
  XNOR2_X1 U342 ( .A(n464), .B(G190GAT), .ZN(n465) );
  XNOR2_X1 U343 ( .A(n492), .B(G43GAT), .ZN(n493) );
  XNOR2_X1 U344 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(G183GAT), .B(KEYINPUT85), .Z(n295) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(KEYINPUT86), .ZN(n294) );
  XNOR2_X1 U348 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U349 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n297) );
  XNOR2_X1 U350 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n296) );
  XNOR2_X1 U351 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U352 ( .A(n299), .B(n298), .Z(n460) );
  XOR2_X1 U353 ( .A(G92GAT), .B(G64GAT), .Z(n326) );
  XOR2_X1 U354 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n301) );
  XNOR2_X1 U355 ( .A(G197GAT), .B(G211GAT), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n303) );
  XOR2_X1 U357 ( .A(G218GAT), .B(KEYINPUT21), .Z(n302) );
  XOR2_X1 U358 ( .A(n303), .B(n302), .Z(n412) );
  INV_X1 U359 ( .A(n412), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n326), .B(n304), .ZN(n306) );
  XNOR2_X1 U361 ( .A(G36GAT), .B(G176GAT), .ZN(n305) );
  XNOR2_X1 U362 ( .A(n306), .B(n305), .ZN(n311) );
  XOR2_X1 U363 ( .A(KEYINPUT97), .B(G204GAT), .Z(n308) );
  NAND2_X1 U364 ( .A1(G226GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U366 ( .A(G8GAT), .B(n309), .Z(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U368 ( .A(n460), .B(n312), .Z(n533) );
  INV_X1 U369 ( .A(n533), .ZN(n513) );
  XOR2_X1 U370 ( .A(G176GAT), .B(G120GAT), .Z(n446) );
  XOR2_X1 U371 ( .A(G99GAT), .B(G85GAT), .Z(n354) );
  XNOR2_X1 U372 ( .A(n446), .B(n354), .ZN(n332) );
  INV_X1 U373 ( .A(G204GAT), .ZN(n313) );
  NAND2_X1 U374 ( .A1(G148GAT), .A2(n313), .ZN(n316) );
  INV_X1 U375 ( .A(G148GAT), .ZN(n314) );
  NAND2_X1 U376 ( .A1(n314), .A2(G204GAT), .ZN(n315) );
  NAND2_X1 U377 ( .A1(n316), .A2(n315), .ZN(n318) );
  XNOR2_X1 U378 ( .A(G106GAT), .B(KEYINPUT69), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n406) );
  XNOR2_X1 U380 ( .A(G71GAT), .B(G57GAT), .ZN(n319) );
  XNOR2_X1 U381 ( .A(n319), .B(KEYINPUT13), .ZN(n385) );
  XNOR2_X1 U382 ( .A(n406), .B(n385), .ZN(n325) );
  XNOR2_X1 U383 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n321) );
  AND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n323) );
  INV_X1 U386 ( .A(KEYINPUT32), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n330) );
  XNOR2_X1 U389 ( .A(G78GAT), .B(n326), .ZN(n328) );
  XOR2_X1 U390 ( .A(n332), .B(n331), .Z(n591) );
  XOR2_X1 U391 ( .A(G197GAT), .B(G113GAT), .Z(n336) );
  XNOR2_X1 U392 ( .A(G169GAT), .B(G15GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n351) );
  XOR2_X1 U394 ( .A(G8GAT), .B(G1GAT), .Z(n373) );
  XOR2_X1 U395 ( .A(n373), .B(G43GAT), .Z(n340) );
  XOR2_X1 U396 ( .A(G29GAT), .B(G36GAT), .Z(n338) );
  XNOR2_X1 U397 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n367) );
  XNOR2_X1 U399 ( .A(n367), .B(G50GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U401 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n342) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U404 ( .A(n344), .B(n343), .Z(n349) );
  XOR2_X1 U405 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n346) );
  XNOR2_X1 U406 ( .A(G22GAT), .B(G141GAT), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n347), .B(KEYINPUT66), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U410 ( .A(n351), .B(n350), .Z(n517) );
  INV_X1 U411 ( .A(n517), .ZN(n586) );
  OR2_X1 U412 ( .A1(n572), .A2(n586), .ZN(n353) );
  XOR2_X1 U413 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n352) );
  XNOR2_X1 U414 ( .A(n353), .B(n352), .ZN(n370) );
  XOR2_X1 U415 ( .A(G50GAT), .B(G162GAT), .Z(n400) );
  XOR2_X1 U416 ( .A(n354), .B(n400), .Z(n356) );
  NAND2_X1 U417 ( .A1(G232GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U419 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n358) );
  XNOR2_X1 U420 ( .A(G190GAT), .B(KEYINPUT9), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U422 ( .A(n360), .B(n359), .Z(n365) );
  XOR2_X1 U423 ( .A(G43GAT), .B(G134GAT), .Z(n450) );
  XOR2_X1 U424 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n362) );
  XNOR2_X1 U425 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n450), .B(n363), .ZN(n364) );
  XNOR2_X1 U428 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U429 ( .A(n366), .B(G92GAT), .Z(n369) );
  XNOR2_X1 U430 ( .A(n367), .B(G106GAT), .ZN(n368) );
  XOR2_X1 U431 ( .A(n369), .B(n368), .Z(n566) );
  INV_X1 U432 ( .A(n566), .ZN(n495) );
  NOR2_X1 U433 ( .A1(n370), .A2(n495), .ZN(n388) );
  XOR2_X1 U434 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n372) );
  XNOR2_X1 U435 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U437 ( .A(G15GAT), .B(G127GAT), .Z(n449) );
  XOR2_X1 U438 ( .A(G211GAT), .B(n449), .Z(n375) );
  XNOR2_X1 U439 ( .A(n373), .B(G183GAT), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U441 ( .A(n377), .B(n376), .Z(n379) );
  NAND2_X1 U442 ( .A1(G231GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U444 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n381) );
  XNOR2_X1 U445 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n380) );
  XNOR2_X1 U446 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U447 ( .A(n383), .B(n382), .Z(n387) );
  XNOR2_X1 U448 ( .A(G22GAT), .B(G155GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n384), .B(G78GAT), .ZN(n407) );
  XNOR2_X1 U450 ( .A(n407), .B(n385), .ZN(n386) );
  XOR2_X1 U451 ( .A(n387), .B(n386), .Z(n596) );
  XOR2_X1 U452 ( .A(n596), .B(KEYINPUT113), .Z(n579) );
  NAND2_X1 U453 ( .A1(n388), .A2(n579), .ZN(n389) );
  XNOR2_X1 U454 ( .A(n389), .B(KEYINPUT47), .ZN(n396) );
  XOR2_X1 U455 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n392) );
  INV_X1 U456 ( .A(n596), .ZN(n390) );
  XOR2_X1 U457 ( .A(KEYINPUT36), .B(n566), .Z(n600) );
  NAND2_X1 U458 ( .A1(n390), .A2(n600), .ZN(n391) );
  XNOR2_X1 U459 ( .A(n392), .B(n391), .ZN(n394) );
  NAND2_X1 U460 ( .A1(n586), .A2(n591), .ZN(n393) );
  NOR2_X1 U461 ( .A1(n394), .A2(n393), .ZN(n395) );
  NOR2_X1 U462 ( .A1(n396), .A2(n395), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n397), .B(KEYINPUT48), .ZN(n543) );
  NOR2_X1 U464 ( .A1(n513), .A2(n543), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n398), .B(KEYINPUT54), .ZN(n582) );
  XOR2_X1 U466 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n402) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n399), .B(KEYINPUT2), .ZN(n426) );
  XNOR2_X1 U469 ( .A(n400), .B(n426), .ZN(n401) );
  XNOR2_X1 U470 ( .A(n402), .B(n401), .ZN(n411) );
  XOR2_X1 U471 ( .A(KEYINPUT90), .B(KEYINPUT93), .Z(n404) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U474 ( .A(n405), .B(KEYINPUT22), .Z(n409) );
  XNOR2_X1 U475 ( .A(n406), .B(n407), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U478 ( .A(n413), .B(n412), .Z(n478) );
  XOR2_X1 U479 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n415) );
  XNOR2_X1 U480 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n451) );
  XOR2_X1 U482 ( .A(n451), .B(KEYINPUT95), .Z(n417) );
  NAND2_X1 U483 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U485 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n419) );
  XNOR2_X1 U486 ( .A(G1GAT), .B(G57GAT), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U489 ( .A(G155GAT), .B(G148GAT), .Z(n423) );
  XNOR2_X1 U490 ( .A(G127GAT), .B(G120GAT), .ZN(n422) );
  XNOR2_X1 U491 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n430) );
  XOR2_X1 U493 ( .A(G85GAT), .B(n426), .Z(n428) );
  XNOR2_X1 U494 ( .A(G29GAT), .B(G162GAT), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U496 ( .A(n430), .B(n429), .Z(n435) );
  XOR2_X1 U497 ( .A(KEYINPUT96), .B(KEYINPUT4), .Z(n432) );
  XNOR2_X1 U498 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n431) );
  XNOR2_X1 U499 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U500 ( .A(G134GAT), .B(n433), .ZN(n434) );
  XOR2_X1 U501 ( .A(n435), .B(n434), .Z(n531) );
  NOR2_X1 U502 ( .A1(n478), .A2(n531), .ZN(n436) );
  XNOR2_X1 U503 ( .A(KEYINPUT120), .B(n437), .ZN(n439) );
  INV_X1 U504 ( .A(n439), .ZN(n438) );
  NAND2_X1 U505 ( .A1(n438), .A2(KEYINPUT55), .ZN(n442) );
  INV_X1 U506 ( .A(KEYINPUT55), .ZN(n440) );
  NAND2_X1 U507 ( .A1(n440), .A2(n439), .ZN(n441) );
  NAND2_X1 U508 ( .A1(n442), .A2(n441), .ZN(n574) );
  XOR2_X1 U509 ( .A(KEYINPUT83), .B(G71GAT), .Z(n444) );
  XNOR2_X1 U510 ( .A(KEYINPUT88), .B(KEYINPUT82), .ZN(n443) );
  XNOR2_X1 U511 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U512 ( .A(n445), .B(KEYINPUT84), .Z(n448) );
  XNOR2_X1 U513 ( .A(n446), .B(G99GAT), .ZN(n447) );
  XNOR2_X1 U514 ( .A(n448), .B(n447), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n450), .B(n449), .ZN(n453) );
  XOR2_X1 U516 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n457) );
  NAND2_X1 U517 ( .A1(G227GAT), .A2(G233GAT), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n457), .B(n456), .ZN(n458) );
  XOR2_X1 U519 ( .A(n459), .B(n458), .Z(n462) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT81), .ZN(n461) );
  INV_X1 U521 ( .A(n571), .ZN(n568) );
  AND2_X1 U522 ( .A1(n568), .A2(n495), .ZN(n463) );
  AND2_X1 U523 ( .A1(n574), .A2(n463), .ZN(n466) );
  AND2_X1 U524 ( .A1(n517), .A2(n591), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n467), .B(KEYINPUT71), .ZN(n500) );
  XOR2_X1 U526 ( .A(KEYINPUT37), .B(KEYINPUT106), .Z(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT107), .B(n468), .ZN(n490) );
  INV_X1 U528 ( .A(n531), .ZN(n581) );
  XOR2_X1 U529 ( .A(n533), .B(KEYINPUT27), .Z(n482) );
  NOR2_X1 U530 ( .A1(n581), .A2(n482), .ZN(n541) );
  XNOR2_X1 U531 ( .A(KEYINPUT28), .B(n478), .ZN(n536) );
  INV_X1 U532 ( .A(n536), .ZN(n545) );
  NAND2_X1 U533 ( .A1(n541), .A2(n545), .ZN(n469) );
  XNOR2_X1 U534 ( .A(KEYINPUT98), .B(n469), .ZN(n471) );
  XOR2_X1 U535 ( .A(KEYINPUT89), .B(n568), .Z(n470) );
  NOR2_X1 U536 ( .A1(n471), .A2(n470), .ZN(n487) );
  NOR2_X1 U537 ( .A1(n513), .A2(n571), .ZN(n472) );
  XOR2_X1 U538 ( .A(KEYINPUT101), .B(n472), .Z(n473) );
  NOR2_X1 U539 ( .A1(n478), .A2(n473), .ZN(n477) );
  XOR2_X1 U540 ( .A(KEYINPUT25), .B(KEYINPUT102), .Z(n475) );
  XOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT26), .Z(n480) );
  NAND2_X1 U542 ( .A1(n478), .A2(n571), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U544 ( .A(KEYINPUT99), .B(n481), .ZN(n583) );
  NOR2_X1 U545 ( .A1(n482), .A2(n583), .ZN(n483) );
  NOR2_X1 U546 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U547 ( .A1(n531), .A2(n485), .ZN(n486) );
  NOR2_X1 U548 ( .A1(n487), .A2(n486), .ZN(n498) );
  NAND2_X1 U549 ( .A1(n596), .A2(n600), .ZN(n488) );
  NOR2_X1 U550 ( .A1(n498), .A2(n488), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n530) );
  XOR2_X1 U552 ( .A(KEYINPUT38), .B(n491), .Z(n515) );
  NOR2_X1 U553 ( .A1(n515), .A2(n571), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n492) );
  NOR2_X1 U555 ( .A1(n495), .A2(n596), .ZN(n496) );
  XOR2_X1 U556 ( .A(KEYINPUT16), .B(n496), .Z(n497) );
  NOR2_X1 U557 ( .A1(n498), .A2(n497), .ZN(n518) );
  INV_X1 U558 ( .A(n518), .ZN(n499) );
  NOR2_X1 U559 ( .A1(n500), .A2(n499), .ZN(n508) );
  NAND2_X1 U560 ( .A1(n531), .A2(n508), .ZN(n504) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n502) );
  XNOR2_X1 U562 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1324GAT) );
  NAND2_X1 U565 ( .A1(n533), .A2(n508), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U567 ( .A(G15GAT), .B(KEYINPUT35), .Z(n507) );
  NAND2_X1 U568 ( .A1(n508), .A2(n568), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1326GAT) );
  NAND2_X1 U570 ( .A1(n508), .A2(n536), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U572 ( .A(G29GAT), .B(KEYINPUT108), .ZN(n512) );
  NOR2_X1 U573 ( .A1(n515), .A2(n581), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n510), .B(KEYINPUT39), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1328GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n515), .ZN(n514) );
  XOR2_X1 U577 ( .A(G36GAT), .B(n514), .Z(G1329GAT) );
  NOR2_X1 U578 ( .A1(n515), .A2(n545), .ZN(n516) );
  XOR2_X1 U579 ( .A(G50GAT), .B(n516), .Z(G1331GAT) );
  NOR2_X1 U580 ( .A1(n517), .A2(n572), .ZN(n528) );
  NAND2_X1 U581 ( .A1(n528), .A2(n518), .ZN(n519) );
  XOR2_X1 U582 ( .A(KEYINPUT110), .B(n519), .Z(n525) );
  NAND2_X1 U583 ( .A1(n525), .A2(n531), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT42), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G57GAT), .B(n521), .ZN(G1332GAT) );
  XOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT111), .Z(n523) );
  NAND2_X1 U587 ( .A1(n525), .A2(n533), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n568), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U592 ( .A1(n536), .A2(n525), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1335GAT) );
  INV_X1 U594 ( .A(n528), .ZN(n529) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n537) );
  NAND2_X1 U596 ( .A1(n537), .A2(n531), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G85GAT), .B(n532), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n537), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n537), .A2(n568), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(G106GAT), .B(n540), .Z(G1339GAT) );
  INV_X1 U606 ( .A(n541), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(KEYINPUT115), .B(n544), .ZN(n557) );
  NOR2_X1 U609 ( .A1(n571), .A2(n557), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n586), .A2(n553), .ZN(n547) );
  XOR2_X1 U612 ( .A(G113GAT), .B(n547), .Z(G1340GAT) );
  NOR2_X1 U613 ( .A1(n572), .A2(n553), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  NOR2_X1 U616 ( .A1(n579), .A2(n553), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(G127GAT), .B(n552), .Z(G1342GAT) );
  NOR2_X1 U620 ( .A1(n566), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(G134GAT), .B(n556), .Z(G1343GAT) );
  OR2_X1 U624 ( .A1(n583), .A2(n557), .ZN(n565) );
  NOR2_X1 U625 ( .A1(n586), .A2(n565), .ZN(n558) );
  XOR2_X1 U626 ( .A(n558), .B(KEYINPUT118), .Z(n559) );
  XNOR2_X1 U627 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  NOR2_X1 U628 ( .A1(n572), .A2(n565), .ZN(n561) );
  XNOR2_X1 U629 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U631 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U632 ( .A1(n596), .A2(n565), .ZN(n564) );
  XNOR2_X1 U633 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n563) );
  XNOR2_X1 U634 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NOR2_X1 U635 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U636 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NAND2_X1 U637 ( .A1(n574), .A2(n568), .ZN(n578) );
  NOR2_X1 U638 ( .A1(n586), .A2(n578), .ZN(n570) );
  XNOR2_X1 U639 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n569) );
  XNOR2_X1 U640 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  NOR2_X1 U641 ( .A1(n572), .A2(n571), .ZN(n573) );
  AND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U643 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n575) );
  XNOR2_X1 U644 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U647 ( .A(G183GAT), .B(n580), .Z(G1350GAT) );
  NAND2_X1 U648 ( .A1(n582), .A2(n581), .ZN(n584) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(KEYINPUT122), .B(n585), .ZN(n601) );
  INV_X1 U651 ( .A(n601), .ZN(n597) );
  NOR2_X1 U652 ( .A1(n586), .A2(n597), .ZN(n590) );
  XOR2_X1 U653 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n588) );
  XNOR2_X1 U654 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n590), .B(n589), .ZN(G1352GAT) );
  NOR2_X1 U657 ( .A1(n591), .A2(n597), .ZN(n595) );
  XOR2_X1 U658 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n593) );
  XNOR2_X1 U659 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n592) );
  XNOR2_X1 U660 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n595), .B(n594), .ZN(G1353GAT) );
  NOR2_X1 U662 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U663 ( .A(G211GAT), .B(n598), .Z(n599) );
  XNOR2_X1 U664 ( .A(KEYINPUT126), .B(n599), .ZN(G1354GAT) );
  XOR2_X1 U665 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n603) );
  NAND2_X1 U666 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U667 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U668 ( .A(G218GAT), .B(n604), .ZN(G1355GAT) );
endmodule

