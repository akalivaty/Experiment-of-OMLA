//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT67), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n476), .B2(new_n462), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n464), .A2(new_n466), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OAI21_X1  g063(.A(G2104), .B1(new_n462), .B2(G114), .ZN(new_n489));
  NOR2_X1   g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT68), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n492), .A2(new_n494), .A3(new_n495), .A4(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(KEYINPUT69), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n499), .A2(new_n464), .A3(new_n466), .A4(new_n462), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n475), .A2(G126), .A3(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n475), .A2(KEYINPUT4), .A3(new_n462), .A4(new_n499), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n497), .A2(new_n502), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G88), .B1(G62), .B2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n515), .A2(new_n521), .ZN(G166));
  AOI22_X1  g097(.A1(new_n512), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(new_n520), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n514), .B1(new_n510), .B2(new_n511), .ZN(new_n525));
  NAND2_X1  g100(.A1(KEYINPUT71), .A2(G51), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT71), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n524), .A2(new_n528), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI21_X1  g107(.A(new_n520), .B1(new_n510), .B2(new_n511), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n520), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n525), .A2(G52), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n520), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT72), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n533), .A2(G81), .B1(new_n525), .B2(G43), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n548), .A3(G651), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n512), .A2(G53), .A3(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n520), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n533), .A2(G91), .B1(new_n562), .B2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G166), .ZN(G303));
  AND2_X1   g140(.A1(new_n517), .A2(new_n519), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n512), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G87), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n567), .A2(KEYINPUT73), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G74), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n509), .B1(new_n520), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n571), .B1(G49), .B2(new_n525), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT73), .B1(new_n567), .B2(new_n568), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n520), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n533), .A2(G86), .B1(G48), .B2(new_n525), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n577), .A2(new_n581), .A3(G651), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n533), .A2(G85), .ZN(new_n584));
  XOR2_X1   g159(.A(KEYINPUT75), .B(G47), .Z(new_n585));
  NAND2_X1  g160(.A1(new_n525), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n566), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n584), .B(new_n586), .C1(new_n509), .C2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OR3_X1    g165(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n520), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n525), .B2(G54), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT10), .B1(new_n567), .B2(new_n590), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT76), .Z(new_n598));
  OAI21_X1  g173(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n589), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  XNOR2_X1  g176(.A(G299), .B(KEYINPUT77), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  NOR2_X1   g181(.A1(new_n551), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n605), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT78), .Z(G323));
  XOR2_X1   g185(.A(G323), .B(KEYINPUT79), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n483), .A2(G135), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  INV_X1    g189(.A(G111), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G2105), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT82), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n613), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(KEYINPUT81), .B1(new_n481), .B2(G123), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n481), .A2(G123), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g197(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2096), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G2100), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n627), .B(new_n629), .Z(new_n630));
  OAI211_X1 g205(.A(new_n624), .B(new_n630), .C1(new_n628), .C2(G2100), .ZN(G156));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2430), .Z(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n641), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n645), .B1(new_n642), .B2(new_n646), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n633), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n651), .A2(new_n647), .A3(new_n632), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n652), .A3(G14), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT85), .Z(G401));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n655), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2096), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n657), .A2(new_n658), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n659), .A3(KEYINPUT17), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(new_n660), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT19), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(KEYINPUT89), .ZN(new_n680));
  INV_X1    g255(.A(new_n678), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n669), .A2(new_n670), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n674), .ZN(new_n685));
  INV_X1    g260(.A(new_n683), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(new_n686), .A3(new_n671), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n679), .A2(new_n682), .A3(new_n684), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT90), .B(G1986), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n692), .ZN(new_n695));
  AND3_X1   g270(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(G229));
  NOR2_X1   g273(.A1(G16), .A2(G23), .ZN(new_n699));
  INV_X1    g274(.A(G288), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G6), .B(G305), .S(G16), .Z(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n703), .A2(new_n706), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT34), .Z(new_n712));
  MUX2_X1   g287(.A(G24), .B(G290), .S(G16), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  INV_X1    g289(.A(G1986), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT35), .B(G1991), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n481), .A2(G119), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n483), .A2(G131), .ZN(new_n722));
  OR2_X1    g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  AOI211_X1 g302(.A(new_n716), .B(new_n717), .C1(new_n718), .C2(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n712), .B(new_n728), .C1(new_n718), .C2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n729), .B(new_n730), .Z(new_n731));
  AND2_X1   g306(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n719), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n719), .ZN(new_n735));
  MUX2_X1   g310(.A(new_n734), .B(new_n735), .S(KEYINPUT99), .Z(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G2078), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT97), .B1(G5), .B2(G16), .ZN(new_n738));
  OR3_X1    g313(.A1(KEYINPUT97), .A2(G5), .A3(G16), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n738), .B(new_n739), .C1(G301), .C2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n740), .A2(G21), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G286), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1966), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n623), .A2(G29), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT31), .B(G11), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT96), .ZN(new_n750));
  INV_X1    g325(.A(G28), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT30), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n750), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n741), .A2(new_n742), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(KEYINPUT98), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n744), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT24), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(G34), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(G34), .ZN(new_n764));
  AOI21_X1  g339(.A(G29), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n478), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n719), .A2(G33), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT25), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n483), .A2(G139), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n771), .B(new_n772), .C1(new_n462), .C2(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT94), .Z(new_n775));
  OAI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(new_n719), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G2072), .Z(new_n777));
  NOR2_X1   g352(.A1(G29), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n483), .A2(G141), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n481), .A2(G129), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n781));
  NAND3_X1  g356(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT26), .Z(new_n783));
  NAND4_X1  g358(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n778), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT27), .B(G1996), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G2078), .B2(new_n736), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n761), .A2(new_n768), .A3(new_n777), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n598), .A2(new_n740), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G4), .B2(new_n740), .ZN(new_n792));
  INV_X1    g367(.A(G1348), .ZN(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n719), .A2(G26), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n481), .A2(G128), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT93), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n483), .A2(G140), .ZN(new_n798));
  NOR2_X1   g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n795), .B1(new_n803), .B2(G29), .ZN(new_n804));
  MUX2_X1   g379(.A(new_n795), .B(new_n804), .S(KEYINPUT28), .Z(new_n805));
  OAI22_X1  g380(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n790), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n794), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n792), .A2(new_n793), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n766), .A2(new_n767), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT95), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n719), .A2(G35), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G162), .B2(new_n719), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT100), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT29), .ZN(new_n815));
  INV_X1    g390(.A(G2090), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n740), .A2(G19), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n551), .B2(new_n740), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(G1341), .Z(new_n820));
  NAND2_X1  g395(.A1(G299), .A2(G16), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n740), .A2(KEYINPUT23), .A3(G20), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT23), .ZN(new_n823));
  INV_X1    g398(.A(G20), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(G16), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n827));
  INV_X1    g402(.A(G1956), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n826), .B(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n815), .B2(new_n816), .ZN(new_n831));
  AND4_X1   g406(.A1(new_n811), .A2(new_n817), .A3(new_n820), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT103), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n809), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n817), .A2(new_n831), .A3(new_n811), .A4(new_n820), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n790), .A2(new_n836), .A3(new_n837), .A4(new_n806), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n838), .A2(KEYINPUT103), .A3(new_n808), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n733), .B1(new_n835), .B2(new_n839), .ZN(G311));
  NOR2_X1   g415(.A1(new_n833), .A2(new_n834), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT103), .B1(new_n838), .B2(new_n808), .ZN(new_n842));
  OAI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(new_n732), .B2(new_n731), .ZN(G150));
  NAND2_X1  g418(.A1(new_n598), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT39), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n550), .A2(KEYINPUT104), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n550), .A2(KEYINPUT104), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n566), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(new_n509), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G55), .B2(new_n525), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n533), .A2(G93), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n847), .A3(new_n848), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n846), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT105), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n854), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(G145));
  XOR2_X1   g440(.A(new_n505), .B(KEYINPUT106), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n623), .B(new_n487), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(new_n478), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n623), .B(G162), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(G160), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n478), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(G160), .ZN(new_n873));
  INV_X1    g448(.A(new_n866), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n483), .A2(G142), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n880), .B(new_n881), .C1(G118), .C2(new_n462), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n481), .A2(G130), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n877), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n802), .A2(new_n725), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n726), .B1(new_n797), .B2(new_n801), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n784), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n784), .B1(new_n885), .B2(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n785), .ZN(new_n892));
  INV_X1    g467(.A(new_n884), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n887), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n775), .B(new_n626), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n890), .B2(new_n894), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n876), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G37), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n890), .A2(new_n894), .ZN(new_n901));
  INV_X1    g476(.A(new_n895), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n871), .A2(new_n875), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n904), .A3(new_n896), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n899), .A2(new_n900), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g482(.A1(new_n854), .A2(G868), .ZN(new_n908));
  XNOR2_X1  g483(.A(G288), .B(G166), .ZN(new_n909));
  XNOR2_X1  g484(.A(G305), .B(G290), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT42), .Z(new_n912));
  XNOR2_X1  g487(.A(new_n858), .B(new_n608), .ZN(new_n913));
  XOR2_X1   g488(.A(G299), .B(new_n597), .Z(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT41), .ZN(new_n915));
  XNOR2_X1  g490(.A(G299), .B(new_n597), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n920), .B1(new_n914), .B2(new_n913), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n912), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  MUX2_X1   g499(.A(new_n923), .B(new_n912), .S(new_n924), .Z(new_n925));
  AOI21_X1  g500(.A(new_n908), .B1(new_n925), .B2(G868), .ZN(G295));
  AOI21_X1  g501(.A(new_n908), .B1(new_n925), .B2(G868), .ZN(G331));
  INV_X1    g502(.A(new_n911), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n524), .A2(new_n528), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n929), .A2(G171), .A3(new_n930), .A4(new_n530), .ZN(new_n931));
  NAND2_X1  g506(.A1(G171), .A2(new_n930), .ZN(new_n932));
  NAND2_X1  g507(.A1(G301), .A2(KEYINPUT109), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(G286), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n857), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n856), .B1(new_n848), .B2(new_n847), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n931), .A2(new_n934), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n855), .A3(new_n857), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n938), .A2(new_n916), .A3(new_n940), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n938), .A2(new_n940), .B1(new_n918), .B2(new_n915), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n928), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n919), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n916), .A3(new_n940), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n911), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n943), .A2(new_n947), .A3(new_n900), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT43), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n943), .A2(new_n947), .A3(new_n950), .A4(new_n900), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT44), .Z(G397));
  XNOR2_X1  g528(.A(new_n802), .B(G2067), .ZN(new_n954));
  INV_X1    g529(.A(G1996), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n784), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n725), .A2(new_n718), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  OAI22_X1  g534(.A1(new_n957), .A2(new_n959), .B1(G2067), .B2(new_n803), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n505), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n473), .A2(G40), .A3(new_n477), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n967), .B(KEYINPUT122), .Z(new_n968));
  INV_X1    g543(.A(new_n966), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n954), .B2(new_n785), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(KEYINPUT123), .B2(KEYINPUT46), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n966), .A2(new_n955), .ZN(new_n972));
  NOR2_X1   g547(.A1(KEYINPUT123), .A2(KEYINPUT46), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n972), .B(new_n973), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n725), .A2(new_n718), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n957), .A2(new_n978), .A3(new_n958), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n966), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n966), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT125), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n968), .B(new_n977), .C1(new_n981), .C2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n505), .B2(new_n961), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n965), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n505), .A2(new_n987), .A3(new_n961), .ZN(new_n990));
  AOI21_X1  g565(.A(G1956), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n473), .A2(G40), .A3(new_n477), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT56), .B(G2072), .ZN(new_n994));
  AND4_X1   g569(.A1(new_n964), .A2(new_n992), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n991), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT57), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT9), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n558), .B(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n563), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n559), .A2(KEYINPUT57), .A3(new_n563), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n505), .A2(new_n987), .A3(new_n961), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1005), .A2(new_n988), .A3(new_n965), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n965), .A2(new_n962), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI22_X1  g583(.A1(new_n1006), .A2(G1348), .B1(new_n1008), .B2(G2067), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1009), .A2(new_n598), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n996), .A2(new_n1003), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1004), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n964), .A2(new_n992), .A3(new_n955), .A4(new_n993), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT58), .B(G1341), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n505), .B2(new_n961), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(new_n965), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(KEYINPUT113), .A3(new_n955), .A4(new_n993), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n551), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1021), .A2(KEYINPUT59), .A3(new_n551), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1003), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT114), .B(new_n1026), .C1(new_n991), .C2(new_n995), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT61), .ZN(new_n1028));
  INV_X1    g603(.A(new_n988), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(new_n992), .A3(new_n990), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n828), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1019), .A2(new_n993), .A3(new_n994), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(KEYINPUT114), .A4(new_n1003), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1027), .A2(new_n1028), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1028), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1024), .B(new_n1025), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT60), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1009), .A2(new_n1037), .ZN(new_n1038));
  OAI221_X1 g613(.A(KEYINPUT60), .B1(new_n1008), .B2(G2067), .C1(new_n1006), .C2(G1348), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n598), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n598), .B2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1012), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT115), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1019), .A2(new_n993), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(G2078), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1030), .A2(new_n742), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1018), .A2(new_n469), .A3(new_n472), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1044), .A2(G2078), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(G40), .A3(new_n993), .A4(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G171), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n505), .A2(new_n1053), .A3(KEYINPUT45), .A4(new_n961), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n993), .A2(KEYINPUT112), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1019), .A2(new_n1054), .A3(new_n1055), .A4(new_n1049), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1046), .A2(G301), .A3(new_n1047), .A4(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(KEYINPUT54), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n515), .B2(new_n521), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT55), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1045), .A2(new_n709), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1006), .A2(new_n816), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1059), .B(new_n1061), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(G8), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1981), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n579), .A2(new_n580), .A3(new_n1069), .A4(new_n582), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1070), .A2(KEYINPUT111), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1070), .B2(KEYINPUT111), .ZN(new_n1073));
  OAI211_X1 g648(.A(G1981), .B(G305), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1073), .ZN(new_n1075));
  NAND2_X1  g650(.A1(G305), .A2(G1981), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1070), .A2(KEYINPUT111), .A3(new_n1071), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1007), .A2(new_n1059), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1074), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n569), .A2(G1976), .A3(new_n572), .A4(new_n573), .ZN(new_n1081));
  XOR2_X1   g656(.A(new_n1081), .B(KEYINPUT110), .Z(new_n1082));
  INV_X1    g657(.A(G1976), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(G288), .B2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1079), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1079), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1081), .B(KEYINPUT110), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT52), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1080), .A2(new_n1085), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1058), .A2(new_n1068), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  INV_X1    g667(.A(G1966), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1055), .A2(new_n964), .A3(new_n992), .A4(new_n1054), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1093), .A2(new_n1094), .B1(new_n1006), .B2(new_n767), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n1095), .B2(new_n1059), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1006), .A2(new_n767), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT116), .A3(G8), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G286), .A2(G8), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1096), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT51), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1104), .B(new_n1101), .C1(new_n1095), .C2(new_n1059), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1099), .A2(G8), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1104), .A4(new_n1101), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1103), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1095), .A2(new_n1101), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1091), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1115));
  AOI21_X1  g690(.A(G301), .B1(new_n1115), .B2(new_n1056), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1051), .A2(G171), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(KEYINPUT119), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT115), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1123), .B(new_n1012), .C1(new_n1036), .C2(new_n1041), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1043), .A2(new_n1113), .A3(new_n1122), .A4(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1090), .A2(new_n1064), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1080), .A2(new_n1083), .A3(new_n700), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1086), .B1(new_n1127), .B2(new_n1070), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1059), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1068), .A2(new_n1090), .A3(G168), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1089), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1133), .A2(KEYINPUT63), .A3(G168), .A4(new_n1129), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n1126), .B(new_n1128), .C1(new_n1132), .C2(new_n1134), .ZN(new_n1135));
  AND3_X1   g710(.A1(new_n1125), .A2(KEYINPUT120), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1111), .B1(new_n1138), .B2(new_n1103), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1133), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1129), .A2(KEYINPUT116), .B1(G8), .B2(G286), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1104), .B1(new_n1143), .B2(new_n1096), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1112), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1116), .B1(new_n1145), .B2(KEYINPUT62), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1137), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1133), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1145), .B2(KEYINPUT62), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT121), .A4(new_n1116), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT120), .B1(new_n1125), .B2(new_n1135), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1136), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n980), .B1(G1986), .B2(G290), .ZN(new_n1155));
  INV_X1    g730(.A(new_n982), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n969), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n986), .B1(new_n1154), .B2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1160));
  AOI211_X1 g734(.A(G227), .B(G229), .C1(new_n949), .C2(new_n951), .ZN(new_n1161));
  AND3_X1   g735(.A1(new_n906), .A2(G319), .A3(new_n653), .ZN(new_n1162));
  AOI21_X1  g736(.A(KEYINPUT126), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g737(.A(G227), .B1(new_n949), .B2(new_n951), .ZN(new_n1164));
  INV_X1    g738(.A(G229), .ZN(new_n1165));
  AND4_X1   g739(.A1(KEYINPUT126), .A2(new_n1164), .A3(new_n1165), .A4(new_n1162), .ZN(new_n1166));
  OAI21_X1  g740(.A(new_n1160), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g744(.A1(new_n1161), .A2(KEYINPUT126), .A3(new_n1162), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n1171), .A3(KEYINPUT127), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n1167), .A2(new_n1172), .ZN(G308));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1171), .ZN(G225));
endmodule


