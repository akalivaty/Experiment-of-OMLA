//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT82), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G116), .ZN(new_n192));
  INV_X1    g006(.A(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT5), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(G113), .B1(new_n192), .B2(KEYINPUT5), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G107), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n202), .A2(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(G101), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  INV_X1    g024(.A(G101), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .A4(new_n203), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  OR2_X1    g027(.A1(new_n201), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(new_n210), .A3(new_n203), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G101), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT4), .A3(new_n212), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n195), .B(new_n196), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n219), .A3(G101), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n190), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g036(.A1(new_n222), .A2(KEYINPUT6), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n214), .A2(new_n221), .A3(new_n189), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n214), .A2(new_n221), .A3(KEYINPUT83), .A4(new_n189), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n223), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G143), .ZN(new_n232));
  INV_X1    g046(.A(G143), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n233), .A2(KEYINPUT64), .A3(G146), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT64), .B1(new_n233), .B2(G146), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  OR2_X1    g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(new_n241), .A2(new_n237), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n239), .A2(G125), .A3(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n233), .A2(G146), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  OAI21_X1  g059(.A(G128), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT66), .B1(new_n236), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n231), .B2(G143), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n233), .A2(KEYINPUT64), .A3(G146), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n245), .A2(G128), .ZN(new_n256));
  OAI22_X1  g070(.A1(new_n247), .A2(new_n255), .B1(new_n241), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G125), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n243), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G224), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G953), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n259), .B(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(G902), .B1(new_n230), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT7), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n259), .A2(new_n264), .A3(new_n261), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n259), .B2(new_n261), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n189), .B(KEYINPUT8), .ZN(new_n267));
  INV_X1    g081(.A(new_n213), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n200), .B(KEYINPUT84), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n197), .B(new_n268), .C1(new_n269), .C2(new_n199), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n270), .B(KEYINPUT85), .Z(new_n271));
  AND2_X1   g085(.A1(new_n201), .A2(new_n213), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n267), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n226), .A2(new_n227), .B1(new_n264), .B2(new_n259), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n263), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n263), .A2(new_n277), .A3(new_n275), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n188), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G237), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n283), .A3(G214), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(G143), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT18), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT18), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n285), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  INV_X1    g104(.A(G140), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(G125), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n258), .A2(G140), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n294), .B(G146), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n288), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n285), .B(new_n286), .ZN(new_n297));
  INV_X1    g111(.A(new_n294), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT16), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT74), .B1(new_n292), .B2(KEYINPUT16), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT16), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n291), .A4(G125), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n299), .A2(G146), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n294), .A2(KEYINPUT86), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT19), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(G146), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n296), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G113), .B(G122), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(new_n202), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n287), .A2(KEYINPUT17), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n297), .B2(KEYINPUT17), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n300), .B(new_n303), .C1(new_n294), .C2(new_n302), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n318));
  OR3_X1    g132(.A1(new_n317), .A2(new_n318), .A3(new_n231), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n304), .A2(new_n318), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n317), .B2(new_n231), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n317), .A2(new_n321), .A3(new_n231), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n319), .B(new_n320), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n312), .B(new_n296), .C1(new_n316), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G475), .ZN(new_n327));
  INV_X1    g141(.A(G902), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT20), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n330), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT87), .B(G475), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n296), .B1(new_n316), .B2(new_n324), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(new_n312), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n335), .B2(G902), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G478), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT15), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G128), .A3(new_n233), .ZN(new_n342));
  XNOR2_X1  g156(.A(G128), .B(G143), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n342), .B(G134), .C1(new_n344), .C2(new_n341), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G134), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G116), .B(G122), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(new_n209), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n343), .B(G134), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n353), .A2(KEYINPUT90), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n209), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT91), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n193), .A2(KEYINPUT14), .A3(G122), .ZN(new_n357));
  INV_X1    g171(.A(new_n350), .ZN(new_n358));
  OAI211_X1 g172(.A(G107), .B(new_n357), .C1(new_n358), .C2(KEYINPUT14), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n353), .A2(KEYINPUT90), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n354), .A2(new_n356), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n352), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT9), .B(G234), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n364), .A2(new_n365), .A3(G953), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n352), .A2(new_n366), .A3(new_n361), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n340), .B1(new_n370), .B2(new_n328), .ZN(new_n371));
  AOI211_X1 g185(.A(G902), .B(new_n339), .C1(new_n368), .C2(new_n369), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n337), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n283), .A2(G952), .ZN(new_n376));
  NAND2_X1  g190(.A1(G234), .A2(G237), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  XOR2_X1   g193(.A(KEYINPUT21), .B(G898), .Z(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(G902), .A3(G953), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n281), .A2(new_n375), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G469), .ZN(new_n387));
  XOR2_X1   g201(.A(G110), .B(G140), .Z(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT80), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n283), .A2(G227), .ZN(new_n390));
  XOR2_X1   g204(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n241), .A2(new_n256), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n393), .B1(new_n241), .B2(new_n246), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n392), .B1(new_n394), .B2(new_n213), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n395), .B(KEYINPUT81), .Z(new_n396));
  AND2_X1   g210(.A1(new_n239), .A2(new_n242), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n220), .A3(new_n217), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n257), .A2(KEYINPUT10), .A3(new_n268), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n348), .A2(G137), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT11), .ZN(new_n402));
  INV_X1    g216(.A(G137), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(G134), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT11), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n348), .B2(G137), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G131), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n402), .A2(new_n405), .A3(new_n286), .A4(new_n407), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(KEYINPUT65), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT65), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n408), .A2(new_n412), .A3(G131), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n400), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n396), .A2(new_n414), .A3(new_n398), .A4(new_n399), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n391), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n236), .A2(KEYINPUT66), .A3(new_n246), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n252), .B1(new_n251), .B2(new_n254), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n393), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n213), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n213), .B2(new_n394), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n415), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(KEYINPUT12), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(KEYINPUT12), .ZN(new_n426));
  AND4_X1   g240(.A1(new_n417), .A2(new_n425), .A3(new_n391), .A4(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n387), .B(new_n328), .C1(new_n418), .C2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n387), .A2(new_n328), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n417), .A2(new_n425), .A3(new_n426), .ZN(new_n431));
  INV_X1    g245(.A(new_n391), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n416), .A2(new_n417), .A3(new_n391), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(G469), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n428), .A2(new_n430), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G221), .B1(new_n364), .B2(G902), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT79), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT92), .B1(new_n386), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n280), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n277), .B1(new_n263), .B2(new_n275), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n187), .B(new_n385), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n436), .A2(new_n438), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .A4(new_n375), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT67), .ZN(new_n448));
  OAI21_X1  g262(.A(G131), .B1(new_n404), .B2(new_n401), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n410), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n257), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT67), .B1(new_n421), .B2(new_n450), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n397), .A2(new_n413), .A3(new_n411), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT30), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n257), .A2(new_n451), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n454), .A3(KEYINPUT30), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n218), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n461));
  INV_X1    g275(.A(new_n218), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n454), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(G101), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n282), .A2(new_n283), .A3(G210), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n460), .A2(new_n461), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n461), .B1(new_n460), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT31), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n474));
  NAND2_X1  g288(.A1(new_n455), .A2(new_n218), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n475), .B2(new_n463), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n464), .A2(KEYINPUT28), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n469), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT31), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n460), .A2(new_n479), .A3(new_n470), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n460), .A2(KEYINPUT69), .A3(new_n479), .A4(new_n470), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n473), .A2(new_n478), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G472), .A2(G902), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT32), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(KEYINPUT32), .A3(new_n485), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n462), .B1(new_n458), .B2(new_n454), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n464), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(KEYINPUT28), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n477), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT29), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n469), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(G902), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n476), .A2(new_n469), .A3(new_n477), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n460), .A2(new_n463), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n497), .B(new_n494), .C1(new_n468), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G472), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n488), .A2(new_n489), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n191), .A2(G128), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n253), .A2(G119), .ZN(new_n504));
  OR3_X1    g318(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT72), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT72), .B1(new_n503), .B2(new_n504), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT24), .B(G110), .Z(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT73), .ZN(new_n510));
  INV_X1    g324(.A(new_n503), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT23), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n510), .B(new_n511), .C1(new_n504), .C2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n253), .B(G119), .C1(KEYINPUT73), .C2(KEYINPUT23), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G110), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n324), .A2(new_n509), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n518));
  OAI221_X1 g332(.A(new_n518), .B1(new_n515), .B2(G110), .C1(new_n507), .C2(new_n508), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n515), .A2(G110), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n508), .B1(new_n505), .B2(new_n506), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT77), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n298), .A2(new_n231), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n519), .A2(new_n522), .A3(new_n304), .A4(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT78), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n517), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT22), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(G137), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n525), .B1(new_n517), .B2(new_n524), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI211_X1 g347(.A(new_n525), .B(new_n530), .C1(new_n517), .C2(new_n524), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n328), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT25), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n537), .B(new_n328), .C1(new_n533), .C2(new_n534), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n365), .B1(G234), .B2(new_n328), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT71), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n539), .A2(G902), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n533), .B2(new_n534), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n440), .A2(new_n447), .A3(new_n502), .A4(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT93), .B(G101), .Z(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(G3));
  NAND2_X1  g362(.A1(KEYINPUT94), .A2(G472), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n484), .A2(new_n328), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n484), .B2(new_n328), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n550), .A2(new_n439), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n545), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n362), .A2(KEYINPUT95), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT33), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n370), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n370), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n556), .A2(G478), .A3(new_n328), .A4(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT96), .B(G478), .ZN(new_n559));
  INV_X1    g373(.A(new_n370), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n559), .B1(new_n560), .B2(G902), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n337), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n553), .A2(new_n443), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT34), .B(G104), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(G6));
  AND3_X1   g380(.A1(new_n331), .A2(new_n332), .A3(new_n336), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n374), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT97), .B1(new_n443), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n337), .A2(new_n373), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n281), .A2(new_n570), .A3(new_n571), .A4(new_n385), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n552), .A3(new_n545), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT35), .B(G107), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT98), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n574), .B(new_n576), .ZN(G9));
  NOR2_X1   g391(.A1(new_n550), .A2(new_n551), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n517), .A2(new_n524), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n579), .B(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n542), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n541), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n440), .A2(new_n447), .A3(new_n578), .A4(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT37), .Z(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G110), .ZN(G12));
  AND2_X1   g404(.A1(new_n502), .A2(new_n281), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n439), .B1(new_n541), .B2(new_n586), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n378), .B1(G900), .B2(new_n382), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n571), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G128), .ZN(G30));
  AND2_X1   g411(.A1(new_n488), .A2(new_n489), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n471), .A2(new_n472), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n469), .B2(new_n491), .ZN(new_n600));
  OAI21_X1  g414(.A(G472), .B1(new_n600), .B2(G902), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n587), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n373), .A2(new_n188), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n337), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n594), .B(KEYINPUT39), .Z(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n445), .A2(KEYINPUT40), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n439), .B2(new_n605), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n279), .A2(new_n280), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT38), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n602), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT102), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G143), .ZN(G45));
  NAND3_X1  g430(.A1(new_n562), .A2(new_n337), .A3(new_n594), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n593), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G146), .ZN(G48));
  OAI21_X1  g434(.A(new_n328), .B1(new_n418), .B2(new_n427), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(G469), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n622), .A2(new_n428), .A3(new_n437), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n443), .A2(new_n563), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n502), .A2(new_n545), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT41), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G113), .ZN(G15));
  NAND4_X1  g441(.A1(new_n573), .A2(new_n502), .A3(new_n545), .A4(new_n623), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT103), .B(G116), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G18));
  AND3_X1   g444(.A1(new_n587), .A2(new_n375), .A3(new_n385), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n502), .A2(new_n631), .A3(new_n281), .A4(new_n623), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G119), .ZN(G21));
  NOR2_X1   g447(.A1(new_n441), .A2(new_n442), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT105), .B1(new_n634), .B2(new_n604), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT105), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n611), .A2(new_n603), .A3(new_n636), .A4(new_n337), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n622), .A2(new_n428), .ZN(new_n639));
  INV_X1    g453(.A(new_n437), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n639), .A2(new_n640), .A3(new_n384), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n484), .A2(new_n328), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n469), .B1(new_n492), .B2(new_n477), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n473), .A2(new_n643), .A3(new_n482), .A4(new_n483), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n485), .B(KEYINPUT104), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n642), .A2(G472), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n638), .A2(new_n641), .A3(new_n545), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G122), .ZN(G24));
  NAND2_X1  g462(.A1(new_n644), .A2(new_n645), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n460), .A2(new_n470), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT68), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n460), .A2(new_n461), .A3(new_n470), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n479), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n482), .A2(new_n483), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(G902), .B1(new_n655), .B2(new_n478), .ZN(new_n656));
  INV_X1    g470(.A(G472), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n587), .B(new_n649), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT106), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n646), .A2(new_n660), .A3(new_n587), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n618), .A2(new_n623), .A3(new_n281), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT107), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n662), .A2(new_n667), .A3(new_n664), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G125), .ZN(G27));
  AND2_X1   g484(.A1(new_n502), .A2(new_n545), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n634), .A2(new_n437), .A3(new_n187), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n433), .A2(KEYINPUT108), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT108), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n431), .A2(new_n674), .A3(new_n432), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n673), .A2(G469), .A3(new_n434), .A4(new_n675), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n676), .A2(new_n428), .A3(new_n430), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n671), .A2(new_n618), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT110), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT32), .B1(new_n484), .B2(new_n485), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT109), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n501), .A2(new_n489), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n544), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n672), .A2(new_n677), .A3(new_n617), .A4(new_n680), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n488), .A2(KEYINPUT109), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n685), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  AND4_X1   g506(.A1(new_n682), .A2(new_n687), .A3(new_n692), .A4(new_n545), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n681), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G131), .ZN(G33));
  NAND3_X1  g509(.A1(new_n671), .A2(new_n595), .A3(new_n678), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G134), .ZN(G36));
  NAND4_X1  g511(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n434), .A4(new_n675), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n433), .A2(new_n434), .ZN(new_n699));
  OAI211_X1 g513(.A(new_n698), .B(G469), .C1(KEYINPUT45), .C2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(KEYINPUT46), .B1(new_n700), .B2(new_n430), .ZN(new_n701));
  INV_X1    g515(.A(new_n428), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(KEYINPUT46), .A3(new_n430), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n437), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n605), .ZN(new_n707));
  INV_X1    g521(.A(new_n562), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n709));
  OAI22_X1  g523(.A1(new_n708), .A2(new_n337), .B1(KEYINPUT111), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n711));
  NAND3_X1  g525(.A1(new_n562), .A2(new_n567), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g527(.A(new_n713), .B(new_n587), .C1(new_n550), .C2(new_n551), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(KEYINPUT44), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n611), .A2(new_n188), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT112), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n707), .A2(new_n716), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G137), .ZN(G39));
  XOR2_X1   g536(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n723));
  OR2_X1    g537(.A1(new_n706), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n725), .B1(new_n705), .B2(new_n437), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n502), .A2(new_n545), .A3(new_n617), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n718), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G140), .ZN(G42));
  AND2_X1   g544(.A1(new_n598), .A2(new_n601), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n545), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n639), .B(KEYINPUT49), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n562), .A2(new_n567), .A3(new_n438), .A4(new_n187), .ZN(new_n734));
  OR4_X1    g548(.A1(new_n612), .A2(new_n732), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n646), .A2(new_n545), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n378), .B1(new_n710), .B2(new_n712), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT115), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(KEYINPUT115), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n737), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n612), .A2(new_n187), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n623), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n741), .A2(KEYINPUT50), .A3(new_n623), .A4(new_n742), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n706), .A2(new_n723), .ZN(new_n748));
  OAI22_X1  g562(.A1(new_n748), .A2(new_n726), .B1(new_n438), .B2(new_n639), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n741), .A2(new_n720), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n740), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n672), .A2(new_n639), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n661), .B2(new_n659), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n747), .A2(new_n751), .A3(new_n757), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n545), .A2(new_n731), .A3(new_n379), .A4(new_n754), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n567), .A3(new_n708), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT116), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n759), .A2(new_n762), .A3(new_n567), .A4(new_n708), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n736), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n756), .B1(new_n749), .B2(new_n750), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(KEYINPUT51), .A3(new_n764), .A4(new_n747), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n766), .A2(new_n376), .A3(new_n768), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n502), .A2(new_n592), .A3(new_n375), .A4(new_n594), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n672), .A2(new_n677), .A3(new_n617), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n770), .A2(new_n718), .B1(new_n662), .B2(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(KEYINPUT53), .A2(new_n694), .A3(new_n696), .A4(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n628), .A2(new_n632), .A3(new_n647), .A4(new_n625), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT114), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n563), .A2(new_n568), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n552), .A2(new_n545), .A3(new_n444), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n546), .A2(new_n588), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n591), .B(new_n592), .C1(new_n595), .C2(new_n618), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n677), .A2(new_n640), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n602), .A2(new_n594), .A3(new_n638), .A4(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n669), .A2(KEYINPUT52), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n667), .B1(new_n662), .B2(new_n664), .ZN(new_n784));
  AOI211_X1 g598(.A(KEYINPUT107), .B(new_n663), .C1(new_n659), .C2(new_n661), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n780), .B(new_n782), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n773), .A2(new_n779), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n778), .A2(new_n774), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n694), .A2(new_n791), .A3(new_n696), .A4(new_n772), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT53), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n741), .A2(new_n281), .A3(new_n623), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n789), .A2(new_n792), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n800), .B2(new_n793), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n769), .A2(new_n796), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  NOR4_X1   g616(.A1(new_n732), .A2(new_n378), .A3(new_n563), .A4(new_n753), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n752), .A2(new_n686), .A3(new_n754), .ZN(new_n804));
  XOR2_X1   g618(.A(new_n804), .B(KEYINPUT48), .Z(new_n805));
  NOR3_X1   g619(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(G952), .A2(G953), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n735), .B1(new_n806), .B2(new_n807), .ZN(G75));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n798), .A2(new_n799), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n773), .A2(new_n779), .A3(new_n789), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n328), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n812), .B2(G210), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n230), .B(new_n262), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT117), .Z(new_n815));
  XOR2_X1   g629(.A(new_n815), .B(KEYINPUT55), .Z(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n809), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(G210), .B(G902), .C1(new_n790), .C2(new_n793), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT56), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n821), .A2(KEYINPUT118), .A3(new_n816), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n283), .A2(G952), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n820), .A3(new_n817), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n819), .A2(KEYINPUT119), .A3(new_n820), .A4(new_n817), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n824), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n823), .A2(new_n829), .ZN(G51));
  NAND2_X1  g644(.A1(new_n430), .A2(KEYINPUT57), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n794), .A2(new_n795), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n810), .A2(new_n811), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n831), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n430), .A2(KEYINPUT57), .ZN(new_n836));
  OAI22_X1  g650(.A1(new_n835), .A2(new_n836), .B1(new_n418), .B2(new_n427), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n794), .A2(new_n328), .A3(new_n700), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n824), .B1(new_n837), .B2(new_n838), .ZN(G54));
  NAND3_X1  g653(.A1(new_n812), .A2(KEYINPUT58), .A3(G475), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n325), .A3(new_n314), .ZN(new_n841));
  INV_X1    g655(.A(new_n824), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n812), .A2(KEYINPUT58), .A3(G475), .A4(new_n326), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(G60));
  NOR2_X1   g658(.A1(new_n832), .A2(new_n834), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n556), .A2(new_n557), .ZN(new_n846));
  NAND2_X1  g660(.A1(G478), .A2(G902), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT59), .Z(new_n848));
  NOR3_X1   g662(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n796), .B2(new_n801), .ZN(new_n850));
  INV_X1    g664(.A(new_n846), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n849), .A2(new_n852), .ZN(G63));
  XNOR2_X1  g667(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n365), .A2(new_n328), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n833), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n533), .A2(new_n534), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n833), .A2(new_n585), .A3(new_n584), .A4(new_n856), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n859), .A2(new_n842), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(G66));
  OAI21_X1  g677(.A(G953), .B1(new_n381), .B2(new_n260), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n791), .B2(G953), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT121), .Z(new_n866));
  OAI221_X1 g680(.A(new_n223), .B1(G898), .B2(new_n283), .C1(new_n228), .C2(new_n229), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n866), .B(new_n867), .ZN(G69));
  NAND3_X1  g682(.A1(new_n707), .A2(new_n638), .A3(new_n686), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n729), .A2(new_n721), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n694), .A2(new_n696), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(KEYINPUT122), .B(new_n780), .C1(new_n784), .C2(new_n785), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n870), .A2(new_n871), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n283), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n457), .A2(new_n459), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n308), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n877), .B(new_n879), .C1(G227), .C2(new_n283), .ZN(new_n880));
  OAI21_X1  g694(.A(G900), .B1(new_n879), .B2(G227), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(G953), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n874), .A2(new_n614), .A3(new_n875), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n874), .A2(KEYINPUT62), .A3(new_n614), .A4(new_n875), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n439), .A2(new_n605), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n671), .A2(new_n888), .A3(new_n718), .A4(new_n776), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n729), .A2(new_n721), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT123), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n893), .B(new_n890), .C1(new_n885), .C2(new_n886), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n283), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n880), .B(new_n882), .C1(new_n895), .C2(new_n879), .ZN(G72));
  NAND2_X1  g710(.A1(G472), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT63), .Z(new_n898));
  INV_X1    g712(.A(new_n791), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n876), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n498), .B(KEYINPUT125), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n469), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT126), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n498), .A2(new_n468), .ZN(new_n905));
  OAI221_X1 g719(.A(new_n898), .B1(new_n599), .B2(new_n905), .C1(new_n800), .C2(new_n793), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n906), .A3(new_n842), .ZN(new_n907));
  INV_X1    g721(.A(new_n898), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n892), .A2(new_n894), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n791), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n901), .B1(new_n910), .B2(KEYINPUT124), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n887), .A2(new_n891), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n893), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n887), .A2(KEYINPUT123), .A3(new_n891), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n791), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n898), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n469), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n907), .B1(new_n911), .B2(new_n918), .ZN(G57));
endmodule


