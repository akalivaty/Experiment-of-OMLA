

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(n694), .A2(n792), .ZN(n728) );
  BUF_X1 U553 ( .A(n554), .Z(n889) );
  INV_X1 U554 ( .A(n728), .ZN(n722) );
  NOR2_X2 U555 ( .A1(G2104), .A2(n540), .ZN(n893) );
  AND2_X1 U556 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U557 ( .A(n756), .B(n755), .ZN(n757) );
  AND2_X1 U558 ( .A1(n541), .A2(G2104), .ZN(n555) );
  BUF_X1 U559 ( .A(n555), .Z(n890) );
  NAND2_X1 U560 ( .A1(n778), .A2(n519), .ZN(n816) );
  INV_X1 U561 ( .A(n820), .ZN(n813) );
  OR2_X1 U562 ( .A1(n775), .A2(n767), .ZN(n518) );
  AND2_X1 U563 ( .A1(n777), .A2(n776), .ZN(n519) );
  AND2_X1 U564 ( .A1(n768), .A2(n518), .ZN(n520) );
  XOR2_X1 U565 ( .A(n733), .B(KEYINPUT103), .Z(n521) );
  XOR2_X1 U566 ( .A(n702), .B(KEYINPUT102), .Z(n522) );
  INV_X1 U567 ( .A(KEYINPUT26), .ZN(n696) );
  NOR2_X1 U568 ( .A1(n700), .A2(n978), .ZN(n701) );
  NOR2_X1 U569 ( .A1(G168), .A2(n732), .ZN(n733) );
  AND2_X1 U570 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U571 ( .A1(G2084), .A2(n728), .ZN(n729) );
  NOR2_X1 U572 ( .A1(n521), .A2(n736), .ZN(n737) );
  NOR2_X1 U573 ( .A1(G1966), .A2(n775), .ZN(n750) );
  INV_X1 U574 ( .A(n973), .ZN(n760) );
  INV_X1 U575 ( .A(KEYINPUT105), .ZN(n755) );
  INV_X1 U576 ( .A(KEYINPUT23), .ZN(n542) );
  NOR2_X1 U577 ( .A1(G164), .A2(G1384), .ZN(n792) );
  INV_X1 U578 ( .A(G2105), .ZN(n540) );
  AND2_X1 U579 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U580 ( .A1(n553), .A2(n552), .ZN(n693) );
  BUF_X1 U581 ( .A(n693), .Z(G160) );
  NOR2_X1 U582 ( .A1(G543), .A2(G651), .ZN(n654) );
  NAND2_X1 U583 ( .A1(G89), .A2(n654), .ZN(n523) );
  XOR2_X1 U584 ( .A(KEYINPUT77), .B(n523), .Z(n524) );
  XNOR2_X1 U585 ( .A(n524), .B(KEYINPUT4), .ZN(n527) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n647) );
  XNOR2_X1 U587 ( .A(G651), .B(KEYINPUT69), .ZN(n531) );
  NOR2_X1 U588 ( .A1(n647), .A2(n531), .ZN(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT70), .B(n525), .ZN(n658) );
  NAND2_X1 U590 ( .A1(G76), .A2(n658), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT5), .ZN(n538) );
  NOR2_X1 U593 ( .A1(n647), .A2(G651), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT65), .B(n529), .Z(n657) );
  NAND2_X1 U595 ( .A1(n657), .A2(G51), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(KEYINPUT78), .ZN(n535) );
  NOR2_X1 U597 ( .A1(G543), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(KEYINPUT1), .B(KEYINPUT71), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n653) );
  NAND2_X1 U600 ( .A1(G63), .A2(n653), .ZN(n534) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(KEYINPUT6), .B(n536), .Z(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U605 ( .A1(n893), .A2(G125), .ZN(n545) );
  INV_X1 U606 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n555), .A2(G101), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n546), .B(KEYINPUT66), .ZN(n547) );
  INV_X1 U611 ( .A(n547), .ZN(n550) );
  NOR2_X1 U612 ( .A1(G2105), .A2(G2104), .ZN(n548) );
  XOR2_X1 U613 ( .A(KEYINPUT17), .B(n548), .Z(n554) );
  NAND2_X1 U614 ( .A1(n554), .A2(G137), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n553) );
  AND2_X1 U616 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  NAND2_X1 U617 ( .A1(G113), .A2(n894), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT67), .B(n551), .ZN(n552) );
  NAND2_X1 U619 ( .A1(G138), .A2(n889), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G102), .A2(n890), .ZN(n556) );
  NAND2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U622 ( .A1(G126), .A2(n893), .ZN(n559) );
  NAND2_X1 U623 ( .A1(G114), .A2(n894), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U625 ( .A1(n561), .A2(n560), .ZN(G164) );
  NAND2_X1 U626 ( .A1(G64), .A2(n653), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G52), .A2(n657), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G90), .A2(n654), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G77), .A2(n658), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT9), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT74), .B(n567), .Z(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(G171) );
  AND2_X1 U635 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U636 ( .A1(n893), .A2(G123), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT18), .ZN(n572) );
  NAND2_X1 U638 ( .A1(G135), .A2(n889), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(KEYINPUT80), .B(n573), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G99), .A2(n890), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G111), .A2(n894), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n925) );
  XNOR2_X1 U645 ( .A(n925), .B(G2096), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n578), .B(KEYINPUT81), .ZN(n579) );
  OR2_X1 U647 ( .A1(G2100), .A2(n579), .ZN(G156) );
  INV_X1 U648 ( .A(G120), .ZN(G236) );
  INV_X1 U649 ( .A(G69), .ZN(G235) );
  INV_X1 U650 ( .A(G108), .ZN(G238) );
  INV_X1 U651 ( .A(G132), .ZN(G219) );
  INV_X1 U652 ( .A(G82), .ZN(G220) );
  NAND2_X1 U653 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U654 ( .A(n580), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U655 ( .A(G223), .ZN(n840) );
  NAND2_X1 U656 ( .A1(n840), .A2(G567), .ZN(n581) );
  XNOR2_X1 U657 ( .A(n581), .B(KEYINPUT11), .ZN(n582) );
  XNOR2_X1 U658 ( .A(KEYINPUT75), .B(n582), .ZN(G234) );
  NAND2_X1 U659 ( .A1(G56), .A2(n653), .ZN(n583) );
  XOR2_X1 U660 ( .A(KEYINPUT14), .B(n583), .Z(n589) );
  NAND2_X1 U661 ( .A1(n654), .A2(G81), .ZN(n584) );
  XNOR2_X1 U662 ( .A(n584), .B(KEYINPUT12), .ZN(n586) );
  NAND2_X1 U663 ( .A1(G68), .A2(n658), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U665 ( .A(KEYINPUT13), .B(n587), .Z(n588) );
  NOR2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n657), .A2(G43), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n978) );
  INV_X1 U669 ( .A(n978), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n592), .A2(G860), .ZN(G153) );
  INV_X1 U671 ( .A(G171), .ZN(G301) );
  NAND2_X1 U672 ( .A1(G66), .A2(n653), .ZN(n594) );
  NAND2_X1 U673 ( .A1(G92), .A2(n654), .ZN(n593) );
  NAND2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G54), .A2(n657), .ZN(n596) );
  NAND2_X1 U676 ( .A1(G79), .A2(n658), .ZN(n595) );
  NAND2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U678 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X1 U679 ( .A(KEYINPUT15), .B(n599), .Z(n981) );
  NOR2_X1 U680 ( .A1(n981), .A2(G868), .ZN(n600) );
  XOR2_X1 U681 ( .A(KEYINPUT76), .B(n600), .Z(n602) );
  NAND2_X1 U682 ( .A1(G868), .A2(G301), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(G284) );
  XOR2_X1 U684 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U685 ( .A1(G65), .A2(n653), .ZN(n604) );
  NAND2_X1 U686 ( .A1(G53), .A2(n657), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G91), .A2(n654), .ZN(n606) );
  NAND2_X1 U689 ( .A1(G78), .A2(n658), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n970) );
  INV_X1 U692 ( .A(n970), .ZN(G299) );
  INV_X1 U693 ( .A(G868), .ZN(n609) );
  NOR2_X1 U694 ( .A1(G286), .A2(n609), .ZN(n611) );
  NOR2_X1 U695 ( .A1(G868), .A2(G299), .ZN(n610) );
  NOR2_X1 U696 ( .A1(n611), .A2(n610), .ZN(G297) );
  INV_X1 U697 ( .A(G559), .ZN(n612) );
  NOR2_X1 U698 ( .A1(G860), .A2(n612), .ZN(n613) );
  XNOR2_X1 U699 ( .A(KEYINPUT79), .B(n613), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n614), .A2(n981), .ZN(n615) );
  XNOR2_X1 U701 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U702 ( .A1(G868), .A2(n978), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n981), .A2(G868), .ZN(n616) );
  NOR2_X1 U704 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U705 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U706 ( .A1(G93), .A2(n654), .ZN(n620) );
  NAND2_X1 U707 ( .A1(G80), .A2(n658), .ZN(n619) );
  NAND2_X1 U708 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U709 ( .A(n621), .B(KEYINPUT83), .ZN(n623) );
  NAND2_X1 U710 ( .A1(G67), .A2(n653), .ZN(n622) );
  NAND2_X1 U711 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n657), .A2(G55), .ZN(n624) );
  XOR2_X1 U713 ( .A(KEYINPUT84), .B(n624), .Z(n625) );
  NOR2_X1 U714 ( .A1(n626), .A2(n625), .ZN(n670) );
  NAND2_X1 U715 ( .A1(G559), .A2(n981), .ZN(n627) );
  XNOR2_X1 U716 ( .A(n627), .B(n978), .ZN(n672) );
  NOR2_X1 U717 ( .A1(G860), .A2(n672), .ZN(n629) );
  XNOR2_X1 U718 ( .A(KEYINPUT82), .B(KEYINPUT85), .ZN(n628) );
  XNOR2_X1 U719 ( .A(n629), .B(n628), .ZN(n630) );
  XOR2_X1 U720 ( .A(n670), .B(n630), .Z(G145) );
  NAND2_X1 U721 ( .A1(G60), .A2(n653), .ZN(n631) );
  XNOR2_X1 U722 ( .A(n631), .B(KEYINPUT72), .ZN(n638) );
  NAND2_X1 U723 ( .A1(G47), .A2(n657), .ZN(n633) );
  NAND2_X1 U724 ( .A1(G72), .A2(n658), .ZN(n632) );
  NAND2_X1 U725 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U726 ( .A1(n654), .A2(G85), .ZN(n634) );
  XOR2_X1 U727 ( .A(KEYINPUT68), .B(n634), .Z(n635) );
  NOR2_X1 U728 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U729 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U730 ( .A(KEYINPUT73), .B(n639), .Z(G290) );
  NAND2_X1 U731 ( .A1(G61), .A2(n653), .ZN(n641) );
  NAND2_X1 U732 ( .A1(G86), .A2(n654), .ZN(n640) );
  NAND2_X1 U733 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n658), .A2(G73), .ZN(n642) );
  XOR2_X1 U735 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U736 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U737 ( .A1(n657), .A2(G48), .ZN(n645) );
  NAND2_X1 U738 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U739 ( .A1(G49), .A2(n657), .ZN(n649) );
  NAND2_X1 U740 ( .A1(G87), .A2(n647), .ZN(n648) );
  NAND2_X1 U741 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U742 ( .A1(n653), .A2(n650), .ZN(n652) );
  NAND2_X1 U743 ( .A1(G651), .A2(G74), .ZN(n651) );
  NAND2_X1 U744 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U745 ( .A1(G62), .A2(n653), .ZN(n656) );
  NAND2_X1 U746 ( .A1(G88), .A2(n654), .ZN(n655) );
  NAND2_X1 U747 ( .A1(n656), .A2(n655), .ZN(n662) );
  NAND2_X1 U748 ( .A1(G50), .A2(n657), .ZN(n660) );
  NAND2_X1 U749 ( .A1(G75), .A2(n658), .ZN(n659) );
  NAND2_X1 U750 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U751 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U752 ( .A(KEYINPUT86), .B(n663), .Z(G303) );
  NOR2_X1 U753 ( .A1(G868), .A2(n670), .ZN(n664) );
  XOR2_X1 U754 ( .A(n664), .B(KEYINPUT88), .Z(n675) );
  XOR2_X1 U755 ( .A(KEYINPUT19), .B(KEYINPUT87), .Z(n665) );
  XNOR2_X1 U756 ( .A(G288), .B(n665), .ZN(n666) );
  XNOR2_X1 U757 ( .A(G305), .B(n666), .ZN(n668) );
  XNOR2_X1 U758 ( .A(n970), .B(G303), .ZN(n667) );
  XNOR2_X1 U759 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U760 ( .A(n670), .B(n669), .Z(n671) );
  XNOR2_X1 U761 ( .A(G290), .B(n671), .ZN(n907) );
  XNOR2_X1 U762 ( .A(n907), .B(n672), .ZN(n673) );
  NAND2_X1 U763 ( .A1(G868), .A2(n673), .ZN(n674) );
  NAND2_X1 U764 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U765 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U766 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U767 ( .A1(G2090), .A2(n677), .ZN(n679) );
  XOR2_X1 U768 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n678) );
  XNOR2_X1 U769 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U770 ( .A1(G2072), .A2(n680), .ZN(G158) );
  XNOR2_X1 U771 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n681) );
  XNOR2_X1 U773 ( .A(KEYINPUT22), .B(n681), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n682), .A2(G96), .ZN(n683) );
  NOR2_X1 U775 ( .A1(G218), .A2(n683), .ZN(n684) );
  XOR2_X1 U776 ( .A(KEYINPUT90), .B(n684), .Z(n847) );
  NAND2_X1 U777 ( .A1(n847), .A2(G2106), .ZN(n689) );
  NOR2_X1 U778 ( .A1(G235), .A2(G236), .ZN(n685) );
  XNOR2_X1 U779 ( .A(n685), .B(KEYINPUT91), .ZN(n686) );
  NOR2_X1 U780 ( .A1(G238), .A2(n686), .ZN(n687) );
  NAND2_X1 U781 ( .A1(G57), .A2(n687), .ZN(n846) );
  NAND2_X1 U782 ( .A1(G567), .A2(n846), .ZN(n688) );
  NAND2_X1 U783 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U784 ( .A(KEYINPUT92), .B(n690), .Z(G319) );
  INV_X1 U785 ( .A(G319), .ZN(n692) );
  NAND2_X1 U786 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n845) );
  NAND2_X1 U788 ( .A1(n845), .A2(G36), .ZN(G176) );
  NAND2_X1 U789 ( .A1(G40), .A2(n693), .ZN(n790) );
  XNOR2_X1 U790 ( .A(n790), .B(KEYINPUT93), .ZN(n694) );
  INV_X1 U791 ( .A(G1996), .ZN(n695) );
  NOR2_X1 U792 ( .A1(n728), .A2(n695), .ZN(n697) );
  XNOR2_X1 U793 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n728), .A2(G1341), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U796 ( .A(n701), .B(KEYINPUT64), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n703), .A2(n981), .ZN(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n981), .ZN(n707) );
  NOR2_X1 U799 ( .A1(G2067), .A2(n728), .ZN(n705) );
  NOR2_X1 U800 ( .A1(n722), .A2(G1348), .ZN(n704) );
  NOR2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n722), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U804 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  AND2_X1 U805 ( .A1(G1956), .A2(n728), .ZN(n709) );
  NOR2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n970), .A2(n716), .ZN(n712) );
  XNOR2_X1 U808 ( .A(KEYINPUT101), .B(KEYINPUT28), .ZN(n711) );
  XNOR2_X1 U809 ( .A(n712), .B(n711), .ZN(n715) );
  AND2_X1 U810 ( .A1(n713), .A2(n715), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n522), .A2(n714), .ZN(n720) );
  INV_X1 U812 ( .A(n715), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n970), .A2(n716), .ZN(n717) );
  OR2_X1 U814 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U815 ( .A(n721), .B(KEYINPUT29), .ZN(n727) );
  NOR2_X1 U816 ( .A1(n722), .A2(G1961), .ZN(n723) );
  XNOR2_X1 U817 ( .A(n723), .B(KEYINPUT100), .ZN(n725) );
  XOR2_X1 U818 ( .A(KEYINPUT25), .B(G2078), .Z(n951) );
  NOR2_X1 U819 ( .A1(n728), .A2(n951), .ZN(n724) );
  NOR2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n734) );
  NOR2_X1 U821 ( .A1(G301), .A2(n734), .ZN(n726) );
  NOR2_X1 U822 ( .A1(n727), .A2(n726), .ZN(n739) );
  NAND2_X1 U823 ( .A1(G8), .A2(n728), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n729), .B(KEYINPUT99), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n751), .A2(G8), .ZN(n730) );
  NOR2_X1 U826 ( .A1(n750), .A2(n730), .ZN(n731) );
  XOR2_X1 U827 ( .A(KEYINPUT30), .B(n731), .Z(n732) );
  NAND2_X1 U828 ( .A1(n734), .A2(G301), .ZN(n735) );
  XOR2_X1 U829 ( .A(KEYINPUT104), .B(n735), .Z(n736) );
  XNOR2_X1 U830 ( .A(n737), .B(KEYINPUT31), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n749) );
  INV_X1 U832 ( .A(n749), .ZN(n740) );
  NAND2_X1 U833 ( .A1(n740), .A2(G286), .ZN(n746) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n775), .ZN(n742) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n728), .ZN(n741) );
  NOR2_X1 U836 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U837 ( .A(KEYINPUT106), .B(n743), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n744), .A2(G303), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U840 ( .A1(n747), .A2(G8), .ZN(n748) );
  XNOR2_X1 U841 ( .A(n748), .B(KEYINPUT32), .ZN(n758) );
  NOR2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n754) );
  INV_X1 U843 ( .A(n751), .ZN(n752) );
  NAND2_X1 U844 ( .A1(G8), .A2(n752), .ZN(n753) );
  NAND2_X1 U845 ( .A1(n754), .A2(n753), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n758), .A2(n757), .ZN(n771) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U848 ( .A1(G303), .A2(G1971), .ZN(n759) );
  NOR2_X1 U849 ( .A1(n766), .A2(n759), .ZN(n980) );
  NAND2_X1 U850 ( .A1(n771), .A2(n980), .ZN(n762) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n973) );
  NOR2_X1 U852 ( .A1(n775), .A2(n760), .ZN(n761) );
  NAND2_X1 U853 ( .A1(n762), .A2(n761), .ZN(n764) );
  INV_X1 U854 ( .A(KEYINPUT33), .ZN(n763) );
  XNOR2_X1 U855 ( .A(n765), .B(KEYINPUT107), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n766), .A2(KEYINPUT33), .ZN(n767) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n985) );
  NAND2_X1 U858 ( .A1(n520), .A2(n985), .ZN(n778) );
  NOR2_X1 U859 ( .A1(G2090), .A2(G303), .ZN(n769) );
  NAND2_X1 U860 ( .A1(G8), .A2(n769), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n772), .A2(n775), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G1981), .A2(G305), .ZN(n773) );
  XOR2_X1 U864 ( .A(n773), .B(KEYINPUT24), .Z(n774) );
  OR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U866 ( .A(G1986), .B(G290), .Z(n974) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NAND2_X1 U868 ( .A1(n894), .A2(G116), .ZN(n779) );
  XOR2_X1 U869 ( .A(KEYINPUT95), .B(n779), .Z(n781) );
  NAND2_X1 U870 ( .A1(n893), .A2(G128), .ZN(n780) );
  NAND2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U872 ( .A(KEYINPUT35), .B(n782), .ZN(n788) );
  NAND2_X1 U873 ( .A1(G140), .A2(n889), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G104), .A2(n890), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n786) );
  XOR2_X1 U876 ( .A(KEYINPUT94), .B(KEYINPUT34), .Z(n785) );
  XNOR2_X1 U877 ( .A(n786), .B(n785), .ZN(n787) );
  NAND2_X1 U878 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U879 ( .A(KEYINPUT36), .B(n789), .Z(n904) );
  OR2_X1 U880 ( .A1(n824), .A2(n904), .ZN(n924) );
  NAND2_X1 U881 ( .A1(n974), .A2(n924), .ZN(n793) );
  XOR2_X1 U882 ( .A(n790), .B(KEYINPUT93), .Z(n791) );
  NOR2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n826) );
  NAND2_X1 U884 ( .A1(n793), .A2(n826), .ZN(n814) );
  NAND2_X1 U885 ( .A1(n890), .A2(G105), .ZN(n794) );
  XNOR2_X1 U886 ( .A(n794), .B(KEYINPUT38), .ZN(n796) );
  NAND2_X1 U887 ( .A1(G117), .A2(n894), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G129), .A2(n893), .ZN(n797) );
  XNOR2_X1 U890 ( .A(KEYINPUT97), .B(n797), .ZN(n798) );
  NOR2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U892 ( .A(n800), .B(KEYINPUT98), .ZN(n802) );
  NAND2_X1 U893 ( .A1(G141), .A2(n889), .ZN(n801) );
  NAND2_X1 U894 ( .A1(n802), .A2(n801), .ZN(n874) );
  NAND2_X1 U895 ( .A1(n874), .A2(G1996), .ZN(n811) );
  NAND2_X1 U896 ( .A1(G95), .A2(n890), .ZN(n804) );
  NAND2_X1 U897 ( .A1(G107), .A2(n894), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n889), .A2(G131), .ZN(n805) );
  XOR2_X1 U900 ( .A(KEYINPUT96), .B(n805), .Z(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U902 ( .A1(n893), .A2(G119), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n873) );
  NAND2_X1 U904 ( .A1(n873), .A2(G1991), .ZN(n810) );
  AND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n935) );
  INV_X1 U906 ( .A(n826), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n935), .A2(n812), .ZN(n820) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n829) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n874), .ZN(n930) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n873), .ZN(n926) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT108), .B(n817), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n926), .A2(n818), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n930), .A2(n821), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n822), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n924), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n824), .A2(n904), .ZN(n923) );
  NAND2_X1 U919 ( .A1(n825), .A2(n923), .ZN(n827) );
  NAND2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U922 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U923 ( .A(G1341), .B(G2454), .ZN(n831) );
  XNOR2_X1 U924 ( .A(n831), .B(G2430), .ZN(n832) );
  XNOR2_X1 U925 ( .A(n832), .B(G1348), .ZN(n838) );
  XOR2_X1 U926 ( .A(G2443), .B(G2427), .Z(n834) );
  XNOR2_X1 U927 ( .A(G2438), .B(G2446), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(n836) );
  XOR2_X1 U929 ( .A(G2451), .B(G2435), .Z(n835) );
  XNOR2_X1 U930 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U931 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U932 ( .A1(n839), .A2(G14), .ZN(n912) );
  XNOR2_X1 U933 ( .A(KEYINPUT109), .B(n912), .ZN(G401) );
  NAND2_X1 U934 ( .A1(G2106), .A2(n840), .ZN(G217) );
  INV_X1 U935 ( .A(G661), .ZN(n842) );
  NAND2_X1 U936 ( .A1(G2), .A2(G15), .ZN(n841) );
  NOR2_X1 U937 ( .A1(n842), .A2(n841), .ZN(n843) );
  XOR2_X1 U938 ( .A(KEYINPUT110), .B(n843), .Z(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(G188) );
  XNOR2_X1 U941 ( .A(G96), .B(KEYINPUT111), .ZN(G221) );
  NOR2_X1 U943 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U944 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U945 ( .A(G1956), .B(KEYINPUT41), .ZN(n857) );
  XOR2_X1 U946 ( .A(G1986), .B(G1976), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1961), .B(G1971), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(G1991), .B(G1981), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1996), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT112), .B(G2474), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(G229) );
  XOR2_X1 U956 ( .A(G2100), .B(G2096), .Z(n859) );
  XNOR2_X1 U957 ( .A(KEYINPUT42), .B(G2678), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U959 ( .A(KEYINPUT43), .B(G2090), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U962 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U963 ( .A(G2078), .B(G2084), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U965 ( .A1(n893), .A2(G124), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G112), .A2(n894), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G136), .A2(n889), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G100), .A2(n890), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U972 ( .A1(n872), .A2(n871), .ZN(G162) );
  XNOR2_X1 U973 ( .A(G160), .B(n925), .ZN(n903) );
  XNOR2_X1 U974 ( .A(G164), .B(n873), .ZN(n877) );
  XNOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n888) );
  NAND2_X1 U978 ( .A1(G130), .A2(n893), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G118), .A2(n894), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n886) );
  XNOR2_X1 U981 ( .A(KEYINPUT45), .B(KEYINPUT114), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n889), .A2(G142), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n890), .A2(G106), .ZN(n880) );
  XOR2_X1 U984 ( .A(KEYINPUT113), .B(n880), .Z(n881) );
  NAND2_X1 U985 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U986 ( .A(n884), .B(n883), .Z(n885) );
  NOR2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U988 ( .A(n888), .B(n887), .Z(n901) );
  NAND2_X1 U989 ( .A1(G139), .A2(n889), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G103), .A2(n890), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U992 ( .A1(G127), .A2(n893), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G115), .A2(n894), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n897), .Z(n898) );
  NOR2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n919) );
  XNOR2_X1 U997 ( .A(n919), .B(G162), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U1002 ( .A(n907), .B(G286), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G171), .B(n981), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n910), .B(n978), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n911), .ZN(G397) );
  NAND2_X1 U1007 ( .A1(n912), .A2(G319), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1012 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1015 ( .A(G164), .B(G2078), .Z(n918) );
  XNOR2_X1 U1016 ( .A(KEYINPUT116), .B(n918), .ZN(n921) );
  XOR2_X1 U1017 ( .A(G2072), .B(n919), .Z(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1019 ( .A(KEYINPUT50), .B(n922), .Z(n940) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n937) );
  NOR2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n933) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(n931), .B(KEYINPUT51), .ZN(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(KEYINPUT115), .B(n938), .ZN(n939) );
  NOR2_X1 U1031 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n941), .ZN(n943) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n942) );
  NAND2_X1 U1034 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1035 ( .A1(n944), .A2(G29), .ZN(n945) );
  XNOR2_X1 U1036 ( .A(n945), .B(KEYINPUT117), .ZN(n968) );
  XNOR2_X1 U1037 ( .A(G2090), .B(G35), .ZN(n961) );
  XOR2_X1 U1038 ( .A(G2072), .B(G33), .Z(n948) );
  XOR2_X1 U1039 ( .A(KEYINPUT118), .B(G26), .Z(n946) );
  XNOR2_X1 U1040 ( .A(n946), .B(G2067), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT119), .B(n949), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(G28), .ZN(n958) );
  XOR2_X1 U1044 ( .A(G1991), .B(G25), .Z(n956) );
  XNOR2_X1 U1045 ( .A(n951), .B(G27), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G32), .B(G1996), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(n954), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n959), .ZN(n960) );
  NOR2_X1 U1052 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n962), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1056 ( .A(KEYINPUT55), .B(n965), .ZN(n966) );
  NOR2_X1 U1057 ( .A1(n966), .A2(G29), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n969), .ZN(n1025) );
  XNOR2_X1 U1060 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1061 ( .A(n970), .B(G1956), .ZN(n972) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n976) );
  NAND2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1065 ( .A1(n976), .A2(n975), .ZN(n993) );
  XOR2_X1 U1066 ( .A(G1341), .B(KEYINPUT122), .Z(n977) );
  XNOR2_X1 U1067 ( .A(n978), .B(n977), .ZN(n979) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n991) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n981), .ZN(n983) );
  XNOR2_X1 U1070 ( .A(G171), .B(G1961), .ZN(n982) );
  NAND2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(KEYINPUT121), .B(n984), .ZN(n989) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(n987), .B(KEYINPUT57), .ZN(n988) );
  NAND2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1079 ( .A1(n995), .A2(n994), .ZN(n1022) );
  INV_X1 U1080 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1081 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n1002) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G22), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(G23), .B(G1976), .ZN(n996) );
  NOR2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1085 ( .A(G1986), .B(KEYINPUT124), .Z(n998) );
  XNOR2_X1 U1086 ( .A(G24), .B(n998), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1002), .B(n1001), .ZN(n1017) );
  XNOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(n1003), .B(G4), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(G6), .B(G1981), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1095 ( .A(KEYINPUT123), .B(G1956), .Z(n1008) );
  XNOR2_X1 U1096 ( .A(G20), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1011), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(G1966), .B(G21), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G1961), .B(G5), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1023), .B(KEYINPUT126), .ZN(n1024) );
  NOR2_X1 U1108 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XOR2_X1 U1109 ( .A(n1026), .B(KEYINPUT127), .Z(n1027) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .ZN(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
  INV_X1 U1112 ( .A(G303), .ZN(G166) );
endmodule

