

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  NOR2_X1 U321 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U322 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U323 ( .A(n345), .B(n344), .ZN(n346) );
  AND2_X1 U324 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U325 ( .A(n468), .B(KEYINPUT106), .ZN(n470) );
  XNOR2_X1 U326 ( .A(n343), .B(n342), .ZN(n462) );
  XNOR2_X1 U327 ( .A(n356), .B(n355), .ZN(n515) );
  XOR2_X1 U328 ( .A(G197GAT), .B(KEYINPUT89), .Z(n289) );
  NOR2_X1 U329 ( .A1(n478), .A2(n409), .ZN(n410) );
  INV_X1 U330 ( .A(KEYINPUT96), .ZN(n344) );
  INV_X1 U331 ( .A(KEYINPUT32), .ZN(n367) );
  XNOR2_X1 U332 ( .A(n335), .B(KEYINPUT22), .ZN(n336) );
  XNOR2_X1 U333 ( .A(n368), .B(n367), .ZN(n369) );
  INV_X1 U334 ( .A(n580), .ZN(n469) );
  XNOR2_X1 U335 ( .A(n337), .B(n336), .ZN(n341) );
  XNOR2_X1 U336 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U337 ( .A(n418), .B(n417), .ZN(n541) );
  NOR2_X1 U338 ( .A1(n441), .A2(n512), .ZN(n564) );
  NOR2_X1 U339 ( .A1(n510), .A2(n482), .ZN(n473) );
  INV_X1 U340 ( .A(G190GAT), .ZN(n445) );
  XNOR2_X1 U341 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U342 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U343 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n477), .B(n476), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G85GAT), .B(G92GAT), .Z(n366) );
  XOR2_X1 U346 ( .A(G106GAT), .B(G99GAT), .Z(n291) );
  XNOR2_X1 U347 ( .A(G162GAT), .B(G218GAT), .ZN(n290) );
  XNOR2_X1 U348 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U349 ( .A(n366), .B(n292), .Z(n294) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U352 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n296) );
  XNOR2_X1 U353 ( .A(KEYINPUT78), .B(G190GAT), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U355 ( .A(n298), .B(n297), .Z(n309) );
  XOR2_X1 U356 ( .A(G36GAT), .B(G43GAT), .Z(n300) );
  XNOR2_X1 U357 ( .A(G29GAT), .B(G50GAT), .ZN(n299) );
  XNOR2_X1 U358 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U359 ( .A(KEYINPUT71), .B(KEYINPUT7), .Z(n302) );
  XNOR2_X1 U360 ( .A(KEYINPUT8), .B(KEYINPUT70), .ZN(n301) );
  XNOR2_X1 U361 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U362 ( .A(n304), .B(n303), .Z(n384) );
  XOR2_X1 U363 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n306) );
  XNOR2_X1 U364 ( .A(G134GAT), .B(KEYINPUT65), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n384), .B(n307), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n478) );
  INV_X1 U368 ( .A(n478), .ZN(n552) );
  XOR2_X1 U369 ( .A(G169GAT), .B(KEYINPUT86), .Z(n311) );
  XNOR2_X1 U370 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U372 ( .A(n312), .B(KEYINPUT17), .Z(n314) );
  XNOR2_X1 U373 ( .A(G190GAT), .B(G176GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n354) );
  XOR2_X1 U375 ( .A(G113GAT), .B(KEYINPUT0), .Z(n316) );
  XNOR2_X1 U376 ( .A(G134GAT), .B(KEYINPUT84), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n423) );
  XOR2_X1 U378 ( .A(KEYINPUT20), .B(n423), .Z(n318) );
  NAND2_X1 U379 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U381 ( .A(KEYINPUT66), .B(KEYINPUT87), .Z(n320) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(KEYINPUT85), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U384 ( .A(n322), .B(n321), .ZN(n326) );
  XNOR2_X1 U385 ( .A(G127GAT), .B(G15GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n323), .B(G183GAT), .ZN(n403) );
  XNOR2_X1 U387 ( .A(G120GAT), .B(G99GAT), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n324), .B(G71GAT), .ZN(n362) );
  XOR2_X1 U389 ( .A(n403), .B(n362), .Z(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n354), .B(n327), .ZN(n525) );
  INV_X1 U392 ( .A(n525), .ZN(n518) );
  XOR2_X1 U393 ( .A(KEYINPUT2), .B(G162GAT), .Z(n329) );
  XNOR2_X1 U394 ( .A(KEYINPUT90), .B(G155GAT), .ZN(n328) );
  XNOR2_X1 U395 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U396 ( .A(KEYINPUT3), .B(n330), .Z(n424) );
  XOR2_X1 U397 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n332) );
  XNOR2_X1 U398 ( .A(G50GAT), .B(G211GAT), .ZN(n331) );
  XNOR2_X1 U399 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n424), .B(n333), .ZN(n343) );
  XNOR2_X1 U401 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n289), .B(n334), .ZN(n347) );
  XOR2_X1 U403 ( .A(G141GAT), .B(G22GAT), .Z(n374) );
  XOR2_X1 U404 ( .A(n347), .B(n374), .Z(n337) );
  NAND2_X1 U405 ( .A1(G228GAT), .A2(G233GAT), .ZN(n335) );
  XOR2_X1 U406 ( .A(G204GAT), .B(G78GAT), .Z(n339) );
  XNOR2_X1 U407 ( .A(G148GAT), .B(G106GAT), .ZN(n338) );
  XNOR2_X1 U408 ( .A(n339), .B(n338), .ZN(n363) );
  XOR2_X1 U409 ( .A(n363), .B(KEYINPUT24), .Z(n340) );
  XNOR2_X1 U410 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U411 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n420) );
  NAND2_X1 U412 ( .A1(G226GAT), .A2(G233GAT), .ZN(n345) );
  XOR2_X1 U413 ( .A(G211GAT), .B(G8GAT), .Z(n393) );
  XOR2_X1 U414 ( .A(n348), .B(n393), .Z(n350) );
  XNOR2_X1 U415 ( .A(G36GAT), .B(G92GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n356) );
  XOR2_X1 U417 ( .A(KEYINPUT97), .B(G204GAT), .Z(n352) );
  XNOR2_X1 U418 ( .A(G183GAT), .B(G64GAT), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U420 ( .A(n354), .B(n353), .Z(n355) );
  INV_X1 U421 ( .A(n515), .ZN(n449) );
  XOR2_X1 U422 ( .A(G64GAT), .B(KEYINPUT75), .Z(n358) );
  XNOR2_X1 U423 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n357) );
  XNOR2_X1 U424 ( .A(n358), .B(n357), .ZN(n402) );
  XOR2_X1 U425 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n360) );
  NAND2_X1 U426 ( .A1(G230GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U428 ( .A(n361), .B(KEYINPUT76), .Z(n365) );
  XNOR2_X1 U429 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n366), .B(G176GAT), .ZN(n368) );
  XOR2_X1 U432 ( .A(n402), .B(n371), .Z(n571) );
  XOR2_X1 U433 ( .A(n571), .B(KEYINPUT41), .Z(n529) );
  XOR2_X1 U434 ( .A(KEYINPUT29), .B(G197GAT), .Z(n373) );
  XNOR2_X1 U435 ( .A(G1GAT), .B(G169GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n375) );
  XOR2_X1 U437 ( .A(n375), .B(n374), .Z(n377) );
  XNOR2_X1 U438 ( .A(G113GAT), .B(G15GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n388) );
  XOR2_X1 U440 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n379) );
  NAND2_X1 U441 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U443 ( .A(n380), .B(KEYINPUT72), .Z(n386) );
  XOR2_X1 U444 ( .A(KEYINPUT68), .B(KEYINPUT73), .Z(n382) );
  XNOR2_X1 U445 ( .A(G8GAT), .B(KEYINPUT69), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U448 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U449 ( .A(n388), .B(n387), .Z(n545) );
  INV_X1 U450 ( .A(n545), .ZN(n566) );
  NAND2_X1 U451 ( .A1(n529), .A2(n566), .ZN(n389) );
  XNOR2_X1 U452 ( .A(KEYINPUT46), .B(n389), .ZN(n408) );
  XOR2_X1 U453 ( .A(G22GAT), .B(G78GAT), .Z(n391) );
  XNOR2_X1 U454 ( .A(G155GAT), .B(G71GAT), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U456 ( .A(n393), .B(n392), .Z(n395) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n407) );
  XOR2_X1 U459 ( .A(KEYINPUT80), .B(KEYINPUT83), .Z(n397) );
  XNOR2_X1 U460 ( .A(KEYINPUT15), .B(KEYINPUT81), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U462 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n399) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(KEYINPUT12), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U465 ( .A(n401), .B(n400), .Z(n405) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n576) );
  XNOR2_X1 U469 ( .A(n576), .B(KEYINPUT116), .ZN(n562) );
  NAND2_X1 U470 ( .A1(n408), .A2(n562), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n410), .B(KEYINPUT47), .ZN(n416) );
  XOR2_X1 U472 ( .A(KEYINPUT36), .B(n478), .Z(n580) );
  NOR2_X1 U473 ( .A1(n580), .A2(n576), .ZN(n411) );
  XOR2_X1 U474 ( .A(KEYINPUT45), .B(n411), .Z(n412) );
  NOR2_X1 U475 ( .A1(n571), .A2(n412), .ZN(n413) );
  XOR2_X1 U476 ( .A(KEYINPUT117), .B(n413), .Z(n414) );
  XNOR2_X1 U477 ( .A(n545), .B(KEYINPUT74), .ZN(n554) );
  NAND2_X1 U478 ( .A1(n414), .A2(n554), .ZN(n415) );
  NAND2_X1 U479 ( .A1(n416), .A2(n415), .ZN(n418) );
  XOR2_X1 U480 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n417) );
  NOR2_X1 U481 ( .A1(n449), .A2(n541), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n441) );
  XOR2_X1 U483 ( .A(KEYINPUT95), .B(G57GAT), .Z(n422) );
  XNOR2_X1 U484 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n422), .B(n421), .ZN(n428) );
  XOR2_X1 U486 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n426) );
  XNOR2_X1 U487 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U489 ( .A(n428), .B(n427), .ZN(n440) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n434) );
  XOR2_X1 U491 ( .A(G141GAT), .B(G148GAT), .Z(n430) );
  XNOR2_X1 U492 ( .A(G120GAT), .B(G127GAT), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U494 ( .A(G29GAT), .B(G85GAT), .Z(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U497 ( .A(KEYINPUT5), .B(G1GAT), .Z(n436) );
  XNOR2_X1 U498 ( .A(KEYINPUT94), .B(KEYINPUT92), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n512) );
  INV_X1 U502 ( .A(n564), .ZN(n442) );
  NOR2_X1 U503 ( .A1(n462), .A2(n442), .ZN(n443) );
  XOR2_X1 U504 ( .A(KEYINPUT55), .B(n443), .Z(n444) );
  NAND2_X1 U505 ( .A1(n518), .A2(n444), .ZN(n561) );
  NOR2_X1 U506 ( .A1(n552), .A2(n561), .ZN(n448) );
  XNOR2_X1 U507 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n446) );
  NOR2_X1 U508 ( .A1(n449), .A2(n525), .ZN(n450) );
  NOR2_X1 U509 ( .A1(n462), .A2(n450), .ZN(n451) );
  XOR2_X1 U510 ( .A(KEYINPUT25), .B(n451), .Z(n456) );
  NAND2_X1 U511 ( .A1(n462), .A2(n525), .ZN(n453) );
  INV_X1 U512 ( .A(KEYINPUT26), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n543) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(n515), .ZN(n460) );
  AND2_X1 U515 ( .A1(n543), .A2(n460), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n454), .B(KEYINPUT100), .ZN(n455) );
  NOR2_X1 U517 ( .A1(n456), .A2(n455), .ZN(n457) );
  XOR2_X1 U518 ( .A(KEYINPUT101), .B(n457), .Z(n458) );
  NOR2_X1 U519 ( .A1(n512), .A2(n458), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n459), .B(KEYINPUT102), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n460), .A2(n512), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT98), .ZN(n542) );
  XNOR2_X1 U523 ( .A(n462), .B(KEYINPUT28), .ZN(n522) );
  NOR2_X1 U524 ( .A1(n542), .A2(n522), .ZN(n527) );
  XNOR2_X1 U525 ( .A(n527), .B(KEYINPUT99), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n518), .B(KEYINPUT88), .ZN(n463) );
  NOR2_X1 U527 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U528 ( .A(KEYINPUT103), .B(n467), .ZN(n480) );
  AND2_X1 U529 ( .A1(n576), .A2(n480), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT37), .ZN(n510) );
  NOR2_X1 U531 ( .A1(n571), .A2(n554), .ZN(n472) );
  XNOR2_X1 U532 ( .A(KEYINPUT77), .B(n472), .ZN(n482) );
  XNOR2_X2 U533 ( .A(n473), .B(KEYINPUT38), .ZN(n496) );
  NAND2_X1 U534 ( .A1(n518), .A2(n496), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n475) );
  INV_X1 U536 ( .A(G43GAT), .ZN(n474) );
  NOR2_X1 U537 ( .A1(n478), .A2(n576), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT16), .ZN(n481) );
  NAND2_X1 U539 ( .A1(n481), .A2(n480), .ZN(n499) );
  NOR2_X1 U540 ( .A1(n482), .A2(n499), .ZN(n489) );
  NAND2_X1 U541 ( .A1(n489), .A2(n512), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n483), .B(KEYINPUT34), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U544 ( .A1(n515), .A2(n489), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n485), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U547 ( .A1(n489), .A2(n518), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  XOR2_X1 U550 ( .A(G22GAT), .B(KEYINPUT105), .Z(n491) );
  NAND2_X1 U551 ( .A1(n489), .A2(n522), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT107), .B(n492), .ZN(n494) );
  NAND2_X1 U555 ( .A1(n496), .A2(n512), .ZN(n493) );
  XOR2_X1 U556 ( .A(n494), .B(n493), .Z(G1328GAT) );
  NAND2_X1 U557 ( .A1(n496), .A2(n515), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n496), .A2(n522), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U561 ( .A(G57GAT), .B(KEYINPUT109), .Z(n501) );
  NAND2_X1 U562 ( .A1(n545), .A2(n529), .ZN(n498) );
  XNOR2_X1 U563 ( .A(KEYINPUT110), .B(n498), .ZN(n511) );
  NOR2_X1 U564 ( .A1(n511), .A2(n499), .ZN(n507) );
  NAND2_X1 U565 ( .A1(n507), .A2(n512), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n501), .B(n500), .ZN(n503) );
  XOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT111), .Z(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n515), .A2(n507), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n507), .A2(n518), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(KEYINPUT112), .ZN(n506) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U575 ( .A1(n507), .A2(n522), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT113), .Z(n514) );
  NOR2_X1 U578 ( .A1(n511), .A2(n510), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n521), .A2(n512), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n515), .A2(n521), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n516), .B(KEYINPUT114), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(n517), .ZN(G1337GAT) );
  XOR2_X1 U584 ( .A(G99GAT), .B(KEYINPUT115), .Z(n520) );
  NAND2_X1 U585 ( .A1(n521), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n541), .A2(n525), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n536) );
  NOR2_X1 U592 ( .A1(n554), .A2(n536), .ZN(n528) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n528), .Z(G1340GAT) );
  INV_X1 U594 ( .A(n529), .ZN(n556) );
  NOR2_X1 U595 ( .A1(n556), .A2(n536), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n533) );
  XNOR2_X1 U599 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n562), .A2(n536), .ZN(n534) );
  XOR2_X1 U602 ( .A(n535), .B(n534), .Z(G1342GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n552), .ZN(n540) );
  XOR2_X1 U604 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n538) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT120), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n544) );
  BUF_X1 U609 ( .A(n543), .Z(n565) );
  NAND2_X1 U610 ( .A1(n544), .A2(n565), .ZN(n551) );
  NOR2_X1 U611 ( .A1(n545), .A2(n551), .ZN(n546) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n556), .A2(n551), .ZN(n548) );
  XNOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n576), .A2(n551), .ZN(n550) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n561), .ZN(n555) );
  XOR2_X1 U622 ( .A(G169GAT), .B(n555), .Z(G1348GAT) );
  NOR2_X1 U623 ( .A1(n561), .A2(n556), .ZN(n560) );
  XOR2_X1 U624 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n558) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n563), .Z(G1350GAT) );
  XOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .Z(n568) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n579) );
  INV_X1 U632 ( .A(n579), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n572), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n574) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .Z(n578) );
  OR2_X1 U642 ( .A1(n579), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

