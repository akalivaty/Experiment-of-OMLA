//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n450, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n602, new_n603, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  INV_X1    g024(.A(G2106), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  AND2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR3_X1    g033(.A1(new_n455), .A2(KEYINPUT67), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT67), .B1(new_n455), .B2(new_n458), .ZN(new_n460));
  OAI211_X1 g035(.A(new_n459), .B(new_n460), .C1(new_n454), .C2(new_n450), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(new_n468), .A3(G137), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT3), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n473), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n467), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n472), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NOR2_X1   g059(.A1(new_n478), .A2(new_n467), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n467), .C2(G112), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n478), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n467), .A2(new_n468), .A3(G138), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT70), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n467), .A2(new_n468), .A3(G138), .A4(new_n494), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n463), .A2(G102), .A3(G2104), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n468), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(new_n463), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n498), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT71), .A3(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OR2_X1    g094(.A1(new_n511), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT72), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n508), .A2(G63), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n517), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n515), .A2(new_n531), .B1(new_n517), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT73), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n508), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(new_n510), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT74), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n534), .A2(new_n539), .A3(new_n536), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n515), .A2(new_n544), .B1(new_n517), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT76), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n550), .A2(new_n554), .ZN(G188));
  AOI22_X1  g130(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n556), .A2(new_n510), .ZN(new_n557));
  INV_X1    g132(.A(new_n515), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G91), .ZN(new_n559));
  OAI211_X1 g134(.A(G53), .B(G543), .C1(new_n512), .C2(new_n513), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  OR2_X1    g138(.A1(new_n508), .A2(G74), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n514), .A2(G543), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(G651), .B1(G49), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n515), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n558), .A2(KEYINPUT77), .A3(G87), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n566), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n510), .B1(new_n573), .B2(new_n517), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n508), .A2(G86), .A3(new_n514), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n510), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n515), .A2(new_n581), .B1(new_n517), .B2(new_n582), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n580), .A2(new_n583), .ZN(G290));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OR3_X1    g160(.A1(new_n515), .A2(KEYINPUT10), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g161(.A(KEYINPUT10), .B1(new_n515), .B2(new_n585), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT79), .B(G66), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n508), .A2(new_n589), .B1(G79), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G54), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n510), .B1(new_n591), .B2(new_n517), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(G171), .B2(new_n595), .ZN(G284));
  OAI21_X1  g172(.A(new_n596), .B1(G171), .B2(new_n595), .ZN(G321));
  NAND2_X1  g173(.A1(G299), .A2(new_n595), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G168), .B2(new_n595), .ZN(G297));
  OAI21_X1  g175(.A(new_n599), .B1(G168), .B2(new_n595), .ZN(G280));
  NOR2_X1   g176(.A1(new_n594), .A2(G559), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(G860), .B2(new_n593), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT80), .Z(G148));
  INV_X1    g179(.A(new_n547), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(new_n595), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n602), .B2(new_n595), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n463), .A2(G2104), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n478), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n610), .B(new_n611), .Z(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(G2100), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n612), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n485), .A2(G123), .ZN(new_n616));
  OAI221_X1 g191(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n467), .C2(G111), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n488), .A2(G135), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT83), .Z(new_n620));
  AND2_X1   g195(.A1(new_n620), .A2(G2096), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n620), .A2(G2096), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT84), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2435), .ZN(new_n626));
  XOR2_X1   g201(.A(G2427), .B(G2438), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT14), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G1341), .B(G1348), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n634), .B(new_n635), .Z(new_n636));
  AND2_X1   g211(.A1(new_n636), .A2(G14), .ZN(G401));
  XNOR2_X1  g212(.A(G2072), .B(G2078), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2100), .Z(new_n645));
  INV_X1    g220(.A(new_n641), .ZN(new_n646));
  OAI21_X1  g221(.A(KEYINPUT17), .B1(new_n646), .B2(new_n639), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n643), .B1(new_n647), .B2(new_n642), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT86), .B(G2096), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(new_n650), .ZN(G227));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n662), .B(new_n663), .C1(new_n661), .C2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(G1981), .B(G1986), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(G229));
  INV_X1    g246(.A(G16), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n672), .A2(G22), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(G303), .B2(G16), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(G1971), .ZN(new_n675));
  NAND4_X1  g250(.A1(new_n566), .A2(G16), .A3(new_n569), .A4(new_n570), .ZN(new_n676));
  OR2_X1    g251(.A1(G16), .A2(G23), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT33), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(G305), .A2(G16), .ZN(new_n681));
  INV_X1    g256(.A(G6), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(G16), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT32), .B(G1981), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n681), .B(new_n684), .C1(new_n682), .C2(G16), .ZN(new_n687));
  NAND4_X1  g262(.A1(new_n675), .A2(new_n680), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n485), .A2(G119), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n488), .A2(new_n692), .A3(G131), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n463), .ZN(new_n694));
  INV_X1    g269(.A(G131), .ZN(new_n695));
  OAI21_X1  g270(.A(KEYINPUT88), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI221_X1 g271(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n467), .C2(G107), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n691), .A2(new_n693), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT89), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT89), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n690), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n690), .A2(G25), .ZN(new_n702));
  OR3_X1    g277(.A1(new_n701), .A2(KEYINPUT90), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT35), .B(G1991), .ZN(new_n704));
  OAI21_X1  g279(.A(KEYINPUT90), .B1(new_n701), .B2(new_n702), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n672), .A2(G24), .ZN(new_n711));
  INV_X1    g286(.A(G290), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n672), .ZN(new_n713));
  INV_X1    g288(.A(G1986), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND4_X1  g290(.A1(new_n689), .A2(new_n709), .A3(new_n710), .A4(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n688), .B2(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n703), .A2(new_n705), .ZN(new_n718));
  INV_X1    g293(.A(new_n704), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(new_n706), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT91), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n716), .A2(new_n722), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n690), .A2(G33), .ZN(new_n728));
  NAND2_X1  g303(.A1(G115), .A2(G2104), .ZN(new_n729));
  INV_X1    g304(.A(G127), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n478), .B2(new_n730), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n731), .A2(new_n481), .B1(new_n488), .B2(G139), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(KEYINPUT25), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n733), .A2(KEYINPUT25), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT95), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n728), .B1(new_n737), .B2(new_n690), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2072), .Z(new_n739));
  NAND3_X1  g314(.A1(new_n672), .A2(KEYINPUT23), .A3(G20), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT23), .ZN(new_n741));
  INV_X1    g316(.A(G20), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(G299), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n740), .B(new_n743), .C1(new_n744), .C2(new_n672), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G1956), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n690), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n485), .A2(G128), .ZN(new_n749));
  OAI221_X1 g324(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n467), .C2(G116), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n488), .A2(G140), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G29), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(KEYINPUT94), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n748), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n758), .A2(new_n759), .B1(G1956), .B2(new_n745), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n672), .A2(G5), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n761), .B(new_n762), .C1(G171), .C2(new_n672), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n739), .A2(new_n746), .A3(new_n760), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n690), .A2(G27), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G164), .B2(new_n690), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n765), .B(new_n766), .S(KEYINPUT100), .Z(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(G2078), .Z(new_n768));
  OR2_X1    g343(.A1(G29), .A2(G32), .ZN(new_n769));
  AOI22_X1  g344(.A1(G129), .A2(new_n485), .B1(new_n488), .B2(G141), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT26), .Z(new_n772));
  INV_X1    g347(.A(G105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n772), .C1(new_n773), .C2(new_n609), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n769), .B1(new_n774), .B2(new_n690), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n619), .A2(new_n690), .ZN(new_n778));
  INV_X1    g353(.A(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT93), .B1(new_n779), .B2(G16), .ZN(new_n780));
  OR3_X1    g355(.A1(new_n779), .A2(KEYINPUT93), .A3(G16), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n780), .B(new_n781), .C1(new_n547), .C2(new_n672), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1341), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n690), .B2(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n768), .A2(new_n777), .A3(new_n778), .A4(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT96), .B(G34), .Z(new_n787));
  INV_X1    g362(.A(KEYINPUT24), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n789), .A2(new_n690), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n793), .B(new_n794), .C1(new_n690), .C2(new_n483), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT98), .Z(new_n798));
  AOI22_X1  g373(.A1(new_n795), .A2(new_n796), .B1(new_n775), .B2(new_n776), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n690), .A2(G35), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G162), .B2(new_n690), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT29), .B(G2090), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n798), .A2(new_n799), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n672), .A2(G4), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n593), .B2(new_n672), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1348), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n764), .A2(new_n786), .A3(new_n804), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n727), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT31), .B(G11), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n716), .A2(new_n722), .A3(new_n726), .ZN(new_n811));
  INV_X1    g386(.A(new_n725), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n723), .A2(new_n724), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g389(.A1(new_n809), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n816));
  NAND2_X1  g391(.A1(G168), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G16), .B2(G21), .ZN(new_n818));
  INV_X1    g393(.A(G1966), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n762), .B1(G171), .B2(new_n672), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G1961), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT99), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n815), .A2(new_n816), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n809), .A2(new_n824), .A3(new_n810), .A4(new_n814), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT101), .B1(new_n826), .B2(new_n820), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n815), .A2(new_n829), .A3(new_n821), .A4(new_n824), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT102), .B1(new_n826), .B2(new_n820), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(G150));
  XNOR2_X1  g407(.A(KEYINPUT103), .B(G93), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n515), .A2(new_n833), .B1(new_n517), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n508), .A2(G67), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n510), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G860), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT37), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n605), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n547), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n593), .A2(G559), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n847), .B(new_n848), .Z(new_n849));
  OAI21_X1  g424(.A(new_n842), .B1(new_n849), .B2(G860), .ZN(G145));
  NAND2_X1  g425(.A1(new_n737), .A2(new_n752), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n737), .A2(new_n752), .ZN(new_n853));
  NAND2_X1  g428(.A1(G114), .A2(G2104), .ZN(new_n854));
  INV_X1    g429(.A(G126), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n478), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G2105), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n857), .A2(new_n496), .A3(new_n499), .A4(new_n497), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n774), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n852), .A2(new_n853), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n737), .A2(new_n752), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n862), .B2(new_n851), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT106), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n860), .B1(new_n852), .B2(new_n853), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n862), .A2(new_n851), .A3(new_n859), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n699), .A2(new_n700), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n485), .A2(G130), .ZN(new_n872));
  OAI221_X1 g447(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n467), .C2(G118), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n488), .A2(G142), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n871), .A2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  INV_X1    g455(.A(new_n870), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n612), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n882), .A3(new_n612), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT107), .B1(new_n869), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n861), .A2(new_n863), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n483), .B(new_n619), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n490), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n864), .A2(new_n868), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n886), .A4(new_n885), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n888), .A2(new_n890), .A3(new_n893), .A4(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n887), .A2(new_n889), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n887), .A2(new_n889), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT108), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n897), .A2(new_n901), .A3(new_n904), .A4(new_n898), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT40), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(G395));
  XNOR2_X1  g483(.A(G288), .B(KEYINPUT110), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n712), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n910), .A2(KEYINPUT111), .ZN(new_n911));
  XNOR2_X1  g486(.A(G305), .B(G303), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(KEYINPUT111), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT42), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n845), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(new_n602), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n593), .B(new_n744), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(KEYINPUT109), .B(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(KEYINPUT41), .B2(new_n921), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n922), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n918), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n840), .A2(new_n595), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G295));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n930), .ZN(G331));
  XNOR2_X1  g507(.A(G171), .B(G286), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n919), .ZN(new_n934));
  XNOR2_X1  g509(.A(G171), .B(G168), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n845), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n934), .A2(new_n936), .A3(new_n925), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n921), .B1(new_n934), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n913), .A2(new_n915), .ZN(new_n940));
  AOI21_X1  g515(.A(G37), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n916), .B1(new_n938), .B2(new_n937), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT43), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n921), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(KEYINPUT41), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n944), .B2(new_n923), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n946), .A2(new_n934), .A3(new_n936), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n916), .B1(new_n938), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n934), .A2(new_n936), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n944), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n934), .A2(new_n936), .A3(new_n925), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n915), .A3(new_n913), .A4(new_n951), .ZN(new_n952));
  AND4_X1   g527(.A1(KEYINPUT43), .A2(new_n948), .A3(new_n952), .A4(new_n898), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT44), .B1(new_n943), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n941), .B2(new_n942), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n955), .A2(new_n948), .A3(new_n952), .A4(new_n898), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n954), .B1(new_n958), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g534(.A(KEYINPUT126), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n498), .B2(new_n501), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT112), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n858), .A2(KEYINPUT112), .A3(new_n961), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n964), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n472), .A2(G40), .A3(new_n482), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n969), .A2(KEYINPUT113), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(KEYINPUT113), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n752), .B(G2067), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT114), .ZN(new_n974));
  INV_X1    g549(.A(G1996), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n774), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n699), .A2(new_n700), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n719), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n719), .B2(new_n978), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(G1986), .B2(G290), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n972), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n575), .A2(new_n577), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n576), .ZN(new_n987));
  OAI21_X1  g562(.A(G1981), .B1(new_n574), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(KEYINPUT49), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g567(.A(KEYINPUT115), .B(G8), .Z(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n963), .B2(new_n968), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n986), .B(new_n988), .C1(new_n990), .C2(KEYINPUT49), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G288), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G1976), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n995), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT52), .ZN(new_n1001));
  INV_X1    g576(.A(G1976), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(new_n995), .A3(new_n1003), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n997), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G303), .A2(G8), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT55), .Z(new_n1007));
  NAND2_X1  g582(.A1(new_n962), .A2(KEYINPUT50), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n858), .A2(new_n1009), .A3(new_n961), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1008), .A2(new_n968), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G2090), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n962), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n858), .A2(KEYINPUT45), .A3(new_n961), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n968), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G1971), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1007), .A2(new_n1020), .A3(G8), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1005), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1007), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1013), .A2(KEYINPUT117), .A3(new_n1019), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n993), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1022), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT62), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1008), .A2(new_n796), .A3(new_n968), .A4(new_n1010), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1017), .A2(new_n819), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n967), .B1(new_n962), .B2(KEYINPUT50), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(KEYINPUT118), .A3(new_n796), .A4(new_n1010), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G286), .A2(new_n993), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT51), .B1(G286), .B2(new_n993), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n993), .B2(new_n1036), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1029), .B(new_n1039), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1017), .A2(G2078), .ZN(new_n1047));
  OAI22_X1  g622(.A1(new_n1047), .A2(KEYINPUT53), .B1(G1961), .B2(new_n1011), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(KEYINPUT53), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1036), .A2(new_n993), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n1043), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1038), .B1(new_n1036), .B2(G8), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1054), .B1(new_n1055), .B2(new_n1040), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1029), .B1(new_n1056), .B2(new_n1039), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1052), .A2(new_n1057), .A3(G301), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n962), .A2(new_n967), .A3(G2067), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1034), .A2(new_n1010), .ZN(new_n1060));
  INV_X1    g635(.A(G1348), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1059), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n594), .B1(new_n1062), .B2(KEYINPUT60), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1348), .B1(new_n1034), .B2(new_n1010), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n1065));
  NOR4_X1   g640(.A1(new_n1064), .A2(new_n1065), .A3(new_n593), .A4(new_n1059), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1063), .A2(new_n1066), .B1(KEYINPUT60), .B2(new_n1062), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1060), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n1070));
  XNOR2_X1  g645(.A(G299), .B(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT56), .B(G2072), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1015), .A2(new_n968), .A3(new_n1016), .A4(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT61), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1069), .A2(new_n1071), .A3(KEYINPUT61), .A4(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1015), .A2(new_n975), .A3(new_n968), .A4(new_n1016), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n962), .B2(new_n967), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n547), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(KEYINPUT120), .A3(new_n547), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT120), .B1(new_n1082), .B2(new_n547), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1084), .B(new_n605), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1092));
  OAI22_X1  g667(.A1(new_n1091), .A2(new_n1092), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1067), .A2(new_n1078), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  AND2_X1   g669(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(new_n1071), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1074), .B(new_n593), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1056), .A2(new_n1039), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G171), .B(KEYINPUT54), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n472), .A2(KEYINPUT122), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n482), .B(G40), .C1(new_n471), .C2(new_n1103), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1102), .A2(new_n1104), .A3(KEYINPUT123), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT123), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(KEYINPUT53), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1016), .ZN(new_n1108));
  NOR4_X1   g683(.A1(new_n966), .A2(new_n1107), .A3(G2078), .A4(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1101), .B1(new_n1048), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n1111));
  XNOR2_X1  g686(.A(G171), .B(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1099), .A2(new_n1100), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1028), .B1(new_n1058), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n997), .A2(new_n1002), .A3(new_n998), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n986), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n995), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1020), .A2(G8), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1005), .A2(new_n1120), .A3(new_n1007), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1053), .A2(G286), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1028), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT63), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT63), .B1(new_n1120), .B2(new_n1007), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1123), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n1022), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1122), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n984), .B1(new_n1116), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n972), .B2(new_n983), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n970), .A2(new_n1134), .A3(new_n971), .A4(new_n982), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT48), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n972), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n980), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1133), .A2(KEYINPUT48), .A3(new_n1135), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT46), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n972), .B2(G1996), .ZN(new_n1144));
  INV_X1    g719(.A(new_n974), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n970), .B(new_n971), .C1(new_n774), .C2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n970), .A2(KEYINPUT46), .A3(new_n975), .A4(new_n971), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT124), .B(KEYINPUT47), .Z(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1149), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n978), .A2(new_n719), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n977), .A2(new_n1154), .B1(G2067), .B2(new_n752), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1139), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1142), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n960), .B1(new_n1132), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1142), .A2(new_n1153), .A3(new_n1156), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT63), .B1(new_n1028), .B2(new_n1123), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1121), .B(new_n1119), .C1(new_n1160), .C2(new_n1129), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1099), .A2(new_n1100), .A3(new_n1114), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1100), .A2(KEYINPUT62), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(G171), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1162), .B1(new_n1164), .B2(new_n1052), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1161), .B1(new_n1028), .B2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(KEYINPUT126), .B(new_n1159), .C1(new_n1166), .C2(new_n984), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1158), .A2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g743(.A1(G401), .A2(G229), .ZN(new_n1170));
  OAI21_X1  g744(.A(new_n1170), .B1(new_n956), .B2(new_n957), .ZN(new_n1171));
  INV_X1    g745(.A(G319), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1172), .A2(G227), .ZN(new_n1173));
  XOR2_X1   g747(.A(new_n1173), .B(KEYINPUT127), .Z(new_n1174));
  NAND2_X1  g748(.A1(new_n902), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1171), .A2(new_n1175), .ZN(G308));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n1177), .B(new_n1170), .C1(new_n956), .C2(new_n957), .ZN(G225));
endmodule


