//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n462), .A2(new_n463), .A3(G137), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT69), .ZN(G160));
  XNOR2_X1  g050(.A(KEYINPUT68), .B(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n463), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n463), .A2(new_n465), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI22_X1  g055(.A1(G124), .A2(new_n478), .B1(new_n480), .B2(G136), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT70), .ZN(G162));
  NAND2_X1  g059(.A1(G126), .A2(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n465), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT71), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n485), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n469), .B2(new_n470), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G138), .B1(new_n469), .B2(new_n470), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n500), .B2(new_n476), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n462), .A2(new_n463), .A3(new_n502), .A4(G138), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n492), .A2(new_n499), .B1(new_n501), .B2(new_n503), .ZN(G164));
  NAND2_X1  g079(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n512), .A2(new_n518), .ZN(G166));
  INV_X1    g094(.A(new_n514), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n522), .B(new_n524), .C1(new_n516), .C2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n521), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n511), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n514), .A2(new_n530), .B1(new_n516), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND2_X1  g109(.A1(new_n509), .A2(G56), .ZN(new_n535));
  INV_X1    g110(.A(G68), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n536), .B2(new_n506), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n511), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n538), .B2(new_n537), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n513), .A2(G543), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n520), .A2(G81), .B1(new_n541), .B2(G43), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  NAND2_X1  g124(.A1(new_n541), .A2(G53), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n541), .A2(new_n552), .A3(G53), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(KEYINPUT9), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  INV_X1    g130(.A(new_n550), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n509), .B(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G651), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n551), .A2(new_n555), .A3(KEYINPUT9), .A4(new_n553), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n520), .A2(G91), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n559), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n520), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n541), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n520), .A2(G86), .B1(new_n541), .B2(G48), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n511), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n511), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n514), .A2(new_n581), .B1(new_n516), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(G66), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n562), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT77), .Z(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G92), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n514), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n592), .A2(new_n595), .B1(G54), .B2(new_n541), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n586), .B1(new_n598), .B2(G868), .ZN(G284));
  XOR2_X1   g174(.A(G284), .B(KEYINPUT78), .Z(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G299), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G297));
  OAI21_X1  g178(.A(new_n602), .B1(new_n601), .B2(G168), .ZN(G280));
  XNOR2_X1  g179(.A(KEYINPUT79), .B(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(G860), .B2(new_n605), .ZN(G148));
  NAND2_X1  g181(.A1(new_n543), .A2(new_n601), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n605), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n601), .ZN(G323));
  XOR2_X1   g185(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n611));
  XNOR2_X1  g186(.A(G323), .B(new_n611), .ZN(G282));
  AOI22_X1  g187(.A1(G123), .A2(new_n478), .B1(new_n480), .B2(G135), .ZN(new_n613));
  OAI221_X1 g188(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT82), .Z(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(G2096), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n463), .A2(new_n466), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT13), .B(G2100), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n617), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT83), .Z(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2443), .B(G2446), .Z(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(G14), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n636), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT85), .Z(new_n645));
  NOR2_X1   g220(.A1(G2072), .A2(G2078), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n442), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(KEYINPUT17), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n643), .B(new_n644), .C1(new_n442), .C2(new_n646), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n645), .A2(new_n649), .A3(new_n643), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n658), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G1981), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G1986), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1991), .B(G1996), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT87), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(G229));
  NOR2_X1   g253(.A1(KEYINPUT94), .A2(G2072), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT25), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n480), .A2(G139), .ZN(new_n683));
  AOI22_X1  g258(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n682), .B(new_n683), .C1(new_n462), .C2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT93), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G29), .ZN(new_n687));
  INV_X1    g262(.A(G29), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(G33), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n679), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(KEYINPUT94), .A2(G2072), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(G32), .ZN(new_n693));
  NAND3_X1  g268(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT26), .Z(new_n695));
  INV_X1    g270(.A(G129), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n477), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n466), .A2(G105), .ZN(new_n698));
  INV_X1    g273(.A(G141), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n479), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n693), .B1(new_n702), .B2(new_n688), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT27), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT95), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n703), .B(new_n705), .Z(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G5), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G171), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1961), .ZN(new_n710));
  INV_X1    g285(.A(G28), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT30), .ZN(new_n712));
  AOI21_X1  g287(.A(G29), .B1(new_n711), .B2(KEYINPUT30), .ZN(new_n713));
  OR2_X1    g288(.A1(KEYINPUT31), .A2(G11), .ZN(new_n714));
  NAND2_X1  g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n616), .B2(new_n688), .ZN(new_n717));
  NAND2_X1  g292(.A1(G160), .A2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(G29), .B1(new_n719), .B2(KEYINPUT24), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(KEYINPUT24), .B2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR4_X1   g299(.A1(new_n706), .A2(new_n710), .A3(new_n717), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n722), .A2(new_n723), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT96), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n707), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n707), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1966), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n688), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n688), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2078), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n692), .A2(new_n725), .A3(new_n727), .A4(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT97), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G35), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G162), .B2(G29), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT29), .B(G2090), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n688), .A2(G26), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT92), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n478), .A2(G128), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n480), .A2(G140), .ZN(new_n746));
  OAI221_X1 g321(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n744), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2067), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n739), .A2(new_n740), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n741), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n707), .A2(G20), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G299), .B2(G16), .ZN(new_n756));
  INV_X1    g331(.A(G1956), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n707), .A2(G19), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n544), .B2(new_n707), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1341), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT91), .Z(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n597), .B2(new_n707), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(G1348), .Z(new_n765));
  NOR4_X1   g340(.A1(new_n752), .A2(new_n758), .A3(new_n761), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n736), .A2(new_n737), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT99), .ZN(new_n768));
  MUX2_X1   g343(.A(G6), .B(G305), .S(G16), .Z(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT32), .B(G1981), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G23), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT90), .Z(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G288), .B2(new_n707), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n707), .A2(G22), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G166), .B2(new_n707), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1971), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n771), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT34), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n707), .A2(G24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n584), .B2(new_n707), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1986), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n688), .A2(G25), .ZN(new_n787));
  AOI22_X1  g362(.A1(G119), .A2(new_n478), .B1(new_n480), .B2(G131), .ZN(new_n788));
  OAI221_X1 g363(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n462), .C2(G107), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n787), .B1(new_n791), .B2(new_n688), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT35), .B(G1991), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT88), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n786), .B1(new_n795), .B2(KEYINPUT89), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(KEYINPUT89), .B2(new_n795), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n782), .A2(new_n783), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT36), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n768), .A2(new_n799), .ZN(G150));
  INV_X1    g375(.A(G150), .ZN(G311));
  INV_X1    g376(.A(G860), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT39), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n598), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(new_n511), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n520), .A2(G93), .B1(new_n541), .B2(G55), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT100), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n544), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n807), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(new_n543), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n805), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(new_n803), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT101), .B1(new_n814), .B2(new_n803), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n802), .B1(new_n803), .B2(new_n814), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT102), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n811), .A2(G860), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(new_n686), .B(new_n702), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n495), .A2(new_n497), .ZN(new_n825));
  AOI211_X1 g400(.A(KEYINPUT103), .B(new_n825), .C1(new_n501), .C2(new_n503), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT103), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n501), .A2(new_n503), .ZN(new_n828));
  INV_X1    g403(.A(new_n825), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n748), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n824), .B(new_n832), .ZN(new_n833));
  AOI22_X1  g408(.A1(G130), .A2(new_n478), .B1(new_n480), .B2(G142), .ZN(new_n834));
  OAI221_X1 g409(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n462), .C2(G118), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n790), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n621), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(KEYINPUT104), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(KEYINPUT104), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n616), .B(G160), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G162), .Z(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n843), .A2(new_n845), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g425(.A(KEYINPUT110), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n584), .B(G288), .Z(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(KEYINPUT109), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(G303), .B(G305), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(KEYINPUT109), .B2(new_n852), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n852), .A2(KEYINPUT109), .ZN(new_n858));
  INV_X1    g433(.A(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n860), .A2(new_n853), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n851), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n853), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n854), .A2(new_n856), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT110), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT42), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n864), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(KEYINPUT42), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n813), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n609), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n874));
  NAND2_X1  g449(.A1(G299), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n566), .A2(new_n567), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n876), .A2(KEYINPUT106), .A3(new_n565), .A4(new_n559), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n598), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(G299), .A2(new_n874), .A3(new_n597), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n873), .B1(new_n880), .B2(KEYINPUT41), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n878), .A2(KEYINPUT107), .A3(new_n882), .A4(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n880), .A2(KEYINPUT41), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(KEYINPUT108), .A3(KEYINPUT41), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n872), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n871), .B(new_n608), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n880), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n869), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n869), .B1(new_n890), .B2(new_n892), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT111), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n869), .A2(new_n890), .A3(KEYINPUT111), .A4(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(G868), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n811), .A2(new_n601), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(G295));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n900), .ZN(G331));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n810), .A2(G301), .A3(new_n812), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G301), .B1(new_n810), .B2(new_n812), .ZN(new_n906));
  OAI21_X1  g481(.A(G286), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(G168), .A3(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n889), .B2(new_n884), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n880), .B1(new_n907), .B2(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n866), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n915));
  INV_X1    g490(.A(new_n910), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n866), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n913), .A2(new_n914), .A3(new_n919), .A4(new_n847), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n880), .B(KEYINPUT41), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n912), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n847), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  AOI211_X1 g498(.A(new_n866), .B(new_n912), .C1(new_n915), .C2(new_n916), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT43), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n903), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT43), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n913), .A2(new_n847), .A3(new_n919), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(KEYINPUT43), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n926), .B1(new_n929), .B2(new_n903), .ZN(G397));
  INV_X1    g505(.A(G138), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n486), .B2(new_n487), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n502), .B1(new_n932), .B2(new_n462), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n500), .A2(new_n476), .A3(KEYINPUT4), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n829), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT103), .ZN(new_n936));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n825), .B1(new_n501), .B2(new_n503), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n827), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(G40), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n468), .A2(new_n943), .A3(new_n473), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1996), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT46), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n748), .B(G2067), .Z(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n702), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n948), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n951), .A2(KEYINPUT126), .A3(new_n954), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(KEYINPUT47), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G290), .A2(G1986), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n948), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n701), .B(new_n949), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n952), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n790), .B(new_n794), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n961), .A2(new_n962), .B1(new_n948), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n791), .A2(new_n794), .ZN(new_n970));
  OAI22_X1  g545(.A1(new_n965), .A2(new_n970), .B1(G2067), .B2(new_n748), .ZN(new_n971));
  AOI22_X1  g546(.A1(new_n963), .A2(new_n969), .B1(new_n948), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n959), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT47), .B1(new_n957), .B2(new_n958), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT125), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT54), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n828), .B2(new_n829), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n981), .A3(new_n944), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(G1961), .ZN(new_n984));
  INV_X1    g559(.A(G2078), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n492), .A2(new_n499), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n828), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n937), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n945), .B1(new_n988), .B2(new_n941), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n941), .A2(G1384), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n831), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n936), .A2(new_n990), .A3(new_n939), .A4(new_n991), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n985), .B(new_n989), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n984), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(KEYINPUT53), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n936), .A2(new_n939), .A3(new_n991), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n1000), .B2(new_n993), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1002), .B1(new_n942), .B2(new_n944), .ZN(new_n1003));
  AOI211_X1 g578(.A(KEYINPUT122), .B(new_n945), .C1(new_n940), .C2(new_n941), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n997), .A2(G301), .A3(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n941), .B1(new_n938), .B2(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n944), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT116), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(new_n944), .C1(new_n979), .C2(KEYINPUT45), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n987), .A2(new_n1012), .A3(new_n991), .ZN(new_n1013));
  INV_X1    g588(.A(new_n991), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT117), .B1(G164), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1009), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(new_n998), .ZN(new_n1018));
  AOI21_X1  g593(.A(G301), .B1(new_n997), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n977), .B1(new_n1006), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1966), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1012), .B1(new_n987), .B2(new_n991), .ZN(new_n1022));
  NOR3_X1   g597(.A1(G164), .A2(KEYINPUT117), .A3(new_n1014), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1011), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1010), .B1(new_n1007), .B2(new_n944), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND4_X1   g601(.A1(new_n723), .A2(new_n978), .A3(new_n981), .A4(new_n944), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(G168), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1027), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(G168), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n1031), .B2(G168), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  OR2_X1    g613(.A1(new_n982), .A2(G2090), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G164), .A2(G1384), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n944), .B1(new_n1040), .B2(KEYINPUT45), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1000), .B2(new_n993), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1039), .B1(new_n1042), .B2(G1971), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT114), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G166), .A2(new_n1034), .ZN(new_n1045));
  XOR2_X1   g620(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1045), .B1(KEYINPUT115), .B2(KEYINPUT55), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1039), .B(new_n1050), .C1(new_n1042), .C2(G1971), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1044), .A2(G8), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n979), .A2(new_n944), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G305), .A2(G1981), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n575), .A2(new_n577), .A3(new_n668), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1054), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1054), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1061), .B(new_n1063), .C1(new_n1062), .C2(G288), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G288), .A2(new_n1062), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT52), .B1(new_n1054), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1060), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n945), .B1(new_n1040), .B2(new_n980), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n980), .B2(new_n979), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1042), .A2(G1971), .B1(G2090), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1049), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1067), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1020), .A2(new_n1038), .A3(new_n1052), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n997), .A2(new_n1018), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT54), .B1(new_n1075), .B2(G171), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n997), .A2(new_n1077), .A3(new_n1005), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n997), .A2(new_n1005), .ZN(new_n1079));
  AOI21_X1  g654(.A(G301), .B1(new_n1079), .B2(KEYINPUT123), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT124), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G286), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1036), .B1(new_n1035), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1030), .A2(KEYINPUT51), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1052), .B(new_n1073), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1080), .A2(new_n1078), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1076), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .A4(new_n1020), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1042), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1069), .A2(new_n757), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1097), .A2(KEYINPUT119), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n1099));
  XNOR2_X1  g674(.A(G299), .B(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n1097), .B2(KEYINPUT119), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1101), .ZN(new_n1102));
  OAI22_X1  g677(.A1(new_n983), .A2(G1348), .B1(G2067), .B2(new_n1053), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n598), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1100), .A2(new_n1096), .A3(new_n1095), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT58), .B(G1341), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n979), .B2(new_n944), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT120), .B(G1996), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1110), .B1(new_n1042), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(new_n543), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1116));
  AOI21_X1  g691(.A(new_n1100), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1116), .B1(new_n1106), .B2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1103), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1103), .B(new_n598), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(KEYINPUT60), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1115), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n1123));
  AOI211_X1 g698(.A(new_n1123), .B(new_n1106), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1108), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1082), .A2(new_n1093), .A3(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1031), .A2(new_n1034), .A3(G286), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1073), .A2(new_n1052), .A3(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1044), .A2(G8), .A3(new_n1051), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1072), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1083), .A2(G8), .A3(G168), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1133), .A2(new_n1067), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1135), .A3(new_n1052), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1073), .A2(new_n1052), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT62), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1033), .A2(new_n1140), .A3(new_n1037), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .A4(new_n1019), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1052), .A2(new_n1067), .ZN(new_n1143));
  INV_X1    g718(.A(G288), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1060), .A2(new_n1062), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1054), .B1(new_n1145), .B2(new_n1056), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1143), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1137), .A2(new_n1142), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1126), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(G290), .A2(G1986), .ZN(new_n1150));
  OR3_X1    g725(.A1(new_n968), .A2(new_n960), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n948), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n976), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1152), .ZN(new_n1154));
  AOI211_X1 g729(.A(KEYINPUT125), .B(new_n1154), .C1(new_n1126), .C2(new_n1148), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n975), .B1(new_n1153), .B2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g731(.A(G319), .ZN(new_n1158));
  OR2_X1    g732(.A1(G227), .A2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g733(.A1(G229), .A2(G401), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1160), .A2(new_n849), .ZN(new_n1161));
  NOR2_X1   g735(.A1(new_n1161), .A2(new_n929), .ZN(G308));
  AND2_X1   g736(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n1163));
  OAI211_X1 g737(.A(new_n849), .B(new_n1160), .C1(new_n1163), .C2(new_n927), .ZN(G225));
endmodule


