

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  OR2_X1 U324 ( .A1(n470), .A2(n469), .ZN(n471) );
  XOR2_X1 U325 ( .A(KEYINPUT28), .B(n554), .Z(n518) );
  XNOR2_X1 U326 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U327 ( .A(n436), .B(n435), .Z(n292) );
  OR2_X1 U328 ( .A1(n573), .A2(n420), .ZN(n410) );
  XNOR2_X1 U329 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n341) );
  NOR2_X1 U330 ( .A1(n578), .A2(n506), .ZN(n507) );
  XOR2_X1 U331 ( .A(G113GAT), .B(KEYINPUT0), .Z(n380) );
  INV_X1 U332 ( .A(n427), .ZN(n389) );
  INV_X1 U333 ( .A(KEYINPUT26), .ZN(n408) );
  AND2_X1 U334 ( .A1(n473), .A2(n497), .ZN(n474) );
  XNOR2_X1 U335 ( .A(n409), .B(n408), .ZN(n531) );
  XNOR2_X1 U336 ( .A(n392), .B(n391), .ZN(n393) );
  NOR2_X1 U337 ( .A1(n573), .A2(n572), .ZN(n584) );
  XOR2_X1 U338 ( .A(n443), .B(n442), .Z(n569) );
  XNOR2_X1 U339 ( .A(KEYINPUT38), .B(n475), .ZN(n481) );
  XOR2_X1 U340 ( .A(KEYINPUT95), .B(G57GAT), .Z(n294) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G148GAT), .Z(n336) );
  XNOR2_X1 U342 ( .A(n380), .B(n336), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U344 ( .A(n295), .B(G85GAT), .Z(n301) );
  XNOR2_X1 U345 ( .A(G1GAT), .B(G127GAT), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n296), .B(G155GAT), .ZN(n447) );
  XOR2_X1 U347 ( .A(G29GAT), .B(KEYINPUT81), .Z(n436) );
  XOR2_X1 U348 ( .A(n447), .B(n436), .Z(n298) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U351 ( .A(G134GAT), .B(n299), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U353 ( .A(KEYINPUT97), .B(KEYINPUT1), .Z(n303) );
  XNOR2_X1 U354 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U356 ( .A(n305), .B(n304), .Z(n314) );
  XNOR2_X1 U357 ( .A(KEYINPUT2), .B(KEYINPUT90), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n306), .B(KEYINPUT3), .ZN(n307) );
  XOR2_X1 U359 ( .A(n307), .B(KEYINPUT91), .Z(n309) );
  XNOR2_X1 U360 ( .A(G141GAT), .B(G162GAT), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n365) );
  XOR2_X1 U362 ( .A(KEYINPUT96), .B(KEYINPUT94), .Z(n311) );
  XNOR2_X1 U363 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n365), .B(n312), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n413) );
  XNOR2_X1 U367 ( .A(KEYINPUT98), .B(n413), .ZN(n552) );
  XOR2_X1 U368 ( .A(G8GAT), .B(G1GAT), .Z(n316) );
  XNOR2_X1 U369 ( .A(G141GAT), .B(G197GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n320) );
  XOR2_X1 U371 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n318) );
  XNOR2_X1 U372 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n317) );
  XNOR2_X1 U373 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U374 ( .A(n320), .B(n319), .Z(n325) );
  XOR2_X1 U375 ( .A(KEYINPUT68), .B(KEYINPUT72), .Z(n322) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U378 ( .A(KEYINPUT69), .B(n323), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n330) );
  XOR2_X1 U380 ( .A(G43GAT), .B(G29GAT), .Z(n328) );
  XNOR2_X1 U381 ( .A(G15GAT), .B(G22GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n326), .B(KEYINPUT71), .ZN(n448) );
  XNOR2_X1 U383 ( .A(G113GAT), .B(n448), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U385 ( .A(n330), .B(n329), .Z(n335) );
  XOR2_X1 U386 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n332) );
  XNOR2_X1 U387 ( .A(G50GAT), .B(G36GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U389 ( .A(KEYINPUT7), .B(n333), .Z(n443) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(n443), .ZN(n334) );
  XOR2_X1 U391 ( .A(n335), .B(n334), .Z(n532) );
  XOR2_X1 U392 ( .A(KEYINPUT31), .B(n336), .Z(n340) );
  XOR2_X1 U393 ( .A(G78GAT), .B(G204GAT), .Z(n338) );
  XNOR2_X1 U394 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n357) );
  XNOR2_X1 U396 ( .A(G176GAT), .B(n357), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n347) );
  INV_X1 U398 ( .A(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G85GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n435) );
  XOR2_X1 U401 ( .A(n435), .B(KEYINPUT77), .Z(n345) );
  NAND2_X1 U402 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U404 ( .A(n347), .B(n346), .Z(n355) );
  XOR2_X1 U405 ( .A(G64GAT), .B(KEYINPUT13), .Z(n349) );
  XNOR2_X1 U406 ( .A(G71GAT), .B(G57GAT), .ZN(n348) );
  XNOR2_X1 U407 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U408 ( .A(KEYINPUT73), .B(n350), .Z(n456) );
  XOR2_X1 U409 ( .A(KEYINPUT78), .B(KEYINPUT33), .Z(n352) );
  XNOR2_X1 U410 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n456), .B(n353), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n578) );
  NOR2_X1 U414 ( .A1(n532), .A2(n578), .ZN(n356) );
  XOR2_X1 U415 ( .A(n356), .B(KEYINPUT79), .Z(n473) );
  XOR2_X1 U416 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n407) );
  XOR2_X1 U417 ( .A(G155GAT), .B(n357), .Z(n359) );
  NAND2_X1 U418 ( .A1(G228GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U419 ( .A(n359), .B(n358), .ZN(n364) );
  XNOR2_X1 U420 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n360), .B(KEYINPUT88), .ZN(n361) );
  XOR2_X1 U422 ( .A(n361), .B(KEYINPUT89), .Z(n363) );
  XNOR2_X1 U423 ( .A(G197GAT), .B(G218GAT), .ZN(n362) );
  XNOR2_X1 U424 ( .A(n363), .B(n362), .ZN(n400) );
  XOR2_X1 U425 ( .A(n364), .B(n400), .Z(n367) );
  XNOR2_X1 U426 ( .A(G50GAT), .B(n365), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n375) );
  XOR2_X1 U428 ( .A(KEYINPUT87), .B(KEYINPUT24), .Z(n369) );
  XNOR2_X1 U429 ( .A(G22GAT), .B(KEYINPUT86), .ZN(n368) );
  XNOR2_X1 U430 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U431 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n371) );
  XNOR2_X1 U432 ( .A(G148GAT), .B(KEYINPUT23), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U434 ( .A(n373), .B(n372), .Z(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n554) );
  XNOR2_X1 U436 ( .A(G176GAT), .B(KEYINPUT18), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n376), .B(KEYINPUT17), .ZN(n377) );
  XOR2_X1 U438 ( .A(n377), .B(KEYINPUT19), .Z(n379) );
  XNOR2_X1 U439 ( .A(G169GAT), .B(G190GAT), .ZN(n378) );
  XOR2_X1 U440 ( .A(n379), .B(n378), .Z(n403) );
  XOR2_X1 U441 ( .A(n380), .B(G120GAT), .Z(n382) );
  NAND2_X1 U442 ( .A1(G227GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n392) );
  XOR2_X1 U444 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n384) );
  XNOR2_X1 U445 ( .A(G99GAT), .B(G183GAT), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U447 ( .A(G127GAT), .B(KEYINPUT83), .Z(n386) );
  XNOR2_X1 U448 ( .A(G15GAT), .B(G71GAT), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n390) );
  XOR2_X1 U451 ( .A(G43GAT), .B(G134GAT), .Z(n427) );
  XOR2_X2 U452 ( .A(n403), .B(n393), .Z(n557) );
  XOR2_X1 U453 ( .A(KEYINPUT77), .B(KEYINPUT99), .Z(n395) );
  NAND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n399) );
  XOR2_X1 U456 ( .A(G64GAT), .B(G92GAT), .Z(n397) );
  XNOR2_X1 U457 ( .A(G36GAT), .B(G204GAT), .ZN(n396) );
  XNOR2_X1 U458 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U459 ( .A(n399), .B(n398), .Z(n402) );
  XOR2_X1 U460 ( .A(G8GAT), .B(G183GAT), .Z(n451) );
  XNOR2_X1 U461 ( .A(n400), .B(n451), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U463 ( .A(n404), .B(n403), .Z(n547) );
  NOR2_X1 U464 ( .A1(n557), .A2(n547), .ZN(n405) );
  NOR2_X1 U465 ( .A1(n554), .A2(n405), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n411) );
  NAND2_X1 U467 ( .A1(n554), .A2(n557), .ZN(n409) );
  INV_X1 U468 ( .A(n531), .ZN(n573) );
  XNOR2_X1 U469 ( .A(n547), .B(KEYINPUT27), .ZN(n420) );
  NAND2_X1 U470 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U471 ( .A(KEYINPUT102), .B(n412), .ZN(n414) );
  NAND2_X1 U472 ( .A1(n414), .A2(n413), .ZN(n417) );
  INV_X1 U473 ( .A(n417), .ZN(n416) );
  INV_X1 U474 ( .A(KEYINPUT103), .ZN(n415) );
  NAND2_X1 U475 ( .A1(n416), .A2(n415), .ZN(n419) );
  NAND2_X1 U476 ( .A1(KEYINPUT103), .A2(n417), .ZN(n418) );
  NAND2_X1 U477 ( .A1(n419), .A2(n418), .ZN(n426) );
  INV_X1 U478 ( .A(n518), .ZN(n424) );
  XOR2_X1 U479 ( .A(KEYINPUT85), .B(n557), .Z(n422) );
  NOR2_X1 U480 ( .A1(n552), .A2(n420), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n421), .B(KEYINPUT100), .ZN(n516) );
  NAND2_X1 U482 ( .A1(n422), .A2(n516), .ZN(n423) );
  NOR2_X1 U483 ( .A1(n424), .A2(n423), .ZN(n425) );
  NOR2_X1 U484 ( .A1(n426), .A2(n425), .ZN(n470) );
  XNOR2_X1 U485 ( .A(n427), .B(G162GAT), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n428), .B(G218GAT), .ZN(n432) );
  XOR2_X1 U487 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n430) );
  XNOR2_X1 U488 ( .A(G106GAT), .B(KEYINPUT80), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n432), .B(n431), .Z(n441) );
  XOR2_X1 U491 ( .A(KEYINPUT64), .B(KEYINPUT11), .Z(n434) );
  XNOR2_X1 U492 ( .A(G190GAT), .B(KEYINPUT9), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n439) );
  NAND2_X1 U494 ( .A1(G232GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n292), .B(n437), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U497 ( .A(n441), .B(n440), .ZN(n442) );
  INV_X1 U498 ( .A(n569), .ZN(n544) );
  XOR2_X1 U499 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n445) );
  NAND2_X1 U500 ( .A1(G231GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U502 ( .A(n446), .B(KEYINPUT15), .Z(n450) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U505 ( .A(n452), .B(n451), .Z(n454) );
  XNOR2_X1 U506 ( .A(G211GAT), .B(G78GAT), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n455) );
  XOR2_X1 U508 ( .A(n456), .B(n455), .Z(n582) );
  NAND2_X1 U509 ( .A1(n544), .A2(n582), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n457), .B(KEYINPUT16), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT82), .ZN(n459) );
  NOR2_X1 U512 ( .A1(n470), .A2(n459), .ZN(n484) );
  NAND2_X1 U513 ( .A1(n473), .A2(n484), .ZN(n467) );
  NOR2_X1 U514 ( .A1(n552), .A2(n467), .ZN(n461) );
  XNOR2_X1 U515 ( .A(KEYINPUT34), .B(KEYINPUT104), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U517 ( .A(G1GAT), .B(n462), .Z(G1324GAT) );
  NOR2_X1 U518 ( .A1(n547), .A2(n467), .ZN(n464) );
  XNOR2_X1 U519 ( .A(G8GAT), .B(KEYINPUT105), .ZN(n463) );
  XNOR2_X1 U520 ( .A(n464), .B(n463), .ZN(G1325GAT) );
  NOR2_X1 U521 ( .A1(n557), .A2(n467), .ZN(n466) );
  XNOR2_X1 U522 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n466), .B(n465), .ZN(G1326GAT) );
  NOR2_X1 U524 ( .A1(n518), .A2(n467), .ZN(n468) );
  XOR2_X1 U525 ( .A(G22GAT), .B(n468), .Z(G1327GAT) );
  XOR2_X1 U526 ( .A(KEYINPUT106), .B(KEYINPUT37), .Z(n472) );
  XOR2_X1 U527 ( .A(KEYINPUT36), .B(n569), .Z(n586) );
  OR2_X1 U528 ( .A1(n582), .A2(n586), .ZN(n469) );
  XOR2_X1 U529 ( .A(n472), .B(n471), .Z(n497) );
  XNOR2_X1 U530 ( .A(n474), .B(KEYINPUT107), .ZN(n475) );
  NOR2_X1 U531 ( .A1(n481), .A2(n552), .ZN(n477) );
  XNOR2_X1 U532 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n477), .B(n476), .ZN(G1328GAT) );
  NOR2_X1 U534 ( .A1(n481), .A2(n547), .ZN(n478) );
  XOR2_X1 U535 ( .A(G36GAT), .B(n478), .Z(G1329GAT) );
  NOR2_X1 U536 ( .A1(n481), .A2(n557), .ZN(n479) );
  XOR2_X1 U537 ( .A(n479), .B(KEYINPUT40), .Z(n480) );
  XNOR2_X1 U538 ( .A(G43GAT), .B(n480), .ZN(G1330GAT) );
  NOR2_X1 U539 ( .A1(n481), .A2(n518), .ZN(n482) );
  XOR2_X1 U540 ( .A(G50GAT), .B(n482), .Z(G1331GAT) );
  XNOR2_X1 U541 ( .A(n578), .B(KEYINPUT41), .ZN(n535) );
  INV_X1 U542 ( .A(n535), .ZN(n563) );
  NAND2_X1 U543 ( .A1(n532), .A2(n563), .ZN(n483) );
  XOR2_X1 U544 ( .A(n483), .B(KEYINPUT108), .Z(n496) );
  NAND2_X1 U545 ( .A1(n484), .A2(n496), .ZN(n492) );
  NOR2_X1 U546 ( .A1(n552), .A2(n492), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G57GAT), .B(n487), .ZN(G1332GAT) );
  NOR2_X1 U550 ( .A1(n547), .A2(n492), .ZN(n488) );
  XOR2_X1 U551 ( .A(KEYINPUT110), .B(n488), .Z(n489) );
  XNOR2_X1 U552 ( .A(G64GAT), .B(n489), .ZN(G1333GAT) );
  NOR2_X1 U553 ( .A1(n557), .A2(n492), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n490) );
  XNOR2_X1 U555 ( .A(n491), .B(n490), .ZN(G1334GAT) );
  NOR2_X1 U556 ( .A1(n518), .A2(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G78GAT), .B(n495), .ZN(G1335GAT) );
  NAND2_X1 U560 ( .A1(n497), .A2(n496), .ZN(n501) );
  NOR2_X1 U561 ( .A1(n552), .A2(n501), .ZN(n498) );
  XOR2_X1 U562 ( .A(G85GAT), .B(n498), .Z(G1336GAT) );
  NOR2_X1 U563 ( .A1(n547), .A2(n501), .ZN(n499) );
  XOR2_X1 U564 ( .A(G92GAT), .B(n499), .Z(G1337GAT) );
  NOR2_X1 U565 ( .A1(n557), .A2(n501), .ZN(n500) );
  XOR2_X1 U566 ( .A(G99GAT), .B(n500), .Z(G1338GAT) );
  NOR2_X1 U567 ( .A1(n518), .A2(n501), .ZN(n502) );
  XOR2_X1 U568 ( .A(KEYINPUT44), .B(n502), .Z(n503) );
  XNOR2_X1 U569 ( .A(G106GAT), .B(n503), .ZN(G1339GAT) );
  INV_X1 U570 ( .A(n532), .ZN(n574) );
  INV_X1 U571 ( .A(n582), .ZN(n541) );
  NOR2_X1 U572 ( .A1(n586), .A2(n541), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n504), .B(KEYINPUT45), .ZN(n505) );
  NAND2_X1 U574 ( .A1(n505), .A2(n532), .ZN(n506) );
  XNOR2_X1 U575 ( .A(KEYINPUT115), .B(n507), .ZN(n514) );
  XOR2_X1 U576 ( .A(KEYINPUT47), .B(KEYINPUT114), .Z(n512) );
  XOR2_X1 U577 ( .A(KEYINPUT113), .B(n582), .Z(n566) );
  NAND2_X1 U578 ( .A1(n574), .A2(n563), .ZN(n508) );
  XOR2_X1 U579 ( .A(KEYINPUT46), .B(n508), .Z(n509) );
  NOR2_X1 U580 ( .A1(n566), .A2(n509), .ZN(n510) );
  NAND2_X1 U581 ( .A1(n510), .A2(n544), .ZN(n511) );
  XNOR2_X1 U582 ( .A(n512), .B(n511), .ZN(n513) );
  NAND2_X1 U583 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n515), .B(KEYINPUT48), .ZN(n548) );
  NAND2_X1 U585 ( .A1(n516), .A2(n548), .ZN(n517) );
  XOR2_X1 U586 ( .A(KEYINPUT116), .B(n517), .Z(n530) );
  NAND2_X1 U587 ( .A1(n518), .A2(n530), .ZN(n519) );
  NOR2_X1 U588 ( .A1(n557), .A2(n519), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n574), .A2(n526), .ZN(n520) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n520), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n522) );
  NAND2_X1 U592 ( .A1(n526), .A2(n563), .ZN(n521) );
  XNOR2_X1 U593 ( .A(n522), .B(n521), .ZN(G1341GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n524) );
  NAND2_X1 U595 ( .A1(n526), .A2(n566), .ZN(n523) );
  XNOR2_X1 U596 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n525), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n528) );
  NAND2_X1 U599 ( .A1(n526), .A2(n569), .ZN(n527) );
  XNOR2_X1 U600 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n529), .ZN(G1343GAT) );
  NAND2_X1 U602 ( .A1(n531), .A2(n530), .ZN(n543) );
  NOR2_X1 U603 ( .A1(n532), .A2(n543), .ZN(n534) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n533) );
  XNOR2_X1 U605 ( .A(n534), .B(n533), .ZN(G1344GAT) );
  NOR2_X1 U606 ( .A1(n535), .A2(n543), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n537) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n536) );
  XNOR2_X1 U609 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U610 ( .A(KEYINPUT52), .B(n538), .ZN(n539) );
  XNOR2_X1 U611 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n541), .A2(n543), .ZN(n542) );
  XOR2_X1 U613 ( .A(G155GAT), .B(n542), .Z(G1346GAT) );
  NOR2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U615 ( .A(KEYINPUT122), .B(n545), .Z(n546) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n546), .ZN(G1347GAT) );
  XNOR2_X1 U617 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n559) );
  INV_X1 U618 ( .A(n547), .ZN(n549) );
  NAND2_X1 U619 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n550), .B(KEYINPUT54), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n551), .B(KEYINPUT123), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n572) );
  NOR2_X1 U623 ( .A1(n554), .A2(n572), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT55), .ZN(n556) );
  NOR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n574), .A2(n568), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT126), .Z(n561) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT125), .B(n562), .Z(n565) );
  NAND2_X1 U632 ( .A1(n568), .A2(n563), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  NAND2_X1 U640 ( .A1(n584), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .ZN(n588) );
  INV_X1 U652 ( .A(n588), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

