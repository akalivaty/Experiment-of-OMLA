//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n558, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1228, new_n1229;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XOR2_X1   g011(.A(new_n436), .B(KEYINPUT66), .Z(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n437), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  OR4_X1    g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(KEYINPUT3), .B2(new_n461), .ZN(new_n462));
  NOR3_X1   g037(.A1(new_n458), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n459), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(new_n459), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g050(.A(KEYINPUT69), .B(new_n459), .C1(new_n462), .C2(new_n463), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n475), .A2(G2105), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n467), .A3(new_n476), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n477), .A2(KEYINPUT70), .A3(G124), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n480), .A2(new_n483), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(new_n467), .A2(G138), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n459), .B(new_n490), .C1(new_n462), .C2(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n468), .A2(new_n459), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n459), .B(new_n497), .C1(new_n462), .C2(new_n463), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n496), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n510), .A2(G651), .B1(G50), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n505), .B(new_n507), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n511), .A2(new_n512), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(G88), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n514), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n513), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n518), .A2(G89), .A3(new_n522), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n508), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G651), .B1(G52), .B2(new_n513), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n518), .A2(G90), .A3(new_n522), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n518), .A2(G81), .A3(new_n522), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n513), .A2(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n505), .A2(new_n507), .A3(G56), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n545), .A2(KEYINPUT72), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT72), .B1(new_n545), .B2(new_n546), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  NOR3_X1   g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n541), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n548), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n545), .A2(KEYINPUT72), .A3(new_n546), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n552), .A2(G651), .A3(new_n553), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n554), .A2(KEYINPUT73), .A3(new_n543), .A4(new_n542), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  OAI211_X1 g137(.A(KEYINPUT74), .B(G543), .C1(new_n515), .C2(new_n516), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n566), .A4(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT75), .B1(new_n569), .B2(new_n549), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n518), .A2(G91), .A3(new_n522), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n508), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n574), .A2(new_n575), .A3(G651), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(new_n576), .ZN(G299));
  OAI21_X1  g152(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n513), .A2(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n518), .A2(new_n522), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(G288));
  AND3_X1   g157(.A1(new_n518), .A2(G86), .A3(new_n522), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n508), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G651), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n513), .A2(G48), .ZN(new_n589));
  AND2_X1   g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n584), .A2(new_n590), .ZN(G305));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n505), .A2(new_n507), .A3(G60), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n593), .A2(KEYINPUT76), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(KEYINPUT76), .B1(new_n593), .B2(new_n594), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n592), .B1(new_n598), .B2(G651), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n593), .A2(new_n594), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n602), .A2(new_n592), .A3(G651), .A4(new_n595), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n518), .A2(G85), .A3(new_n522), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n513), .A2(G47), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n605), .A2(KEYINPUT78), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT78), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n599), .A2(new_n604), .B1(new_n607), .B2(new_n608), .ZN(G290));
  NAND3_X1  g184(.A1(new_n518), .A2(G92), .A3(new_n522), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT80), .B(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n508), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(G54), .B2(new_n513), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n518), .A2(new_n522), .A3(new_n616), .A4(G92), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n611), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n611), .A2(new_n615), .A3(new_n617), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G868), .ZN(new_n625));
  NOR2_X1   g200(.A1(G171), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(KEYINPUT79), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(KEYINPUT79), .B2(new_n626), .ZN(G321));
  XOR2_X1   g203(.A(G321), .B(KEYINPUT82), .Z(G284));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  XOR2_X1   g207(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n623), .B1(new_n634), .B2(G860), .ZN(G148));
  INV_X1    g210(.A(new_n556), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(new_n625), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n619), .A2(new_n622), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n638), .A2(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n637), .B1(new_n639), .B2(new_n625), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n482), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n477), .A2(G123), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT85), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2096), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n649));
  NOR3_X1   g224(.A1(new_n458), .A2(new_n461), .A3(G2105), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2100), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2435), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2438), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1341), .B(G1348), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(G14), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n671), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT18), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n672), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n672), .B(KEYINPUT17), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n677), .B(new_n674), .C1(new_n671), .C2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n671), .A2(new_n678), .A3(new_n673), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n676), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2100), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT19), .Z(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n691), .A2(new_n692), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n694), .B(new_n695), .C1(new_n692), .C2(new_n691), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(G1986), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT22), .B(G1981), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  INV_X1    g278(.A(KEYINPUT94), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT92), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G24), .ZN(new_n707));
  INV_X1    g282(.A(G290), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(new_n706), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G1986), .ZN(new_n710));
  INV_X1    g285(.A(G1986), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n711), .B(new_n707), .C1(new_n708), .C2(new_n706), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n706), .A2(G6), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G305), .B2(G16), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT88), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT32), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n706), .B1(new_n584), .B2(new_n590), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n716), .B1(new_n719), .B2(new_n713), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(G16), .A2(G23), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT89), .Z(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G288), .B2(new_n706), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1971), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n706), .B1(new_n514), .B2(new_n523), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n706), .A2(G22), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT90), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT91), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n728), .A2(KEYINPUT91), .A3(new_n730), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n727), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n733), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n735), .A2(G1971), .A3(new_n731), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n721), .A2(new_n726), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n710), .B(new_n712), .C1(new_n737), .C2(KEYINPUT34), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n482), .A2(G131), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n477), .A2(G119), .ZN(new_n742));
  OR2_X1    g317(.A1(G95), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT35), .B(G1991), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n705), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n710), .A2(new_n712), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n734), .A2(new_n736), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT34), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n752), .A2(new_n753), .A3(new_n721), .A4(new_n726), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n751), .A2(new_n754), .A3(KEYINPUT92), .A4(new_n748), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n737), .A2(KEYINPUT34), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n704), .B1(new_n756), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(KEYINPUT94), .B(new_n759), .C1(new_n750), .C2(new_n755), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n762), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n482), .A2(G141), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n477), .A2(G129), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT97), .Z(new_n770));
  XOR2_X1   g345(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND4_X1  g348(.A1(new_n767), .A2(new_n768), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(new_n739), .ZN(new_n775));
  NOR2_X1   g350(.A1(G29), .A2(G32), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT27), .B(G1996), .Z(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  OR2_X1    g354(.A1(G5), .A2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G301), .B2(new_n706), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n777), .A2(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n706), .A2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G168), .B2(new_n706), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1966), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n781), .A2(new_n779), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n642), .A2(new_n643), .A3(G29), .A4(new_n645), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT31), .B(G11), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(G28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(G28), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n790), .A2(new_n791), .A3(new_n739), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n786), .A2(new_n787), .A3(new_n788), .A4(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT99), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G1966), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n784), .B(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT99), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n787), .A2(new_n788), .A3(new_n792), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n796), .A2(new_n797), .A3(new_n786), .A4(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n778), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n775), .B2(new_n776), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n782), .A2(new_n794), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n739), .A2(G27), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G164), .B2(new_n739), .ZN(new_n805));
  INV_X1    g380(.A(G2078), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n482), .A2(G139), .ZN(new_n808));
  NAND2_X1  g383(.A1(G115), .A2(G2104), .ZN(new_n809));
  INV_X1    g384(.A(G127), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n493), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G2105), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT25), .Z(new_n814));
  NAND3_X1  g389(.A1(new_n808), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n808), .A2(KEYINPUT96), .A3(new_n812), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G29), .ZN(new_n820));
  INV_X1    g395(.A(G2072), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n739), .A2(G33), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n821), .B1(new_n820), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g400(.A1(KEYINPUT24), .A2(G34), .ZN(new_n826));
  NOR2_X1   g401(.A1(KEYINPUT24), .A2(G34), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n826), .A2(new_n827), .A3(G29), .ZN(new_n828));
  INV_X1    g403(.A(G160), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(G29), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G2084), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n803), .A2(new_n807), .A3(new_n825), .A4(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n802), .A2(new_n824), .A3(new_n823), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n835), .A2(KEYINPUT100), .A3(new_n807), .A4(new_n831), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n739), .A2(G35), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n487), .B2(G29), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT29), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n840));
  INV_X1    g415(.A(G2090), .ZN(new_n841));
  AND3_X1   g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT23), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n706), .A2(G20), .ZN(new_n844));
  AOI22_X1  g419(.A1(G299), .A2(G16), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(G1956), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT95), .B(G1341), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n636), .A2(G16), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n706), .A2(G19), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(new_n848), .A3(new_n850), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(new_n853), .C1(new_n839), .C2(new_n841), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n840), .B1(new_n839), .B2(new_n841), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n842), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n834), .A2(new_n836), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  OAI22_X1  g433(.A1(new_n761), .A2(new_n763), .B1(KEYINPUT93), .B2(KEYINPUT36), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n739), .A2(G26), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n482), .A2(G140), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n477), .A2(G128), .ZN(new_n862));
  NOR2_X1   g437(.A1(G104), .A2(G2105), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n861), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n860), .B1(new_n865), .B2(G29), .ZN(new_n866));
  MUX2_X1   g441(.A(new_n860), .B(new_n866), .S(KEYINPUT28), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G2067), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n766), .A2(new_n858), .A3(new_n859), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n706), .A2(G4), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n623), .B2(new_n706), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G1348), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n869), .A2(new_n872), .ZN(G311));
  NOR2_X1   g448(.A1(new_n761), .A2(new_n763), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n857), .B1(new_n874), .B2(new_n765), .ZN(new_n875));
  INV_X1    g450(.A(new_n872), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n875), .A2(new_n868), .A3(new_n859), .A4(new_n876), .ZN(G150));
  NAND2_X1  g452(.A1(G80), .A2(G543), .ZN(new_n878));
  INV_X1    g453(.A(G67), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n508), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G651), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n513), .A2(G55), .ZN(new_n882));
  INV_X1    g457(.A(G93), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n881), .B(new_n882), .C1(new_n580), .C2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(G860), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT37), .Z(new_n886));
  NAND2_X1  g461(.A1(new_n623), .A2(G559), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT38), .ZN(new_n888));
  INV_X1    g463(.A(new_n884), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n889), .B1(new_n551), .B2(new_n555), .ZN(new_n890));
  INV_X1    g465(.A(new_n544), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n884), .B1(new_n891), .B2(new_n554), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n888), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(KEYINPUT102), .A3(KEYINPUT39), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G860), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n895), .B2(KEYINPUT39), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT102), .B1(new_n895), .B2(KEYINPUT39), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  NOR4_X1   g478(.A1(new_n897), .A2(new_n899), .A3(new_n900), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n886), .B1(new_n902), .B2(new_n904), .ZN(G145));
  XNOR2_X1  g480(.A(new_n646), .B(G160), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(new_n487), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n482), .A2(G142), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n908), .B(KEYINPUT106), .Z(new_n909));
  OR2_X1    g484(.A1(G106), .A2(G2105), .ZN(new_n910));
  INV_X1    g485(.A(G118), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n461), .B1(new_n911), .B2(G2105), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n477), .A2(G130), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n745), .B(new_n651), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n914), .B(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  AND3_X1   g492(.A1(new_n498), .A2(new_n917), .A3(new_n500), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n917), .B1(new_n498), .B2(new_n500), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n496), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n865), .B(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n817), .A2(KEYINPUT105), .A3(new_n818), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n774), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n920), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n865), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n819), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(KEYINPUT105), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n774), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n922), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n916), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n907), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n916), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n925), .A2(new_n916), .A3(new_n932), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(KEYINPUT107), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n940), .A3(new_n907), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n605), .A2(new_n606), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT78), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n605), .A2(KEYINPUT78), .A3(new_n606), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n602), .A2(G651), .A3(new_n595), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT77), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n603), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n951), .A2(G288), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G288), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n946), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(G305), .B(G303), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G288), .ZN(new_n960));
  NAND2_X1  g535(.A1(G290), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(G288), .A3(new_n954), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(KEYINPUT108), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n958), .B(new_n946), .C1(new_n955), .C2(new_n956), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT42), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(KEYINPUT42), .A3(new_n965), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n894), .A2(new_n639), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT41), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n620), .A2(G299), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n620), .A2(G299), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n618), .A2(new_n631), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n620), .A2(G299), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n975), .A2(KEYINPUT41), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n893), .B1(G559), .B2(new_n638), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n970), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n970), .A2(new_n979), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n972), .A2(new_n973), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n969), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n969), .A2(new_n983), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n625), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n889), .A2(G868), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(G295));
  XNOR2_X1  g564(.A(new_n988), .B(KEYINPUT109), .ZN(G331));
  NAND3_X1  g565(.A1(G286), .A2(new_n538), .A3(new_n537), .ZN(new_n991));
  NAND3_X1  g566(.A1(G301), .A2(new_n531), .A3(new_n530), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n556), .A2(new_n884), .ZN(new_n994));
  INV_X1    g569(.A(new_n892), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n991), .A2(new_n992), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n890), .A2(new_n997), .A3(new_n892), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n978), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(new_n995), .A3(new_n993), .ZN(new_n1000));
  INV_X1    g575(.A(new_n982), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n890), .B2(new_n892), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n965), .A3(new_n964), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n964), .A2(new_n965), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1006), .A2(new_n999), .A3(new_n1003), .ZN(new_n1007));
  INV_X1    g582(.A(G37), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n1011));
  AOI21_X1  g586(.A(G37), .B1(new_n1004), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1006), .A2(KEYINPUT111), .A3(new_n999), .A4(new_n1003), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n1005), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1010), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT112), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT112), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1019), .A3(KEYINPUT43), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1022));
  AND3_X1   g597(.A1(new_n1021), .A2(KEYINPUT113), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT113), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1015), .B1(new_n1023), .B2(new_n1024), .ZN(G397));
  AND2_X1   g600(.A1(new_n865), .A2(G2067), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n865), .A2(G2067), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n1028));
  OR3_X1    g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1030));
  INV_X1    g605(.A(G1996), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n774), .B(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT114), .B(G1384), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n920), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G40), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n829), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT116), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1033), .A2(new_n1042), .A3(new_n1039), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n745), .A2(new_n747), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n745), .A2(new_n747), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1039), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(G290), .B(G1986), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1039), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT62), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n920), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n466), .A2(new_n1038), .A3(new_n471), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n494), .B1(KEYINPUT4), .B2(new_n491), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n498), .A2(new_n500), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1053), .A2(new_n1054), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G2084), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n501), .A2(new_n1062), .A3(KEYINPUT45), .A4(new_n1052), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT45), .B(new_n1052), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT120), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1056), .A2(KEYINPUT104), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n498), .A2(new_n917), .A3(new_n500), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(G1384), .B1(new_n1070), .B2(new_n496), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1067), .B(new_n1054), .C1(new_n1071), .C2(KEYINPUT45), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n920), .A2(new_n1054), .A3(new_n1052), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1054), .A2(KEYINPUT45), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(KEYINPUT119), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1066), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1061), .B1(new_n1076), .B2(G1966), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT123), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1061), .B(new_n1079), .C1(new_n1076), .C2(G1966), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(KEYINPUT51), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1066), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1060), .B1(new_n1084), .B2(new_n795), .ZN(new_n1085));
  OAI21_X1  g660(.A(G168), .B1(new_n1085), .B2(KEYINPUT51), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(G8), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1078), .A2(G168), .A3(new_n1080), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1050), .B(new_n1087), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1081), .A2(G8), .A3(new_n1086), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1090), .B1(new_n1088), .B2(G8), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT62), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G8), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1071), .B2(new_n1054), .ZN(new_n1096));
  INV_X1    g671(.A(G1981), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n584), .A2(new_n590), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n588), .A2(new_n589), .ZN(new_n1099));
  OAI21_X1  g674(.A(G1981), .B1(new_n1099), .B2(new_n583), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT49), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1098), .A2(new_n1100), .A3(KEYINPUT49), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1096), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n960), .A2(G1976), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1073), .A2(new_n1106), .A3(G8), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT52), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(new_n960), .B2(G1976), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1105), .B(new_n1108), .C1(new_n1107), .C2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n920), .A2(KEYINPUT45), .A3(new_n1034), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1057), .A2(new_n1036), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1054), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n727), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1053), .A2(new_n1058), .A3(new_n841), .A4(new_n1054), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1095), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(KEYINPUT117), .A2(KEYINPUT55), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1119));
  NAND2_X1  g694(.A1(G303), .A2(G8), .ZN(new_n1120));
  MUX2_X1   g695(.A(new_n1118), .B(new_n1119), .S(new_n1120), .Z(new_n1121));
  AOI21_X1  g696(.A(new_n1111), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1051), .B1(new_n920), .B2(new_n1052), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1051), .B(new_n1052), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1054), .ZN(new_n1126));
  OR3_X1    g701(.A1(new_n1124), .A2(new_n1126), .A3(G2090), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1095), .B1(new_n1127), .B2(new_n1115), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1123), .B1(new_n1128), .B2(new_n1121), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1121), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1127), .A2(new_n1115), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT118), .B(new_n1130), .C1(new_n1131), .C2(new_n1095), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1122), .A2(new_n1129), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n806), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1114), .B2(G2078), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT124), .B(G1961), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1059), .A2(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1133), .A2(new_n1140), .A3(G301), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1091), .A2(new_n1094), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1117), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1143), .A2(new_n1111), .A3(new_n1130), .ZN(new_n1144));
  INV_X1    g719(.A(G1976), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1105), .A2(new_n1145), .A3(new_n960), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1098), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1096), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT63), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1077), .A2(G8), .A3(G168), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1133), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1149), .B1(new_n1143), .B2(new_n1130), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1122), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1152), .B1(new_n1154), .B2(new_n1150), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1150), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1156), .A2(KEYINPUT121), .A3(new_n1122), .A4(new_n1153), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1151), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(G301), .B(KEYINPUT54), .Z(new_n1159));
  NOR2_X1   g734(.A1(new_n1135), .A2(G2078), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1037), .A2(new_n1054), .A3(new_n1112), .A4(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1139), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1122), .A2(new_n1132), .A3(new_n1129), .A4(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1140), .A2(new_n1159), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT58), .B(G1341), .Z(new_n1167));
  NAND2_X1  g742(.A1(new_n1073), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT122), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1073), .A2(new_n1170), .A3(new_n1167), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1169), .B(new_n1171), .C1(G1996), .C2(new_n1114), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n556), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(KEYINPUT59), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1172), .A2(new_n1175), .A3(new_n556), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G1956), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1179));
  XOR2_X1   g754(.A(G299), .B(KEYINPUT57), .Z(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT56), .B(G2072), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1112), .A2(new_n1113), .A3(new_n1054), .A4(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1180), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1185));
  OAI21_X1  g760(.A(KEYINPUT61), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1180), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1183), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1186), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(G1348), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1059), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT60), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1073), .A2(G2067), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1194), .A2(new_n623), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1194), .A2(new_n638), .A3(new_n1196), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n638), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1199));
  OAI21_X1  g774(.A(KEYINPUT60), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1177), .A2(new_n1192), .A3(new_n1197), .A4(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1199), .A2(new_n1183), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1201), .A2(new_n1202), .A3(new_n1189), .ZN(new_n1203));
  OAI211_X1 g778(.A(new_n1148), .B(new_n1158), .C1(new_n1166), .C2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1049), .B1(new_n1142), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1047), .A2(KEYINPUT126), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1041), .A2(new_n1207), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1039), .A2(new_n711), .A3(new_n708), .ZN(new_n1209));
  XOR2_X1   g784(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1210));
  XNOR2_X1  g785(.A(new_n1209), .B(new_n1210), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1206), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1039), .B1(new_n1213), .B2(new_n1027), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1039), .A2(new_n1031), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT46), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1029), .A2(new_n930), .A3(new_n1030), .ZN(new_n1217));
  AND3_X1   g792(.A1(new_n1217), .A2(KEYINPUT125), .A3(new_n1039), .ZN(new_n1218));
  AOI21_X1  g793(.A(KEYINPUT125), .B1(new_n1217), .B2(new_n1039), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1216), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1220), .A2(KEYINPUT47), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT47), .ZN(new_n1222));
  OAI211_X1 g797(.A(new_n1222), .B(new_n1216), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n1212), .A2(new_n1214), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1205), .A2(new_n1225), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g801(.A(new_n683), .B1(new_n666), .B2(new_n667), .ZN(new_n1228));
  AOI21_X1  g802(.A(new_n1228), .B1(new_n942), .B2(new_n943), .ZN(new_n1229));
  NAND4_X1  g803(.A1(new_n1229), .A2(new_n702), .A3(G319), .A4(new_n1021), .ZN(G225));
  INV_X1    g804(.A(G225), .ZN(G308));
endmodule


