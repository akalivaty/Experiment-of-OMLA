

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750;

  XOR2_X1 U365 ( .A(n706), .B(n705), .Z(n367) );
  XNOR2_X1 U366 ( .A(n393), .B(n362), .ZN(n621) );
  NAND2_X1 U367 ( .A1(n343), .A2(n610), .ZN(n393) );
  XNOR2_X1 U368 ( .A(n573), .B(KEYINPUT1), .ZN(n663) );
  INV_X1 U369 ( .A(G125), .ZN(n484) );
  INV_X1 U370 ( .A(G104), .ZN(n403) );
  XNOR2_X2 U371 ( .A(n402), .B(n401), .ZN(n724) );
  XOR2_X2 U372 ( .A(KEYINPUT15), .B(G902), .Z(n524) );
  XOR2_X2 U373 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n364) );
  XNOR2_X2 U374 ( .A(n342), .B(KEYINPUT39), .ZN(n596) );
  NAND2_X1 U375 ( .A1(n345), .A2(n478), .ZN(n342) );
  XNOR2_X2 U376 ( .A(KEYINPUT4), .B(KEYINPUT68), .ZN(n733) );
  XNOR2_X2 U377 ( .A(n585), .B(KEYINPUT41), .ZN(n674) );
  XNOR2_X2 U378 ( .A(n436), .B(n528), .ZN(n623) );
  XNOR2_X1 U379 ( .A(n517), .B(KEYINPUT91), .ZN(n428) );
  NOR2_X1 U380 ( .A1(n607), .A2(n577), .ZN(n417) );
  AND2_X2 U381 ( .A1(n591), .A2(n745), .ZN(n349) );
  AND2_X2 U382 ( .A1(n383), .A2(n381), .ZN(n380) );
  XNOR2_X2 U383 ( .A(n347), .B(n595), .ZN(n346) );
  AND2_X2 U384 ( .A1(n575), .A2(n678), .ZN(n345) );
  XOR2_X2 U385 ( .A(G472), .B(n540), .Z(n617) );
  XNOR2_X2 U386 ( .A(n398), .B(n434), .ZN(n721) );
  XNOR2_X1 U387 ( .A(n428), .B(n518), .ZN(n541) );
  INV_X4 U388 ( .A(G953), .ZN(n737) );
  NOR2_X1 U389 ( .A1(n578), .A2(n579), .ZN(n369) );
  NOR2_X1 U390 ( .A1(n632), .A2(G902), .ZN(n540) );
  XNOR2_X1 U391 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n452) );
  XNOR2_X1 U392 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n453) );
  XNOR2_X1 U393 ( .A(n369), .B(n458), .ZN(n348) );
  NOR2_X1 U394 ( .A1(n656), .A2(n433), .ZN(n432) );
  BUF_X1 U395 ( .A(n747), .Z(n748) );
  XNOR2_X1 U396 ( .A(n443), .B(n363), .ZN(n747) );
  XNOR2_X1 U397 ( .A(n620), .B(KEYINPUT99), .ZN(n635) );
  XNOR2_X1 U398 ( .A(n616), .B(KEYINPUT31), .ZN(n651) );
  NAND2_X1 U399 ( .A1(n396), .A2(n395), .ZN(n478) );
  XNOR2_X1 U400 ( .A(n617), .B(n464), .ZN(n624) );
  XOR2_X1 U401 ( .A(n632), .B(KEYINPUT62), .Z(n365) );
  XNOR2_X1 U402 ( .A(n491), .B(n359), .ZN(n490) );
  XNOR2_X1 U403 ( .A(n548), .B(n547), .ZN(n449) );
  XNOR2_X1 U404 ( .A(n736), .B(n533), .ZN(n547) );
  XNOR2_X1 U405 ( .A(n403), .B(G110), .ZN(n402) );
  XNOR2_X1 U406 ( .A(n453), .B(n452), .ZN(n451) );
  XNOR2_X1 U407 ( .A(n733), .B(n404), .ZN(n450) );
  XNOR2_X1 U408 ( .A(KEYINPUT67), .B(G101), .ZN(n404) );
  XNOR2_X1 U409 ( .A(G107), .B(KEYINPUT78), .ZN(n401) );
  NAND2_X1 U410 ( .A1(n343), .A2(n657), .ZN(n445) );
  XNOR2_X2 U411 ( .A(n439), .B(n364), .ZN(n343) );
  AND2_X2 U412 ( .A1(n596), .A2(n646), .ZN(n588) );
  NAND2_X1 U413 ( .A1(n346), .A2(n432), .ZN(n405) );
  NAND2_X1 U414 ( .A1(n349), .A2(n348), .ZN(n347) );
  NOR2_X2 U415 ( .A1(n586), .A2(n564), .ZN(n644) );
  BUF_X1 U416 ( .A(n663), .Z(n350) );
  INV_X1 U417 ( .A(n655), .ZN(n433) );
  XNOR2_X1 U418 ( .A(n592), .B(n563), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n592), .B(n563), .ZN(n603) );
  NAND2_X1 U420 ( .A1(n351), .A2(n602), .ZN(n352) );
  NAND2_X1 U421 ( .A1(n603), .A2(n602), .ZN(n439) );
  XNOR2_X2 U422 ( .A(n353), .B(n354), .ZN(n749) );
  NAND2_X1 U423 ( .A1(n469), .A2(n621), .ZN(n353) );
  XNOR2_X1 U424 ( .A(KEYINPUT65), .B(n614), .ZN(n354) );
  NAND2_X1 U425 ( .A1(n380), .A2(n379), .ZN(n382) );
  NOR2_X1 U426 ( .A1(G237), .A2(G902), .ZN(n504) );
  INV_X1 U427 ( .A(G469), .ZN(n474) );
  NAND2_X1 U428 ( .A1(G214), .A2(n554), .ZN(n677) );
  XNOR2_X1 U429 ( .A(n463), .B(KEYINPUT108), .ZN(n593) );
  NAND2_X1 U430 ( .A1(n465), .A2(n624), .ZN(n463) );
  OR2_X1 U431 ( .A1(n710), .A2(G902), .ZN(n407) );
  XNOR2_X1 U432 ( .A(n566), .B(n459), .ZN(n409) );
  INV_X1 U433 ( .A(KEYINPUT88), .ZN(n459) );
  NAND2_X1 U434 ( .A1(n388), .A2(n387), .ZN(n386) );
  INV_X1 U435 ( .A(n651), .ZN(n388) );
  INV_X1 U436 ( .A(n635), .ZN(n387) );
  NAND2_X1 U437 ( .A1(G237), .A2(G234), .ZN(n509) );
  INV_X1 U438 ( .A(KEYINPUT75), .ZN(n458) );
  NAND2_X1 U439 ( .A1(n574), .A2(n483), .ZN(n481) );
  XOR2_X1 U440 ( .A(KEYINPUT72), .B(G119), .Z(n497) );
  INV_X1 U441 ( .A(KEYINPUT45), .ZN(n434) );
  NAND2_X1 U442 ( .A1(n382), .A2(n399), .ZN(n398) );
  XNOR2_X1 U443 ( .A(n414), .B(n413), .ZN(n412) );
  XNOR2_X1 U444 ( .A(KEYINPUT102), .B(G122), .ZN(n414) );
  XNOR2_X1 U445 ( .A(G107), .B(G116), .ZN(n413) );
  XNOR2_X1 U446 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n411) );
  XNOR2_X1 U447 ( .A(n378), .B(n454), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n456), .B(n455), .ZN(n454) );
  XNOR2_X1 U449 ( .A(n451), .B(n546), .ZN(n378) );
  NAND2_X1 U450 ( .A1(n375), .A2(n374), .ZN(n373) );
  NOR2_X1 U451 ( .A1(n418), .A2(KEYINPUT36), .ZN(n374) );
  AND2_X1 U452 ( .A1(n372), .A2(n376), .ZN(n371) );
  AND2_X1 U453 ( .A1(n617), .A2(n558), .ZN(n559) );
  INV_X1 U454 ( .A(G478), .ZN(n461) );
  OR2_X1 U455 ( .A1(n713), .A2(G902), .ZN(n408) );
  XNOR2_X1 U456 ( .A(n527), .B(n526), .ZN(n528) );
  INV_X1 U457 ( .A(KEYINPUT25), .ZN(n526) );
  INV_X1 U458 ( .A(KEYINPUT6), .ZN(n464) );
  BUF_X1 U459 ( .A(n350), .Z(n427) );
  INV_X1 U460 ( .A(KEYINPUT64), .ZN(n442) );
  NOR2_X1 U461 ( .A1(G953), .A2(G237), .ZN(n545) );
  INV_X1 U462 ( .A(KEYINPUT48), .ZN(n595) );
  XNOR2_X1 U463 ( .A(n390), .B(n389), .ZN(n400) );
  INV_X1 U464 ( .A(KEYINPUT105), .ZN(n389) );
  NAND2_X1 U465 ( .A1(n386), .A2(n391), .ZN(n390) );
  NAND2_X1 U466 ( .A1(n385), .A2(n384), .ZN(n379) );
  NOR2_X1 U467 ( .A1(n749), .A2(n397), .ZN(n384) );
  XNOR2_X1 U468 ( .A(n493), .B(n514), .ZN(n544) );
  XNOR2_X1 U469 ( .A(n476), .B(KEYINPUT71), .ZN(n549) );
  INV_X1 U470 ( .A(G137), .ZN(n476) );
  XNOR2_X1 U471 ( .A(n457), .B(G104), .ZN(n456) );
  INV_X1 U472 ( .A(G113), .ZN(n457) );
  XNOR2_X1 U473 ( .A(G143), .B(G122), .ZN(n455) );
  XNOR2_X1 U474 ( .A(n544), .B(n358), .ZN(n731) );
  XNOR2_X1 U475 ( .A(n549), .B(n475), .ZN(n732) );
  INV_X1 U476 ( .A(KEYINPUT97), .ZN(n475) );
  XOR2_X1 U477 ( .A(KEYINPUT95), .B(KEYINPUT17), .Z(n503) );
  XNOR2_X1 U478 ( .A(n492), .B(n501), .ZN(n491) );
  XNOR2_X1 U479 ( .A(n493), .B(n500), .ZN(n492) );
  INV_X1 U480 ( .A(KEYINPUT94), .ZN(n447) );
  NAND2_X1 U481 ( .A1(n664), .A2(n663), .ZN(n615) );
  INV_X1 U482 ( .A(KEYINPUT93), .ZN(n561) );
  NOR2_X1 U483 ( .A1(n574), .A2(n531), .ZN(n558) );
  XNOR2_X1 U484 ( .A(n352), .B(n364), .ZN(n394) );
  INV_X1 U485 ( .A(KEYINPUT5), .ZN(n536) );
  XNOR2_X1 U486 ( .A(G137), .B(G131), .ZN(n537) );
  INV_X1 U487 ( .A(n450), .ZN(n535) );
  INV_X1 U488 ( .A(G146), .ZN(n533) );
  XNOR2_X1 U489 ( .A(n732), .B(n358), .ZN(n551) );
  INV_X1 U490 ( .A(n677), .ZN(n446) );
  XNOR2_X1 U491 ( .A(n471), .B(n470), .ZN(n469) );
  INV_X1 U492 ( .A(KEYINPUT86), .ZN(n470) );
  INV_X1 U493 ( .A(n624), .ZN(n472) );
  XNOR2_X1 U494 ( .A(n572), .B(n571), .ZN(n575) );
  NAND2_X1 U495 ( .A1(n480), .A2(n479), .ZN(n395) );
  AND2_X1 U496 ( .A1(n482), .A2(n481), .ZN(n396) );
  XNOR2_X1 U497 ( .A(n498), .B(KEYINPUT16), .ZN(n499) );
  INV_X1 U498 ( .A(G122), .ZN(n498) );
  XNOR2_X1 U499 ( .A(n736), .B(n410), .ZN(n543) );
  XNOR2_X1 U500 ( .A(n412), .B(n411), .ZN(n410) );
  XNOR2_X1 U501 ( .A(n587), .B(n437), .ZN(n746) );
  XNOR2_X1 U502 ( .A(KEYINPUT42), .B(KEYINPUT110), .ZN(n437) );
  NOR2_X1 U503 ( .A1(n370), .A2(n355), .ZN(n594) );
  NAND2_X1 U504 ( .A1(n444), .A2(n357), .ZN(n443) );
  NOR2_X1 U505 ( .A1(n626), .A2(n625), .ZN(n633) );
  INV_X1 U506 ( .A(KEYINPUT60), .ZN(n422) );
  INV_X1 U507 ( .A(KEYINPUT56), .ZN(n429) );
  AND2_X1 U508 ( .A1(n593), .A2(KEYINPUT36), .ZN(n355) );
  XOR2_X1 U509 ( .A(KEYINPUT13), .B(G475), .Z(n356) );
  XOR2_X1 U510 ( .A(n607), .B(KEYINPUT84), .Z(n357) );
  XNOR2_X1 U511 ( .A(G131), .B(G140), .ZN(n358) );
  XOR2_X1 U512 ( .A(n503), .B(n502), .Z(n359) );
  NOR2_X1 U513 ( .A1(n427), .A2(n658), .ZN(n360) );
  AND2_X1 U514 ( .A1(n575), .A2(n478), .ZN(n361) );
  XOR2_X1 U515 ( .A(KEYINPUT22), .B(KEYINPUT74), .Z(n362) );
  XNOR2_X1 U516 ( .A(KEYINPUT35), .B(KEYINPUT83), .ZN(n363) );
  XOR2_X1 U517 ( .A(n709), .B(n708), .Z(n366) );
  XNOR2_X1 U518 ( .A(n731), .B(n377), .ZN(n710) );
  XOR2_X1 U519 ( .A(n710), .B(n711), .Z(n368) );
  NAND2_X1 U520 ( .A1(n373), .A2(n371), .ZN(n370) );
  NAND2_X1 U521 ( .A1(n418), .A2(KEYINPUT36), .ZN(n372) );
  INV_X1 U522 ( .A(n593), .ZN(n375) );
  INV_X1 U523 ( .A(n612), .ZN(n376) );
  NAND2_X1 U524 ( .A1(n749), .A2(n397), .ZN(n381) );
  NAND2_X1 U525 ( .A1(n392), .A2(n397), .ZN(n383) );
  INV_X1 U526 ( .A(n392), .ZN(n385) );
  INV_X1 U527 ( .A(n409), .ZN(n391) );
  NAND2_X1 U528 ( .A1(n747), .A2(n639), .ZN(n392) );
  XNOR2_X2 U529 ( .A(n576), .B(n581), .ZN(n678) );
  INV_X1 U530 ( .A(KEYINPUT44), .ZN(n397) );
  AND2_X1 U531 ( .A1(n400), .A2(n627), .ZN(n399) );
  XNOR2_X2 U532 ( .A(n532), .B(G134), .ZN(n736) );
  XNOR2_X2 U533 ( .A(G143), .B(G128), .ZN(n532) );
  XNOR2_X2 U534 ( .A(n450), .B(n724), .ZN(n548) );
  NOR2_X2 U535 ( .A1(n721), .A2(n405), .ZN(n629) );
  XNOR2_X1 U536 ( .A(n405), .B(n739), .ZN(n738) );
  XNOR2_X2 U537 ( .A(n406), .B(KEYINPUT103), .ZN(n646) );
  NAND2_X1 U538 ( .A1(n570), .A2(n582), .ZN(n406) );
  XNOR2_X2 U539 ( .A(n407), .B(n356), .ZN(n582) );
  XNOR2_X2 U540 ( .A(n408), .B(n461), .ZN(n570) );
  NOR2_X1 U541 ( .A1(n409), .A2(KEYINPUT47), .ZN(n567) );
  BUF_X1 U542 ( .A(n539), .Z(n415) );
  BUF_X1 U543 ( .A(n715), .Z(n416) );
  OR2_X2 U544 ( .A1(n646), .A2(n650), .ZN(n460) );
  AND2_X1 U545 ( .A1(n558), .A2(n646), .ZN(n465) );
  XNOR2_X1 U546 ( .A(n445), .B(n606), .ZN(n444) );
  BUF_X1 U547 ( .A(n592), .Z(n418) );
  INV_X1 U548 ( .A(n717), .ZN(n486) );
  NAND2_X1 U549 ( .A1(n462), .A2(G472), .ZN(n440) );
  XNOR2_X1 U550 ( .A(n440), .B(n365), .ZN(n419) );
  NAND2_X1 U551 ( .A1(n419), .A2(n486), .ZN(n420) );
  XNOR2_X1 U552 ( .A(n707), .B(n367), .ZN(n435) );
  XNOR2_X1 U553 ( .A(n420), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U554 ( .A(n421), .B(KEYINPUT123), .ZN(G54) );
  NAND2_X1 U555 ( .A1(n424), .A2(n486), .ZN(n421) );
  XNOR2_X1 U556 ( .A(n423), .B(n422), .ZN(G60) );
  NAND2_X1 U557 ( .A1(n425), .A2(n486), .ZN(n423) );
  XNOR2_X1 U558 ( .A(n477), .B(n366), .ZN(n424) );
  XNOR2_X1 U559 ( .A(n712), .B(n368), .ZN(n425) );
  XNOR2_X1 U560 ( .A(n426), .B(n442), .ZN(n441) );
  NOR2_X1 U561 ( .A1(n630), .A2(n631), .ZN(n426) );
  NAND2_X2 U562 ( .A1(n580), .A2(n677), .ZN(n562) );
  NOR2_X1 U563 ( .A1(n750), .A2(n746), .ZN(n590) );
  NOR2_X1 U564 ( .A1(n715), .A2(G902), .ZN(n436) );
  XNOR2_X1 U565 ( .A(n430), .B(n429), .ZN(G51) );
  NAND2_X1 U566 ( .A1(n435), .A2(n486), .ZN(n430) );
  NAND2_X1 U567 ( .A1(n431), .A2(n569), .ZN(n579) );
  NAND2_X1 U568 ( .A1(n568), .A2(n644), .ZN(n431) );
  XNOR2_X1 U569 ( .A(n543), .B(n542), .ZN(n713) );
  XNOR2_X2 U570 ( .A(n726), .B(n548), .ZN(n494) );
  XNOR2_X2 U571 ( .A(G113), .B(KEYINPUT3), .ZN(n496) );
  BUF_X2 U572 ( .A(n629), .Z(n695) );
  XNOR2_X2 U573 ( .A(n438), .B(n497), .ZN(n539) );
  XNOR2_X2 U574 ( .A(n496), .B(G116), .ZN(n438) );
  NOR2_X4 U575 ( .A1(n697), .A2(n441), .ZN(n462) );
  XNOR2_X2 U576 ( .A(n628), .B(KEYINPUT79), .ZN(n697) );
  OR2_X1 U577 ( .A1(n427), .A2(n446), .ZN(n555) );
  XNOR2_X1 U578 ( .A(n350), .B(n447), .ZN(n612) );
  NAND2_X1 U579 ( .A1(n622), .A2(n448), .ZN(n626) );
  INV_X1 U580 ( .A(n427), .ZN(n448) );
  XNOR2_X1 U581 ( .A(n449), .B(n552), .ZN(n709) );
  INV_X1 U582 ( .A(n566), .ZN(n679) );
  XNOR2_X2 U583 ( .A(n460), .B(KEYINPUT104), .ZN(n566) );
  NAND2_X1 U584 ( .A1(n462), .A2(G210), .ZN(n707) );
  NAND2_X1 U585 ( .A1(n462), .A2(G469), .ZN(n477) );
  NAND2_X1 U586 ( .A1(n462), .A2(G475), .ZN(n712) );
  NAND2_X1 U587 ( .A1(n462), .A2(G478), .ZN(n489) );
  NAND2_X1 U588 ( .A1(n462), .A2(G217), .ZN(n714) );
  XNOR2_X1 U589 ( .A(n468), .B(n466), .ZN(n632) );
  XNOR2_X1 U590 ( .A(n535), .B(n467), .ZN(n466) );
  XNOR2_X1 U591 ( .A(n538), .B(n534), .ZN(n467) );
  XNOR2_X1 U592 ( .A(n415), .B(n547), .ZN(n468) );
  NOR2_X1 U593 ( .A1(n709), .A2(G902), .ZN(n553) );
  NAND2_X1 U594 ( .A1(n473), .A2(n472), .ZN(n471) );
  XNOR2_X1 U595 ( .A(n613), .B(KEYINPUT106), .ZN(n473) );
  XNOR2_X2 U596 ( .A(n553), .B(n474), .ZN(n573) );
  NOR2_X1 U597 ( .A1(n574), .A2(n483), .ZN(n479) );
  INV_X1 U598 ( .A(n618), .ZN(n480) );
  NAND2_X1 U599 ( .A1(n618), .A2(n483), .ZN(n482) );
  INV_X1 U600 ( .A(KEYINPUT80), .ZN(n483) );
  XNOR2_X2 U601 ( .A(n484), .B(G146), .ZN(n493) );
  XNOR2_X1 U602 ( .A(n485), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U603 ( .A1(n487), .A2(n486), .ZN(n485) );
  XNOR2_X1 U604 ( .A(n489), .B(n488), .ZN(n487) );
  INV_X1 U605 ( .A(n713), .ZN(n488) );
  XNOR2_X2 U606 ( .A(n494), .B(n490), .ZN(n704) );
  XNOR2_X2 U607 ( .A(n539), .B(n499), .ZN(n726) );
  XNOR2_X1 U608 ( .A(n521), .B(n495), .ZN(n522) );
  XNOR2_X2 U609 ( .A(n588), .B(KEYINPUT40), .ZN(n750) );
  BUF_X1 U610 ( .A(n580), .Z(n576) );
  NOR2_X2 U611 ( .A1(n609), .A2(n623), .ZN(n664) );
  XOR2_X1 U612 ( .A(n520), .B(n519), .Z(n495) );
  XNOR2_X1 U613 ( .A(KEYINPUT92), .B(KEYINPUT46), .ZN(n589) );
  XNOR2_X1 U614 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U615 ( .A(KEYINPUT30), .B(KEYINPUT109), .ZN(n571) );
  XNOR2_X1 U616 ( .A(n523), .B(n522), .ZN(n715) );
  NOR2_X1 U617 ( .A1(G952), .A2(n737), .ZN(n717) );
  INV_X1 U618 ( .A(n532), .ZN(n500) );
  XOR2_X1 U619 ( .A(KEYINPUT82), .B(KEYINPUT18), .Z(n501) );
  NAND2_X1 U620 ( .A1(G224), .A2(n737), .ZN(n502) );
  NOR2_X2 U621 ( .A1(n704), .A2(n524), .ZN(n506) );
  XNOR2_X1 U622 ( .A(n504), .B(KEYINPUT77), .ZN(n554) );
  NAND2_X1 U623 ( .A1(G210), .A2(n554), .ZN(n505) );
  XNOR2_X2 U624 ( .A(n506), .B(n505), .ZN(n580) );
  NOR2_X1 U625 ( .A1(G900), .A2(n737), .ZN(n507) );
  NAND2_X1 U626 ( .A1(n507), .A2(G902), .ZN(n508) );
  NAND2_X1 U627 ( .A1(G952), .A2(n737), .ZN(n598) );
  NAND2_X1 U628 ( .A1(n508), .A2(n598), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n509), .B(KEYINPUT14), .ZN(n600) );
  NAND2_X1 U630 ( .A1(n510), .A2(n600), .ZN(n574) );
  XOR2_X1 U631 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n512) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(KEYINPUT98), .ZN(n511) );
  XNOR2_X1 U633 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U634 ( .A(KEYINPUT23), .B(n513), .Z(n516) );
  XNOR2_X1 U635 ( .A(KEYINPUT10), .B(KEYINPUT70), .ZN(n514) );
  XNOR2_X1 U636 ( .A(n549), .B(n544), .ZN(n515) );
  XNOR2_X1 U637 ( .A(n515), .B(n516), .ZN(n523) );
  XOR2_X1 U638 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n518) );
  NAND2_X1 U639 ( .A1(G234), .A2(n737), .ZN(n517) );
  NAND2_X1 U640 ( .A1(G221), .A2(n541), .ZN(n521) );
  XOR2_X1 U641 ( .A(G140), .B(G119), .Z(n520) );
  BUF_X1 U642 ( .A(G128), .Z(n643) );
  XNOR2_X1 U643 ( .A(n643), .B(G110), .ZN(n519) );
  INV_X1 U644 ( .A(n524), .ZN(n631) );
  NAND2_X1 U645 ( .A1(G234), .A2(n631), .ZN(n525) );
  XNOR2_X1 U646 ( .A(KEYINPUT20), .B(n525), .ZN(n529) );
  NAND2_X1 U647 ( .A1(G217), .A2(n529), .ZN(n527) );
  NAND2_X1 U648 ( .A1(n529), .A2(G221), .ZN(n530) );
  XOR2_X1 U649 ( .A(KEYINPUT21), .B(n530), .Z(n659) );
  NAND2_X1 U650 ( .A1(n623), .A2(n659), .ZN(n531) );
  AND2_X1 U651 ( .A1(n545), .A2(G210), .ZN(n534) );
  NAND2_X1 U652 ( .A1(n541), .A2(G217), .ZN(n542) );
  NAND2_X1 U653 ( .A1(n545), .A2(G214), .ZN(n546) );
  NAND2_X1 U654 ( .A1(G227), .A2(n737), .ZN(n550) );
  XNOR2_X1 U655 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U656 ( .A1(n593), .A2(n555), .ZN(n556) );
  XNOR2_X1 U657 ( .A(n556), .B(KEYINPUT43), .ZN(n557) );
  NOR2_X1 U658 ( .A1(n576), .A2(n557), .ZN(n656) );
  NOR2_X1 U659 ( .A1(n582), .A2(n570), .ZN(n650) );
  XNOR2_X1 U660 ( .A(KEYINPUT28), .B(n559), .ZN(n560) );
  NAND2_X1 U661 ( .A1(n560), .A2(n573), .ZN(n586) );
  XNOR2_X2 U662 ( .A(n562), .B(n561), .ZN(n592) );
  XOR2_X1 U663 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n563) );
  INV_X1 U664 ( .A(n351), .ZN(n564) );
  NAND2_X1 U665 ( .A1(n566), .A2(n644), .ZN(n565) );
  NAND2_X1 U666 ( .A1(n565), .A2(KEYINPUT47), .ZN(n569) );
  XNOR2_X1 U667 ( .A(n567), .B(KEYINPUT76), .ZN(n568) );
  INV_X1 U668 ( .A(n570), .ZN(n583) );
  NAND2_X1 U669 ( .A1(n583), .A2(n582), .ZN(n607) );
  NAND2_X1 U670 ( .A1(n617), .A2(n677), .ZN(n572) );
  INV_X1 U671 ( .A(n659), .ZN(n609) );
  NAND2_X1 U672 ( .A1(n573), .A2(n664), .ZN(n618) );
  NAND2_X1 U673 ( .A1(n576), .A2(n361), .ZN(n577) );
  XOR2_X1 U674 ( .A(KEYINPUT89), .B(n417), .Z(n578) );
  INV_X1 U675 ( .A(KEYINPUT38), .ZN(n581) );
  NOR2_X1 U676 ( .A1(n583), .A2(n582), .ZN(n608) );
  AND2_X1 U677 ( .A1(n677), .A2(n608), .ZN(n584) );
  AND2_X1 U678 ( .A1(n678), .A2(n584), .ZN(n585) );
  NOR2_X1 U679 ( .A1(n586), .A2(n674), .ZN(n587) );
  XNOR2_X1 U680 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U681 ( .A(KEYINPUT111), .B(n594), .ZN(n745) );
  NAND2_X1 U682 ( .A1(n596), .A2(n650), .ZN(n655) );
  NOR2_X1 U683 ( .A1(G898), .A2(n737), .ZN(n597) );
  XNOR2_X1 U684 ( .A(KEYINPUT96), .B(n597), .ZN(n728) );
  NAND2_X1 U685 ( .A1(n728), .A2(G902), .ZN(n599) );
  AND2_X1 U686 ( .A1(n599), .A2(n598), .ZN(n601) );
  INV_X1 U687 ( .A(n600), .ZN(n690) );
  NOR2_X1 U688 ( .A1(n601), .A2(n690), .ZN(n602) );
  XNOR2_X1 U689 ( .A(n615), .B(KEYINPUT107), .ZN(n604) );
  NAND2_X1 U690 ( .A1(n604), .A2(n624), .ZN(n605) );
  XNOR2_X1 U691 ( .A(n605), .B(KEYINPUT33), .ZN(n657) );
  INV_X1 U692 ( .A(KEYINPUT34), .ZN(n606) );
  INV_X1 U693 ( .A(n608), .ZN(n676) );
  NOR2_X1 U694 ( .A1(n609), .A2(n676), .ZN(n610) );
  INV_X1 U695 ( .A(n623), .ZN(n658) );
  AND2_X1 U696 ( .A1(n621), .A2(n360), .ZN(n611) );
  INV_X1 U697 ( .A(n617), .ZN(n662) );
  NAND2_X1 U698 ( .A1(n611), .A2(n662), .ZN(n639) );
  NOR2_X1 U699 ( .A1(n658), .A2(n612), .ZN(n613) );
  XOR2_X1 U700 ( .A(KEYINPUT85), .B(KEYINPUT32), .Z(n614) );
  NOR2_X1 U701 ( .A1(n662), .A2(n615), .ZN(n670) );
  NAND2_X1 U702 ( .A1(n394), .A2(n670), .ZN(n616) );
  NOR2_X1 U703 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n394), .A2(n619), .ZN(n620) );
  BUF_X1 U705 ( .A(n621), .Z(n622) );
  OR2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U707 ( .A(n633), .ZN(n627) );
  NAND2_X1 U708 ( .A1(KEYINPUT2), .A2(n695), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(KEYINPUT2), .ZN(n630) );
  XOR2_X1 U710 ( .A(G101), .B(n633), .Z(G3) );
  NAND2_X1 U711 ( .A1(n635), .A2(n646), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(G104), .ZN(G6) );
  XOR2_X1 U713 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n637) );
  NAND2_X1 U714 ( .A1(n635), .A2(n650), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U716 ( .A(G107), .B(n638), .ZN(G9) );
  XNOR2_X1 U717 ( .A(n639), .B(G110), .ZN(G12) );
  XOR2_X1 U718 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n641) );
  NAND2_X1 U719 ( .A1(n644), .A2(n650), .ZN(n640) );
  XNOR2_X1 U720 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n643), .B(n642), .ZN(G30) );
  XOR2_X1 U722 ( .A(n417), .B(G143), .Z(G45) );
  NAND2_X1 U723 ( .A1(n644), .A2(n646), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n645), .B(G146), .ZN(G48) );
  XOR2_X1 U725 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n648) );
  NAND2_X1 U726 ( .A1(n651), .A2(n646), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(G113), .B(n649), .ZN(G15) );
  XOR2_X1 U729 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n653) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U732 ( .A(G116), .B(n654), .ZN(G18) );
  XNOR2_X1 U733 ( .A(G134), .B(n655), .ZN(G36) );
  XOR2_X1 U734 ( .A(G140), .B(n656), .Z(G42) );
  INV_X1 U735 ( .A(n657), .ZN(n684) );
  OR2_X1 U736 ( .A1(n684), .A2(n674), .ZN(n701) );
  NOR2_X1 U737 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n660), .B(KEYINPUT49), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n664), .A2(n427), .ZN(n665) );
  XNOR2_X1 U741 ( .A(n665), .B(KEYINPUT50), .ZN(n666) );
  NOR2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U743 ( .A(KEYINPUT117), .B(n668), .Z(n669) );
  NOR2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U745 ( .A(KEYINPUT51), .B(n671), .Z(n672) );
  XNOR2_X1 U746 ( .A(n672), .B(KEYINPUT118), .ZN(n673) );
  NOR2_X1 U747 ( .A1(n674), .A2(n673), .ZN(n687) );
  NOR2_X1 U748 ( .A1(n678), .A2(n677), .ZN(n675) );
  NOR2_X1 U749 ( .A1(n676), .A2(n675), .ZN(n683) );
  NAND2_X1 U750 ( .A1(n678), .A2(n677), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U752 ( .A(KEYINPUT119), .B(n681), .Z(n682) );
  NOR2_X1 U753 ( .A1(n683), .A2(n682), .ZN(n685) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U756 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U758 ( .A1(n691), .A2(G952), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT120), .ZN(n693) );
  NAND2_X1 U760 ( .A1(n693), .A2(n737), .ZN(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT2), .B(KEYINPUT87), .Z(n694) );
  NOR2_X1 U762 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U766 ( .A(n702), .B(KEYINPUT121), .ZN(n703) );
  XNOR2_X1 U767 ( .A(KEYINPUT53), .B(n703), .ZN(G75) );
  XOR2_X1 U768 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n706) );
  XNOR2_X1 U769 ( .A(n704), .B(KEYINPUT55), .ZN(n705) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n708) );
  XOR2_X1 U771 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n711) );
  XNOR2_X1 U772 ( .A(n416), .B(n714), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n717), .A2(n716), .ZN(G66) );
  NAND2_X1 U774 ( .A1(G224), .A2(G953), .ZN(n718) );
  XNOR2_X1 U775 ( .A(n718), .B(KEYINPUT126), .ZN(n719) );
  XNOR2_X1 U776 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  AND2_X1 U777 ( .A1(n720), .A2(G898), .ZN(n723) );
  NOR2_X1 U778 ( .A1(G953), .A2(n721), .ZN(n722) );
  NOR2_X1 U779 ( .A1(n723), .A2(n722), .ZN(n730) );
  XOR2_X1 U780 ( .A(G101), .B(n724), .Z(n725) );
  XNOR2_X1 U781 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U782 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U783 ( .A(n730), .B(n729), .Z(G69) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n734) );
  XNOR2_X1 U785 ( .A(n733), .B(n734), .ZN(n735) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(n739) );
  NAND2_X1 U787 ( .A1(n738), .A2(n737), .ZN(n743) );
  XNOR2_X1 U788 ( .A(G227), .B(n739), .ZN(n740) );
  NAND2_X1 U789 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n741), .A2(G953), .ZN(n742) );
  NAND2_X1 U791 ( .A1(n743), .A2(n742), .ZN(G72) );
  XOR2_X1 U792 ( .A(G125), .B(KEYINPUT37), .Z(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(G27) );
  XOR2_X1 U794 ( .A(G137), .B(n746), .Z(G39) );
  XNOR2_X1 U795 ( .A(G122), .B(n748), .ZN(G24) );
  XOR2_X1 U796 ( .A(n749), .B(G119), .Z(G21) );
  XOR2_X1 U797 ( .A(n750), .B(G131), .Z(G33) );
endmodule

