//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n451), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OR2_X1    g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT68), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(new_n463), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n474), .B1(new_n469), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n465), .A2(G2104), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n476), .A2(G2105), .B1(G101), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n473), .A2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n470), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n469), .A2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g059(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G112), .B2(new_n465), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n480), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  OAI22_X1  g065(.A1(new_n466), .A2(new_n489), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n491));
  XOR2_X1   g066(.A(KEYINPUT70), .B(KEYINPUT4), .Z(new_n492));
  NAND3_X1  g067(.A1(new_n470), .A2(G138), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n465), .A2(G114), .ZN(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n481), .B2(G126), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT6), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT71), .B1(new_n503), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(new_n501), .A3(KEYINPUT6), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(G50), .A3(G543), .ZN(new_n508));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(G88), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  AND2_X1   g089(.A1(G75), .A2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(G651), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n508), .A2(new_n512), .A3(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  AOI21_X1  g093(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n522), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n519), .A2(G63), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n504), .A2(new_n506), .ZN(new_n525));
  INV_X1    g100(.A(new_n502), .ZN(new_n526));
  NAND4_X1  g101(.A1(new_n525), .A2(G89), .A3(new_n526), .A4(new_n511), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n525), .A2(G51), .A3(G543), .A4(new_n526), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n501), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT72), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n507), .A2(G52), .A3(G543), .ZN(new_n533));
  INV_X1    g108(.A(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n507), .A2(new_n511), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n509), .B2(new_n510), .ZN(new_n539));
  AND2_X1   g114(.A1(G68), .A2(G543), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n525), .A2(G43), .A3(G543), .A4(new_n526), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n541), .B(new_n542), .C1(new_n535), .C2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  AND2_X1   g126(.A1(G53), .A2(G543), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n525), .A2(KEYINPUT75), .A3(new_n526), .A4(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(KEYINPUT74), .A2(KEYINPUT75), .A3(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n507), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n525), .A2(new_n526), .A3(new_n552), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n555), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n555), .A2(new_n560), .A3(KEYINPUT76), .A4(new_n557), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n507), .A2(G91), .A3(new_n511), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n509), .A2(KEYINPUT77), .A3(new_n510), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  AND2_X1   g143(.A1(KEYINPUT5), .A2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(KEYINPUT5), .A2(G543), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n566), .B1(new_n573), .B2(new_n501), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT78), .B1(new_n565), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  AOI211_X1 g152(.A(new_n577), .B(new_n574), .C1(new_n563), .C2(new_n564), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  NAND3_X1  g155(.A1(new_n524), .A2(new_n527), .A3(new_n528), .ZN(G286));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  OAI211_X1 g157(.A(new_n582), .B(G651), .C1(new_n511), .C2(G74), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n569), .B2(new_n570), .ZN(new_n584));
  NAND2_X1  g159(.A1(G74), .A2(G651), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(KEYINPUT79), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n507), .A2(G49), .A3(G543), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n507), .A2(G87), .A3(new_n511), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  NAND3_X1  g165(.A1(new_n507), .A2(G48), .A3(G543), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n507), .A2(G86), .A3(new_n511), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n509), .B2(new_n510), .ZN(new_n594));
  AND2_X1   g169(.A1(G73), .A2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n591), .A2(new_n592), .A3(new_n596), .ZN(G305));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n509), .B2(new_n510), .ZN(new_n599));
  AND2_X1   g174(.A1(G72), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n525), .A2(G85), .A3(new_n526), .A4(new_n511), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n525), .A2(G47), .A3(G543), .A4(new_n526), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n567), .B2(new_n571), .ZN(new_n607));
  AND2_X1   g182(.A1(G79), .A2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n507), .A2(G54), .A3(G543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n609), .A2(KEYINPUT80), .A3(new_n610), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g190(.A1(new_n507), .A2(G92), .A3(new_n511), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(KEYINPUT10), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n613), .A2(new_n614), .B1(new_n617), .B2(new_n618), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n605), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n605), .B1(new_n626), .B2(G868), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT82), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n626), .B1(new_n634), .B2(G860), .ZN(G148));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n544), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n625), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n636), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n464), .A2(new_n477), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n470), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n481), .A2(G123), .ZN(new_n646));
  OR2_X1    g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n647), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT83), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n651), .ZN(G156));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2430), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n659));
  OAI22_X1  g234(.A1(new_n658), .A2(new_n659), .B1(new_n654), .B2(new_n655), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2451), .B(G2454), .Z(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2443), .B(G2446), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(G401));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT86), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n676), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2072), .B(G2078), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n677), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n681), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1961), .B(G1966), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT20), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n689), .A2(new_n690), .ZN(new_n694));
  NOR3_X1   g269(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(new_n688), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(G229));
  NAND2_X1  g278(.A1(new_n470), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n481), .A2(G119), .ZN(new_n705));
  OR2_X1    g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT89), .B(G29), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G25), .B(new_n708), .S(new_n710), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G16), .A2(G24), .ZN(new_n715));
  AND3_X1   g290(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G16), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1986), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G23), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT92), .ZN(new_n722));
  NAND2_X1  g297(.A1(G288), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n587), .A2(KEYINPUT92), .A3(new_n588), .A4(new_n589), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(new_n720), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT93), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT33), .B(G1976), .Z(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(KEYINPUT93), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n720), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n720), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1971), .ZN(new_n735));
  NOR2_X1   g310(.A1(G6), .A2(G16), .ZN(new_n736));
  INV_X1    g311(.A(G305), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G16), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT32), .B(G1981), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n735), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n732), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n730), .B1(new_n728), .B2(new_n731), .ZN(new_n744));
  OR3_X1    g319(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n748));
  AOI21_X1  g323(.A(new_n719), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n748), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n745), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT36), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n749), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n720), .A2(G4), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n625), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT95), .B(G1348), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n720), .A2(G19), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n545), .B2(new_n720), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1341), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n470), .A2(G140), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n481), .A2(G128), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n465), .A2(G116), .ZN(new_n766));
  OAI21_X1  g341(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G29), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n709), .A2(G26), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2067), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n759), .A2(new_n760), .A3(new_n763), .A4(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n720), .A2(G20), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT101), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G299), .B2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n710), .A2(G35), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G162), .B2(new_n710), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT29), .Z(new_n786));
  INV_X1    g361(.A(G2090), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n470), .A2(G141), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n481), .A2(G129), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n477), .A2(G105), .ZN(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT26), .Z(new_n793));
  NAND4_X1  g368(.A1(new_n789), .A2(new_n790), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G32), .B(new_n794), .S(G29), .Z(new_n795));
  XOR2_X1   g370(.A(KEYINPUT27), .B(G1996), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT99), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n795), .B(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n649), .A2(new_n709), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT31), .B(G11), .Z(new_n800));
  INV_X1    g375(.A(G29), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(G28), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT100), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n803), .A2(KEYINPUT100), .B1(new_n802), .B2(G28), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n788), .A2(new_n798), .A3(new_n799), .A4(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT24), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(G34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(G34), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n709), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G160), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n801), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2084), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n709), .A2(G27), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G164), .B2(new_n709), .ZN(new_n816));
  INV_X1    g391(.A(G2078), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n807), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(G171), .A2(new_n720), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G5), .B2(new_n720), .ZN(new_n822));
  INV_X1    g397(.A(G1961), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n465), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  NAND3_X1  g402(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT25), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G139), .B2(new_n470), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT97), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G29), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n801), .A2(G33), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(G2072), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(G2072), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n824), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n822), .A2(new_n823), .B1(new_n786), .B2(new_n787), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n720), .A2(G21), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G168), .B2(new_n720), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(G1966), .ZN(new_n842));
  AND2_X1   g417(.A1(new_n841), .A2(G1966), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AND4_X1   g419(.A1(new_n783), .A2(new_n820), .A3(new_n838), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n777), .A2(new_n778), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT102), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n777), .A2(new_n848), .A3(new_n778), .A4(new_n845), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n753), .A2(new_n755), .B1(new_n847), .B2(new_n849), .ZN(G311));
  NAND2_X1  g425(.A1(new_n753), .A2(new_n755), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(G150));
  NAND2_X1  g428(.A1(new_n626), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n509), .B2(new_n510), .ZN(new_n857));
  AND2_X1   g432(.A1(G80), .A2(G543), .ZN(new_n858));
  OAI21_X1  g433(.A(G651), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT103), .B(G55), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n525), .A2(G543), .A3(new_n526), .A4(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G93), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n861), .C1(new_n535), .C2(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n544), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n544), .A2(new_n863), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n855), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  AOI21_X1  g444(.A(G860), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n863), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT37), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(G145));
  XOR2_X1   g449(.A(new_n708), .B(KEYINPUT106), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n642), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n768), .B(KEYINPUT105), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n832), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n832), .A2(new_n878), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n876), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n491), .A2(new_n885), .A3(new_n493), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n885), .B1(new_n491), .B2(new_n493), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n498), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n794), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n470), .A2(G142), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n481), .A2(G130), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n465), .A2(G118), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n889), .A2(new_n894), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n884), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n881), .A2(new_n895), .A3(new_n883), .A4(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n487), .B(new_n649), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n812), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n904), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n905), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n908), .A2(KEYINPUT40), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT40), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(G395));
  NAND2_X1  g487(.A1(new_n638), .A2(new_n867), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n866), .B1(new_n625), .B2(G559), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n620), .B1(new_n576), .B2(new_n578), .ZN(new_n916));
  AND4_X1   g491(.A1(new_n525), .A2(new_n526), .A3(new_n552), .A4(new_n556), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT74), .B1(new_n507), .B2(new_n552), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT76), .B1(new_n919), .B2(new_n555), .ZN(new_n920));
  AND4_X1   g495(.A1(KEYINPUT76), .A2(new_n555), .A3(new_n557), .A4(new_n560), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n575), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n577), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n565), .A2(KEYINPUT78), .A3(new_n575), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n622), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT41), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n916), .A2(new_n925), .A3(KEYINPUT41), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n915), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n916), .A2(new_n925), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n928), .B(KEYINPUT108), .C1(new_n915), .C2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  NAND2_X1  g507(.A1(G290), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n716), .A2(KEYINPUT109), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n725), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n933), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n723), .A3(new_n724), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(G303), .A2(G305), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(G303), .A2(G305), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(KEYINPUT110), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  INV_X1    g518(.A(new_n941), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n943), .B1(new_n944), .B2(new_n939), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n944), .A2(new_n939), .A3(new_n943), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n935), .A2(new_n947), .A3(new_n937), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n949), .A2(KEYINPUT111), .A3(KEYINPUT112), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n725), .B(new_n936), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n942), .A2(new_n945), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n951), .B(new_n948), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT42), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT42), .B1(new_n949), .B2(KEYINPUT112), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OR3_X1    g536(.A1(new_n915), .A2(KEYINPUT108), .A3(new_n930), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n956), .A2(KEYINPUT113), .A3(new_n958), .ZN(new_n963));
  AND4_X1   g538(.A1(new_n931), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n963), .A2(new_n961), .B1(new_n931), .B2(new_n962), .ZN(new_n965));
  OAI21_X1  g540(.A(G868), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n863), .A2(new_n636), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(G295));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n967), .ZN(G331));
  INV_X1    g544(.A(KEYINPUT117), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT114), .B(KEYINPUT44), .Z(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n951), .B1(new_n946), .B2(new_n948), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n955), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G168), .A2(KEYINPUT115), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n976));
  NAND2_X1  g551(.A1(G286), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n544), .A2(new_n863), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n544), .A2(new_n863), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n977), .B(new_n975), .C1(new_n864), .C2(new_n865), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G301), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n981), .A2(new_n982), .A3(G171), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n929), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT41), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n576), .A2(new_n578), .A3(new_n620), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n622), .B1(new_n923), .B2(new_n924), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n916), .A2(new_n925), .A3(KEYINPUT41), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n986), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n993), .B2(KEYINPUT116), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n984), .A2(new_n985), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n927), .B2(new_n926), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n974), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n930), .A2(new_n995), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n993), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n955), .A2(new_n973), .ZN(new_n1003));
  AOI21_X1  g578(.A(G37), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1000), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n974), .B1(new_n993), .B2(new_n1001), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n996), .A2(new_n1003), .A3(new_n987), .ZN(new_n1008));
  INV_X1    g583(.A(G37), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT43), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n972), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1000), .B1(new_n999), .B2(new_n1004), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1006), .A2(new_n1008), .A3(new_n1000), .A4(new_n1009), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT44), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n970), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1001), .B1(new_n996), .B2(new_n997), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n993), .A2(KEYINPUT116), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1003), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n1020), .A2(KEYINPUT43), .A3(new_n1010), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1000), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n971), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT43), .B1(new_n1020), .B2(new_n1010), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(KEYINPUT44), .A3(new_n1014), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1023), .A2(KEYINPUT117), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1017), .A2(new_n1026), .ZN(G397));
  NOR2_X1   g602(.A1(new_n622), .A2(KEYINPUT125), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n473), .A2(G40), .A3(new_n478), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n888), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n773), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n888), .A2(new_n1035), .A3(new_n1029), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n499), .A2(new_n1029), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1030), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n758), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1034), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT60), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1028), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1044), .A2(new_n758), .B1(new_n1033), .B2(new_n773), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n620), .B(KEYINPUT125), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(KEYINPUT60), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1043), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n922), .A2(KEYINPUT57), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n574), .A2(new_n561), .A3(KEYINPUT57), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1956), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1035), .B1(new_n888), .B2(new_n1029), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1031), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT45), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1030), .B1(new_n1037), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1053), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1053), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(KEYINPUT61), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1996), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1058), .A2(new_n1060), .A3(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  NAND2_X1  g644(.A1(new_n1032), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n544), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n1071), .B(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT61), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1065), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1075), .B1(new_n1076), .B2(new_n1063), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1049), .A2(new_n1066), .A3(new_n1074), .A4(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1045), .A2(new_n620), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1065), .B1(new_n1079), .B2(new_n1063), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1058), .A2(new_n1060), .A3(new_n817), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n888), .A2(new_n1029), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1059), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n1029), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1084), .A2(G2078), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1087), .A2(new_n1031), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1044), .A2(new_n823), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G171), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT127), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT127), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1092), .A2(new_n1095), .A3(G171), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1087), .A2(new_n1031), .A3(new_n1058), .A4(new_n1089), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1085), .A2(new_n1098), .A3(new_n1091), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1082), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1087), .A2(new_n1031), .A3(new_n1088), .ZN(new_n1102));
  INV_X1    g677(.A(G1966), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1044), .A2(G2084), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(G168), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(KEYINPUT126), .A2(KEYINPUT51), .ZN(new_n1107));
  OR2_X1    g682(.A1(KEYINPUT126), .A2(KEYINPUT51), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1106), .A2(G8), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G2084), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1102), .A2(new_n1103), .B1(new_n1039), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1112), .A2(G8), .A3(G286), .ZN(new_n1113));
  INV_X1    g688(.A(G8), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1111), .B2(G168), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1109), .B(new_n1113), .C1(new_n1115), .C2(new_n1107), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n726), .A2(G1976), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1032), .A2(new_n1117), .A3(new_n1118), .A4(G8), .ZN(new_n1119));
  INV_X1    g694(.A(G288), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(G1976), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1117), .A2(new_n1032), .A3(G8), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(G305), .B(G1981), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT49), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n1127), .B(KEYINPUT122), .Z(new_n1128));
  NAND2_X1  g703(.A1(new_n1032), .A2(G8), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1119), .A2(new_n1124), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1055), .A2(new_n1056), .A3(G2090), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1971), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1134));
  OAI21_X1  g709(.A(G8), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(G303), .A2(G8), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT55), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1124), .A2(new_n1119), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1137), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1044), .A2(G2090), .ZN(new_n1141));
  OAI211_X1 g716(.A(G8), .B(new_n1140), .C1(new_n1141), .C2(new_n1134), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1132), .A2(new_n1138), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1085), .A2(new_n1090), .A3(new_n1091), .A4(G301), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1082), .B1(new_n1099), .B2(G171), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1081), .A2(new_n1101), .A3(new_n1116), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1116), .A2(KEYINPUT62), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1143), .B1(new_n1096), .B2(new_n1094), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1106), .A2(G8), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(KEYINPUT126), .A3(KEYINPUT51), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1151), .A2(new_n1152), .A3(new_n1109), .A4(new_n1113), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1148), .A2(new_n1149), .A3(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1129), .B(KEYINPUT123), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1156));
  INV_X1    g731(.A(G1976), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1120), .ZN(new_n1158));
  OR2_X1    g733(.A1(G305), .A2(G1981), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1155), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1142), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1132), .A2(new_n1139), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1111), .A2(new_n1114), .A3(G286), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1143), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(G8), .B1(new_n1141), .B2(new_n1134), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1168), .B2(new_n1137), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1162), .A2(new_n1142), .A3(new_n1165), .A4(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1147), .A2(new_n1154), .A3(new_n1163), .A4(new_n1171), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n1087), .A2(KEYINPUT118), .A3(new_n1030), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT118), .B1(new_n1087), .B2(new_n1030), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(G290), .A2(G1986), .ZN(new_n1177));
  AND2_X1   g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT119), .Z(new_n1180));
  XNOR2_X1  g755(.A(new_n768), .B(G2067), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1176), .A2(KEYINPUT120), .A3(new_n1181), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n794), .B(G1996), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1184), .A2(new_n1185), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n713), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n708), .A2(new_n1188), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n708), .A2(new_n1188), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1176), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g766(.A1(new_n1180), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1172), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT48), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1187), .A2(new_n1195), .A3(new_n1191), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT46), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1176), .A2(new_n1197), .A3(new_n1067), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT46), .B1(new_n1175), .B2(G1996), .ZN(new_n1199));
  OR2_X1    g774(.A1(new_n1181), .A2(new_n794), .ZN(new_n1200));
  AOI22_X1  g775(.A1(new_n1198), .A2(new_n1199), .B1(new_n1176), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT47), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1196), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n768), .A2(G2067), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1175), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NOR2_X1   g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1193), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g785(.A(G319), .ZN(new_n1212));
  OR2_X1    g786(.A1(G227), .A2(new_n1212), .ZN(new_n1213));
  NOR3_X1   g787(.A1(G401), .A2(G229), .A3(new_n1213), .ZN(new_n1214));
  AND3_X1   g788(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n905), .ZN(new_n1215));
  AOI21_X1  g789(.A(KEYINPUT107), .B1(new_n903), .B2(new_n905), .ZN(new_n1216));
  OAI221_X1 g790(.A(new_n1214), .B1(new_n1021), .B2(new_n1022), .C1(new_n1215), .C2(new_n1216), .ZN(G225));
  INV_X1    g791(.A(G225), .ZN(G308));
endmodule


