

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755;

  XNOR2_X1 U379 ( .A(n417), .B(n367), .ZN(n570) );
  XNOR2_X2 U380 ( .A(n547), .B(n428), .ZN(n561) );
  NAND2_X2 U381 ( .A1(n406), .A2(n402), .ZN(n383) );
  NOR2_X1 U382 ( .A1(n398), .A2(n585), .ZN(n586) );
  XNOR2_X1 U383 ( .A(n372), .B(n551), .ZN(n398) );
  NAND2_X1 U384 ( .A1(n550), .A2(n685), .ZN(n372) );
  INV_X1 U385 ( .A(G146), .ZN(n409) );
  BUF_X1 U386 ( .A(n751), .Z(n358) );
  XNOR2_X1 U387 ( .A(n424), .B(n366), .ZN(n751) );
  XNOR2_X1 U388 ( .A(n738), .B(n409), .ZN(n479) );
  NOR2_X1 U389 ( .A1(n665), .A2(n626), .ZN(n456) );
  XNOR2_X1 U390 ( .A(n625), .B(n369), .ZN(n665) );
  NAND2_X1 U391 ( .A1(n751), .A2(KEYINPUT44), .ZN(n592) );
  AND2_X1 U392 ( .A1(n433), .A2(n438), .ZN(n437) );
  AND2_X1 U393 ( .A1(n615), .A2(n599), .ZN(n610) );
  XNOR2_X1 U394 ( .A(n450), .B(n477), .ZN(n382) );
  XNOR2_X1 U395 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U396 ( .A1(n627), .A2(KEYINPUT2), .ZN(n458) );
  INV_X1 U397 ( .A(n472), .ZN(n531) );
  XNOR2_X1 U398 ( .A(KEYINPUT4), .B(G131), .ZN(n476) );
  INV_X2 U399 ( .A(G953), .ZN(n745) );
  BUF_X1 U400 ( .A(n397), .Z(n359) );
  XNOR2_X2 U401 ( .A(G101), .B(G104), .ZN(n399) );
  XNOR2_X2 U402 ( .A(n401), .B(G110), .ZN(n400) );
  INV_X2 U403 ( .A(KEYINPUT74), .ZN(n401) );
  XNOR2_X2 U404 ( .A(n540), .B(n539), .ZN(n550) );
  XNOR2_X2 U405 ( .A(n400), .B(n399), .ZN(n534) );
  NOR2_X1 U406 ( .A1(n655), .A2(n657), .ZN(n691) );
  NAND2_X1 U407 ( .A1(n373), .A2(n476), .ZN(n376) );
  AND2_X1 U408 ( .A1(n475), .A2(n377), .ZN(n375) );
  AND2_X1 U409 ( .A1(n587), .A2(KEYINPUT33), .ZN(n445) );
  OR2_X1 U410 ( .A1(G237), .A2(G902), .ZN(n537) );
  XNOR2_X1 U411 ( .A(n501), .B(G475), .ZN(n502) );
  NAND2_X1 U412 ( .A1(n381), .A2(n404), .ZN(n449) );
  INV_X1 U413 ( .A(n382), .ZN(n381) );
  INV_X1 U414 ( .A(KEYINPUT84), .ZN(n465) );
  XNOR2_X1 U415 ( .A(G902), .B(KEYINPUT15), .ZN(n626) );
  INV_X1 U416 ( .A(G472), .ZN(n405) );
  NAND2_X1 U417 ( .A1(G902), .A2(G472), .ZN(n407) );
  XNOR2_X1 U418 ( .A(n409), .B(n392), .ZN(n391) );
  INV_X1 U419 ( .A(G125), .ZN(n392) );
  INV_X1 U420 ( .A(KEYINPUT6), .ZN(n419) );
  XNOR2_X1 U421 ( .A(n544), .B(KEYINPUT30), .ZN(n415) );
  XNOR2_X1 U422 ( .A(n600), .B(n412), .ZN(n411) );
  INV_X1 U423 ( .A(KEYINPUT101), .ZN(n412) );
  XNOR2_X1 U424 ( .A(n527), .B(n526), .ZN(n670) );
  XNOR2_X1 U425 ( .A(n525), .B(KEYINPUT25), .ZN(n526) );
  XNOR2_X1 U426 ( .A(n384), .B(n485), .ZN(n628) );
  XNOR2_X1 U427 ( .A(n479), .B(n536), .ZN(n384) );
  XNOR2_X1 U428 ( .A(G101), .B(G116), .ZN(n483) );
  XOR2_X1 U429 ( .A(G140), .B(KEYINPUT11), .Z(n495) );
  XNOR2_X1 U430 ( .A(G122), .B(KEYINPUT12), .ZN(n494) );
  XNOR2_X1 U431 ( .A(G143), .B(G131), .ZN(n492) );
  XOR2_X1 U432 ( .A(G104), .B(G113), .Z(n493) );
  NAND2_X1 U433 ( .A1(n581), .A2(n459), .ZN(n668) );
  NOR2_X1 U434 ( .A1(n420), .A2(n554), .ZN(n430) );
  XNOR2_X1 U435 ( .A(n553), .B(n364), .ZN(n420) );
  XNOR2_X1 U436 ( .A(n598), .B(n597), .ZN(n615) );
  INV_X1 U437 ( .A(KEYINPUT22), .ZN(n597) );
  INV_X1 U438 ( .A(KEYINPUT1), .ZN(n448) );
  NOR2_X1 U439 ( .A1(G952), .A2(n745), .ZN(n729) );
  XNOR2_X1 U440 ( .A(KEYINPUT99), .B(n543), .ZN(n657) );
  NOR2_X1 U441 ( .A1(n660), .A2(n650), .ZN(n564) );
  INV_X1 U442 ( .A(n691), .ZN(n396) );
  XOR2_X1 U443 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n511) );
  XOR2_X1 U444 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n481) );
  INV_X1 U445 ( .A(KEYINPUT75), .ZN(n426) );
  XNOR2_X1 U446 ( .A(n532), .B(n455), .ZN(n454) );
  INV_X1 U447 ( .A(KEYINPUT17), .ZN(n455) );
  XNOR2_X1 U448 ( .A(KEYINPUT18), .B(KEYINPUT4), .ZN(n388) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n505) );
  XNOR2_X1 U450 ( .A(n394), .B(KEYINPUT69), .ZN(n552) );
  NAND2_X1 U451 ( .A1(n395), .A2(n671), .ZN(n394) );
  NOR2_X1 U452 ( .A1(n670), .A2(n545), .ZN(n395) );
  NOR2_X2 U453 ( .A1(n616), .A2(n593), .ZN(n673) );
  AND2_X1 U454 ( .A1(n408), .A2(n407), .ZN(n406) );
  NAND2_X1 U455 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n478), .B(G119), .ZN(n536) );
  XNOR2_X1 U457 ( .A(G113), .B(KEYINPUT3), .ZN(n478) );
  XNOR2_X1 U458 ( .A(G128), .B(G119), .ZN(n517) );
  INV_X1 U459 ( .A(G134), .ZN(n473) );
  XOR2_X1 U460 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n488) );
  XNOR2_X1 U461 ( .A(n416), .B(G107), .ZN(n535) );
  XNOR2_X1 U462 ( .A(G122), .B(G116), .ZN(n416) );
  XNOR2_X1 U463 ( .A(n380), .B(n385), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n387), .B(n386), .ZN(n385) );
  XNOR2_X1 U465 ( .A(n531), .B(n391), .ZN(n386) );
  XNOR2_X1 U466 ( .A(n454), .B(n388), .ZN(n387) );
  XNOR2_X1 U467 ( .A(n556), .B(n421), .ZN(n557) );
  INV_X1 U468 ( .A(KEYINPUT105), .ZN(n421) );
  INV_X1 U469 ( .A(KEYINPUT76), .ZN(n428) );
  NOR2_X1 U470 ( .A1(n415), .A2(n545), .ZN(n546) );
  XNOR2_X1 U471 ( .A(n628), .B(KEYINPUT62), .ZN(n629) );
  XNOR2_X1 U472 ( .A(n390), .B(n389), .ZN(n380) );
  XNOR2_X1 U473 ( .A(n536), .B(n533), .ZN(n389) );
  XNOR2_X1 U474 ( .A(n534), .B(n535), .ZN(n390) );
  XOR2_X1 U475 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n533) );
  XNOR2_X1 U476 ( .A(n500), .B(n414), .ZN(n715) );
  XNOR2_X1 U477 ( .A(n515), .B(n499), .ZN(n414) );
  NOR2_X1 U478 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X1 U479 ( .A(KEYINPUT98), .B(n504), .ZN(n655) );
  NOR2_X1 U480 ( .A1(n571), .A2(n542), .ZN(n504) );
  XNOR2_X1 U481 ( .A(n463), .B(n462), .ZN(n754) );
  INV_X1 U482 ( .A(KEYINPUT100), .ZN(n462) );
  NOR2_X1 U483 ( .A1(n674), .A2(n616), .ZN(n464) );
  XNOR2_X1 U484 ( .A(n725), .B(n429), .ZN(n728) );
  XNOR2_X1 U485 ( .A(n452), .B(n451), .ZN(G75) );
  XNOR2_X1 U486 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n451) );
  NAND2_X1 U487 ( .A1(n708), .A2(n453), .ZN(n452) );
  AND2_X1 U488 ( .A1(n707), .A2(n745), .ZN(n453) );
  XNOR2_X1 U489 ( .A(n393), .B(G128), .ZN(n649) );
  INV_X1 U490 ( .A(KEYINPUT29), .ZN(n393) );
  AND2_X1 U491 ( .A1(n566), .A2(n365), .ZN(n360) );
  INV_X1 U492 ( .A(n670), .ZN(n616) );
  XOR2_X1 U493 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n361) );
  NAND2_X1 U494 ( .A1(n674), .A2(n673), .ZN(n602) );
  XOR2_X1 U495 ( .A(KEYINPUT70), .B(G469), .Z(n362) );
  AND2_X1 U496 ( .A1(n664), .A2(n663), .ZN(n363) );
  XNOR2_X1 U497 ( .A(KEYINPUT28), .B(KEYINPUT102), .ZN(n364) );
  XNOR2_X1 U498 ( .A(KEYINPUT47), .B(KEYINPUT67), .ZN(n365) );
  XOR2_X1 U499 ( .A(n591), .B(KEYINPUT35), .Z(n366) );
  XOR2_X1 U500 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n367) );
  XOR2_X1 U501 ( .A(KEYINPUT0), .B(KEYINPUT88), .Z(n368) );
  INV_X1 U502 ( .A(G902), .ZN(n404) );
  INV_X1 U503 ( .A(KEYINPUT34), .ZN(n447) );
  XOR2_X1 U504 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n369) );
  XOR2_X1 U505 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n370) );
  XOR2_X1 U506 ( .A(KEYINPUT68), .B(KEYINPUT48), .Z(n371) );
  BUF_X1 U507 ( .A(n724), .Z(n720) );
  BUF_X1 U508 ( .A(n550), .Z(n562) );
  NOR2_X1 U509 ( .A1(n557), .A2(n372), .ZN(n559) );
  INV_X1 U510 ( .A(n476), .ZN(n377) );
  NAND2_X1 U511 ( .A1(n474), .A2(n475), .ZN(n373) );
  AND2_X1 U512 ( .A1(n474), .A2(n475), .ZN(n423) );
  NAND2_X1 U513 ( .A1(n376), .A2(n374), .ZN(n738) );
  NAND2_X1 U514 ( .A1(n474), .A2(n375), .ZN(n374) );
  NOR2_X1 U515 ( .A1(n436), .A2(n435), .ZN(n434) );
  NAND2_X1 U516 ( .A1(n378), .A2(n437), .ZN(n590) );
  NAND2_X1 U517 ( .A1(n434), .A2(n440), .ZN(n378) );
  NAND2_X1 U518 ( .A1(n397), .A2(n626), .ZN(n540) );
  AND2_X2 U519 ( .A1(n379), .A2(n363), .ZN(n742) );
  XNOR2_X1 U520 ( .A(n579), .B(n371), .ZN(n379) );
  NOR2_X1 U521 ( .A1(n719), .A2(G902), .ZN(n491) );
  XNOR2_X1 U522 ( .A(n422), .B(n489), .ZN(n719) );
  NAND2_X1 U523 ( .A1(n380), .A2(n735), .ZN(n736) );
  XNOR2_X1 U524 ( .A(n382), .B(KEYINPUT57), .ZN(n709) );
  INV_X1 U525 ( .A(n383), .ZN(n618) );
  NAND2_X1 U526 ( .A1(n383), .A2(n685), .ZN(n544) );
  NAND2_X1 U527 ( .A1(n552), .A2(n383), .ZN(n553) );
  XNOR2_X2 U528 ( .A(n383), .B(n419), .ZN(n587) );
  NOR2_X1 U529 ( .A1(n679), .A2(n383), .ZN(n680) );
  NAND2_X1 U530 ( .A1(n628), .A2(G472), .ZN(n408) );
  XNOR2_X1 U531 ( .A(n391), .B(KEYINPUT10), .ZN(n515) );
  NAND2_X1 U532 ( .A1(n651), .A2(n396), .ZN(n555) );
  XNOR2_X1 U533 ( .A(n359), .B(n468), .ZN(n635) );
  NOR2_X1 U534 ( .A1(n574), .A2(n398), .ZN(n651) );
  OR2_X1 U535 ( .A1(n628), .A2(n403), .ZN(n402) );
  NAND2_X1 U536 ( .A1(n445), .A2(n444), .ZN(n439) );
  XNOR2_X2 U537 ( .A(n410), .B(n370), .ZN(n750) );
  NAND2_X1 U538 ( .A1(n570), .A2(n655), .ZN(n410) );
  NAND2_X1 U539 ( .A1(n546), .A2(n411), .ZN(n547) );
  NAND2_X1 U540 ( .A1(n413), .A2(n458), .ZN(n460) );
  NAND2_X1 U541 ( .A1(n456), .A2(n457), .ZN(n413) );
  XNOR2_X1 U542 ( .A(n503), .B(n502), .ZN(n572) );
  AND2_X2 U543 ( .A1(n460), .A2(n668), .ZN(n724) );
  NAND2_X1 U544 ( .A1(n610), .A2(n464), .ZN(n463) );
  XNOR2_X1 U545 ( .A(n516), .B(n361), .ZN(n427) );
  NAND2_X1 U546 ( .A1(n561), .A2(n686), .ZN(n417) );
  AND2_X2 U547 ( .A1(n418), .A2(n673), .ZN(n600) );
  INV_X1 U548 ( .A(n554), .ZN(n418) );
  INV_X1 U549 ( .A(n479), .ZN(n450) );
  NAND2_X1 U550 ( .A1(n682), .A2(n461), .ZN(n603) );
  NAND2_X1 U551 ( .A1(n528), .A2(n587), .ZN(n556) );
  XNOR2_X1 U552 ( .A(n535), .B(n423), .ZN(n422) );
  XNOR2_X1 U553 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U554 ( .A1(n590), .A2(n589), .ZN(n424) );
  NAND2_X1 U555 ( .A1(n425), .A2(n624), .ZN(n625) );
  XNOR2_X1 U556 ( .A(n466), .B(n465), .ZN(n425) );
  XNOR2_X1 U557 ( .A(n742), .B(n426), .ZN(n457) );
  XNOR2_X1 U558 ( .A(n519), .B(n427), .ZN(n522) );
  XNOR2_X1 U559 ( .A(n727), .B(n726), .ZN(n429) );
  XNOR2_X1 U560 ( .A(n430), .B(KEYINPUT103), .ZN(n574) );
  XNOR2_X1 U561 ( .A(n431), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U562 ( .A1(n718), .A2(n729), .ZN(n431) );
  NAND2_X1 U563 ( .A1(n651), .A2(n360), .ZN(n567) );
  NAND2_X1 U564 ( .A1(n432), .A2(n447), .ZN(n433) );
  NAND2_X1 U565 ( .A1(n461), .A2(n439), .ZN(n432) );
  INV_X1 U566 ( .A(n461), .ZN(n435) );
  NAND2_X1 U567 ( .A1(n439), .A2(KEYINPUT34), .ZN(n436) );
  NAND2_X1 U568 ( .A1(n441), .A2(n447), .ZN(n438) );
  NAND2_X1 U569 ( .A1(n440), .A2(n439), .ZN(n703) );
  INV_X1 U570 ( .A(n441), .ZN(n440) );
  NAND2_X1 U571 ( .A1(n443), .A2(n442), .ZN(n441) );
  NAND2_X1 U572 ( .A1(n599), .A2(n446), .ZN(n442) );
  NAND2_X1 U573 ( .A1(n602), .A2(n446), .ZN(n443) );
  INV_X1 U574 ( .A(n602), .ZN(n444) );
  INV_X1 U575 ( .A(KEYINPUT33), .ZN(n446) );
  XNOR2_X2 U576 ( .A(n554), .B(n448), .ZN(n674) );
  XNOR2_X2 U577 ( .A(n449), .B(n362), .ZN(n554) );
  NOR2_X2 U578 ( .A1(n750), .A2(n753), .ZN(n576) );
  INV_X1 U579 ( .A(n665), .ZN(n459) );
  INV_X1 U580 ( .A(n594), .ZN(n461) );
  XNOR2_X1 U581 ( .A(n586), .B(n368), .ZN(n594) );
  NAND2_X1 U582 ( .A1(n467), .A2(n620), .ZN(n466) );
  XNOR2_X1 U583 ( .A(n609), .B(KEYINPUT85), .ZN(n467) );
  XNOR2_X1 U584 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X2 U585 ( .A1(n637), .A2(n729), .ZN(n639) );
  XNOR2_X1 U586 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n468) );
  XNOR2_X1 U587 ( .A(n538), .B(KEYINPUT77), .ZN(n539) );
  XNOR2_X1 U588 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n558) );
  INV_X1 U589 ( .A(KEYINPUT59), .ZN(n714) );
  INV_X1 U590 ( .A(n588), .ZN(n589) );
  XNOR2_X1 U591 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U592 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X2 U593 ( .A1(n631), .A2(n729), .ZN(n634) );
  XNOR2_X1 U594 ( .A(G137), .B(G140), .ZN(n514) );
  XNOR2_X1 U595 ( .A(G107), .B(n514), .ZN(n470) );
  NAND2_X1 U596 ( .A1(G227), .A2(n745), .ZN(n469) );
  XNOR2_X1 U597 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U598 ( .A(n534), .B(n471), .ZN(n477) );
  XNOR2_X2 U599 ( .A(G143), .B(G128), .ZN(n472) );
  NAND2_X1 U600 ( .A1(n472), .A2(G134), .ZN(n475) );
  NAND2_X1 U601 ( .A1(n473), .A2(n531), .ZN(n474) );
  NOR2_X1 U602 ( .A1(G953), .A2(G237), .ZN(n498) );
  NAND2_X1 U603 ( .A1(n498), .A2(G210), .ZN(n480) );
  XNOR2_X1 U604 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U605 ( .A(n482), .B(G137), .Z(n484) );
  XNOR2_X1 U606 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U607 ( .A1(G234), .A2(n745), .ZN(n486) );
  XOR2_X1 U608 ( .A(KEYINPUT8), .B(n486), .Z(n520) );
  NAND2_X1 U609 ( .A1(G217), .A2(n520), .ZN(n487) );
  XNOR2_X1 U610 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U611 ( .A(KEYINPUT97), .B(G478), .ZN(n490) );
  XNOR2_X1 U612 ( .A(n491), .B(n490), .ZN(n571) );
  XNOR2_X1 U613 ( .A(n493), .B(n492), .ZN(n497) );
  XNOR2_X1 U614 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U615 ( .A(n497), .B(n496), .Z(n500) );
  NAND2_X1 U616 ( .A1(G214), .A2(n498), .ZN(n499) );
  NOR2_X1 U617 ( .A1(G902), .A2(n715), .ZN(n503) );
  XNOR2_X1 U618 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n501) );
  INV_X1 U619 ( .A(n572), .ZN(n542) );
  XNOR2_X1 U620 ( .A(n505), .B(KEYINPUT14), .ZN(n506) );
  NAND2_X1 U621 ( .A1(G952), .A2(n506), .ZN(n702) );
  NOR2_X1 U622 ( .A1(G953), .A2(n702), .ZN(n584) );
  NAND2_X1 U623 ( .A1(G902), .A2(n506), .ZN(n507) );
  XOR2_X1 U624 ( .A(KEYINPUT90), .B(n507), .Z(n508) );
  NAND2_X1 U625 ( .A1(G953), .A2(n508), .ZN(n582) );
  NOR2_X1 U626 ( .A1(G900), .A2(n582), .ZN(n509) );
  NOR2_X1 U627 ( .A1(n584), .A2(n509), .ZN(n545) );
  NAND2_X1 U628 ( .A1(G234), .A2(n626), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n511), .B(n510), .ZN(n524) );
  NAND2_X1 U630 ( .A1(G221), .A2(n524), .ZN(n512) );
  XOR2_X1 U631 ( .A(KEYINPUT94), .B(n512), .Z(n513) );
  XOR2_X1 U632 ( .A(KEYINPUT21), .B(n513), .Z(n593) );
  INV_X1 U633 ( .A(n593), .ZN(n671) );
  XNOR2_X1 U634 ( .A(n515), .B(n514), .ZN(n739) );
  XOR2_X1 U635 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n516) );
  XOR2_X1 U636 ( .A(KEYINPUT80), .B(G110), .Z(n518) );
  XNOR2_X1 U637 ( .A(n517), .B(n518), .ZN(n519) );
  NAND2_X1 U638 ( .A1(G221), .A2(n520), .ZN(n521) );
  XNOR2_X1 U639 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U640 ( .A(n739), .B(n523), .ZN(n727) );
  NOR2_X1 U641 ( .A1(n727), .A2(G902), .ZN(n527) );
  NAND2_X1 U642 ( .A1(G217), .A2(n524), .ZN(n525) );
  AND2_X1 U643 ( .A1(n655), .A2(n552), .ZN(n528) );
  NOR2_X1 U644 ( .A1(n674), .A2(n556), .ZN(n529) );
  NAND2_X1 U645 ( .A1(G214), .A2(n537), .ZN(n685) );
  NAND2_X1 U646 ( .A1(n529), .A2(n685), .ZN(n530) );
  XNOR2_X1 U647 ( .A(n530), .B(KEYINPUT43), .ZN(n541) );
  NAND2_X1 U648 ( .A1(G224), .A2(n745), .ZN(n532) );
  NAND2_X1 U649 ( .A1(G210), .A2(n537), .ZN(n538) );
  INV_X1 U650 ( .A(n562), .ZN(n548) );
  NAND2_X1 U651 ( .A1(n541), .A2(n548), .ZN(n664) );
  NAND2_X1 U652 ( .A1(n571), .A2(n542), .ZN(n543) );
  XNOR2_X1 U653 ( .A(KEYINPUT38), .B(KEYINPUT73), .ZN(n549) );
  XOR2_X1 U654 ( .A(n549), .B(n548), .Z(n686) );
  NAND2_X1 U655 ( .A1(n657), .A2(n570), .ZN(n663) );
  XOR2_X1 U656 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n551) );
  NAND2_X1 U657 ( .A1(n555), .A2(KEYINPUT47), .ZN(n565) );
  INV_X1 U658 ( .A(n674), .ZN(n612) );
  NOR2_X1 U659 ( .A1(n612), .A2(n560), .ZN(n660) );
  NAND2_X1 U660 ( .A1(n571), .A2(n572), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U662 ( .A1(n588), .A2(n563), .ZN(n650) );
  NAND2_X1 U663 ( .A1(n565), .A2(n564), .ZN(n569) );
  XOR2_X1 U664 ( .A(n691), .B(KEYINPUT79), .Z(n605) );
  INV_X1 U665 ( .A(n605), .ZN(n566) );
  XOR2_X1 U666 ( .A(KEYINPUT72), .B(n567), .Z(n568) );
  NOR2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n578) );
  NAND2_X1 U668 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U669 ( .A1(n572), .A2(n571), .ZN(n596) );
  INV_X1 U670 ( .A(n596), .ZN(n688) );
  NOR2_X1 U671 ( .A1(n690), .A2(n688), .ZN(n573) );
  XNOR2_X1 U672 ( .A(n573), .B(KEYINPUT41), .ZN(n704) );
  NOR2_X1 U673 ( .A1(n704), .A2(n574), .ZN(n575) );
  XNOR2_X1 U674 ( .A(n575), .B(KEYINPUT42), .ZN(n753) );
  XNOR2_X1 U675 ( .A(n576), .B(KEYINPUT46), .ZN(n577) );
  NAND2_X1 U676 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U677 ( .A1(n742), .A2(KEYINPUT2), .ZN(n580) );
  XNOR2_X1 U678 ( .A(n580), .B(KEYINPUT81), .ZN(n581) );
  NOR2_X1 U679 ( .A1(n582), .A2(G898), .ZN(n583) );
  NOR2_X1 U680 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U681 ( .A(n587), .ZN(n599) );
  INV_X1 U682 ( .A(KEYINPUT82), .ZN(n591) );
  XNOR2_X1 U683 ( .A(n592), .B(KEYINPUT86), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U685 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U686 ( .A1(n600), .A2(n618), .ZN(n601) );
  NOR2_X1 U687 ( .A1(n435), .A2(n601), .ZN(n644) );
  NOR2_X1 U688 ( .A1(n618), .A2(n602), .ZN(n682) );
  XNOR2_X1 U689 ( .A(KEYINPUT31), .B(n603), .ZN(n658) );
  NOR2_X1 U690 ( .A1(n644), .A2(n658), .ZN(n604) );
  NOR2_X1 U691 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U692 ( .A1(n754), .A2(n606), .ZN(n607) );
  NAND2_X1 U693 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n616), .A2(n610), .ZN(n611) );
  XNOR2_X1 U695 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n613) );
  XNOR2_X1 U696 ( .A(n614), .B(n613), .ZN(n752) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U698 ( .A1(n674), .A2(n617), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n647) );
  NAND2_X1 U700 ( .A1(n752), .A2(n647), .ZN(n621) );
  NAND2_X1 U701 ( .A1(KEYINPUT44), .A2(n621), .ZN(n620) );
  INV_X1 U702 ( .A(n621), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n358), .A2(KEYINPUT44), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  INV_X1 U705 ( .A(n626), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n724), .A2(G472), .ZN(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT89), .B(KEYINPUT106), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(KEYINPUT63), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n634), .B(n633), .ZN(G57) );
  NAND2_X1 U710 ( .A1(n724), .A2(G210), .ZN(n636) );
  XNOR2_X1 U711 ( .A(KEYINPUT56), .B(KEYINPUT120), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(G51) );
  NAND2_X1 U713 ( .A1(n655), .A2(n644), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n640), .B(G104), .ZN(G6) );
  XOR2_X1 U715 ( .A(KEYINPUT27), .B(KEYINPUT109), .Z(n642) );
  XNOR2_X1 U716 ( .A(G107), .B(KEYINPUT108), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n642), .B(n641), .ZN(n643) );
  XOR2_X1 U718 ( .A(KEYINPUT26), .B(n643), .Z(n646) );
  NAND2_X1 U719 ( .A1(n644), .A2(n657), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(G9) );
  XNOR2_X1 U721 ( .A(G110), .B(n647), .ZN(G12) );
  NAND2_X1 U722 ( .A1(n651), .A2(n657), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(G30) );
  XOR2_X1 U724 ( .A(G143), .B(n650), .Z(G45) );
  AND2_X1 U725 ( .A1(n655), .A2(n651), .ZN(n653) );
  XNOR2_X1 U726 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U728 ( .A(G146), .B(n654), .ZN(G48) );
  NAND2_X1 U729 ( .A1(n658), .A2(n655), .ZN(n656) );
  XNOR2_X1 U730 ( .A(G113), .B(n656), .ZN(G15) );
  NAND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(G116), .ZN(G18) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT112), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(KEYINPUT37), .ZN(n662) );
  XNOR2_X1 U735 ( .A(G125), .B(n662), .ZN(G27) );
  XNOR2_X1 U736 ( .A(G134), .B(n663), .ZN(G36) );
  XNOR2_X1 U737 ( .A(G140), .B(n664), .ZN(G42) );
  NAND2_X1 U738 ( .A1(n742), .A2(n459), .ZN(n667) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n666) );
  NAND2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n708) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U743 ( .A(KEYINPUT49), .B(n672), .ZN(n678) );
  XNOR2_X1 U744 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n676) );
  NOR2_X1 U745 ( .A1(n673), .A2(n674), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n676), .B(n675), .ZN(n677) );
  NAND2_X1 U747 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT114), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U750 ( .A(KEYINPUT51), .B(n683), .Z(n684) );
  NOR2_X1 U751 ( .A1(n704), .A2(n684), .ZN(n697) );
  NOR2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U754 ( .A(KEYINPUT115), .B(n689), .Z(n694) );
  NOR2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U756 ( .A(KEYINPUT116), .B(n692), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U758 ( .A1(n695), .A2(n703), .ZN(n696) );
  NOR2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n700) );
  XNOR2_X1 U760 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n698) );
  XNOR2_X1 U761 ( .A(n698), .B(KEYINPUT52), .ZN(n699) );
  XOR2_X1 U762 ( .A(n700), .B(n699), .Z(n701) );
  NOR2_X1 U763 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U764 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U765 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U766 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n710), .B(n709), .ZN(n712) );
  NAND2_X1 U768 ( .A1(n720), .A2(G469), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U770 ( .A1(n729), .A2(n713), .ZN(G54) );
  NAND2_X1 U771 ( .A1(n724), .A2(G475), .ZN(n717) );
  XNOR2_X1 U772 ( .A(n719), .B(KEYINPUT122), .ZN(n722) );
  NAND2_X1 U773 ( .A1(G478), .A2(n720), .ZN(n721) );
  XNOR2_X1 U774 ( .A(n722), .B(n721), .ZN(n723) );
  NOR2_X1 U775 ( .A1(n723), .A2(n729), .ZN(G63) );
  XOR2_X1 U776 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n726) );
  NAND2_X1 U777 ( .A1(n720), .A2(G217), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(G66) );
  XOR2_X1 U779 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n731) );
  NAND2_X1 U780 ( .A1(G224), .A2(G953), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n731), .B(n730), .ZN(n732) );
  NAND2_X1 U782 ( .A1(n732), .A2(G898), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n459), .A2(n745), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n734), .A2(n733), .ZN(n737) );
  OR2_X1 U785 ( .A1(n745), .A2(G898), .ZN(n735) );
  XOR2_X1 U786 ( .A(n737), .B(n736), .Z(G69) );
  XOR2_X1 U787 ( .A(n738), .B(n739), .Z(n743) );
  XOR2_X1 U788 ( .A(G227), .B(n743), .Z(n740) );
  NOR2_X1 U789 ( .A1(n745), .A2(n740), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n741), .A2(G900), .ZN(n748) );
  XNOR2_X1 U791 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U792 ( .A(n744), .B(KEYINPUT126), .ZN(n746) );
  NAND2_X1 U793 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U795 ( .A(n749), .B(KEYINPUT127), .ZN(G72) );
  XOR2_X1 U796 ( .A(n750), .B(G131), .Z(G33) );
  XOR2_X1 U797 ( .A(n358), .B(G122), .Z(G24) );
  XNOR2_X1 U798 ( .A(G119), .B(n752), .ZN(G21) );
  XOR2_X1 U799 ( .A(G137), .B(n753), .Z(G39) );
  XNOR2_X1 U800 ( .A(G101), .B(KEYINPUT107), .ZN(n755) );
  XNOR2_X1 U801 ( .A(n755), .B(n754), .ZN(G3) );
endmodule

