//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n540, new_n541, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(new_n451));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  AND2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(G2104), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR3_X1   g037(.A1(new_n462), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n463));
  OAI21_X1  g038(.A(G101), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI211_X1 g041(.A(G137), .B(new_n460), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n460), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  NOR2_X1   g047(.A1(new_n465), .A2(new_n466), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n460), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n475), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  OAI211_X1 g056(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n460), .A2(G114), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(G138), .B(new_n460), .C1(new_n465), .C2(new_n466), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT4), .ZN(new_n487));
  OR2_X1    g062(.A1(new_n465), .A2(new_n466), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G138), .A4(new_n460), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(new_n487), .B2(new_n490), .ZN(G164));
  INV_X1    g066(.A(KEYINPUT5), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G543), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  INV_X1    g069(.A(G543), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(KEYINPUT5), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n492), .A2(KEYINPUT69), .A3(G543), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n496), .A2(new_n497), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n495), .A2(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n503), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n501), .A2(new_n511), .ZN(G166));
  INV_X1    g087(.A(new_n509), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G89), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n498), .A2(G63), .A3(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n504), .A2(G51), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n514), .A2(new_n515), .A3(new_n517), .A4(new_n518), .ZN(G286));
  INV_X1    g094(.A(G286), .ZN(G168));
  AOI22_X1  g095(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n500), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n504), .A2(G52), .ZN(new_n523));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n509), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(G171));
  INV_X1    g101(.A(KEYINPUT70), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n506), .A2(G56), .A3(new_n507), .ZN(new_n528));
  NAND2_X1  g103(.A1(G68), .A2(G543), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n500), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n506), .A2(G81), .A3(new_n508), .A4(new_n507), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n504), .A2(G43), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n527), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NOR3_X1   g110(.A1(new_n530), .A2(new_n533), .A3(new_n527), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND4_X1  g116(.A1(G319), .A2(G483), .A3(G661), .A4(new_n541), .ZN(G188));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n509), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n498), .A2(KEYINPUT71), .A3(new_n508), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G91), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT72), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n544), .A2(new_n548), .A3(G91), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n492), .A2(KEYINPUT69), .A3(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT69), .B1(new_n492), .B2(G543), .ZN(new_n552));
  OAI211_X1 g127(.A(G65), .B(new_n507), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(KEYINPUT6), .A2(G651), .ZN(new_n556));
  NOR2_X1   g131(.A1(KEYINPUT6), .A2(G651), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n504), .A2(new_n560), .A3(G53), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n555), .A2(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n550), .A2(new_n562), .ZN(G299));
  OR2_X1    g138(.A1(new_n522), .A2(new_n525), .ZN(G301));
  INV_X1    g139(.A(G166), .ZN(G303));
  AND4_X1   g140(.A1(KEYINPUT71), .A2(new_n506), .A3(new_n507), .A4(new_n508), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT71), .B1(new_n498), .B2(new_n508), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G87), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n498), .A2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n504), .A2(G49), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n504), .A2(KEYINPUT73), .A3(G49), .ZN(new_n574));
  AOI22_X1  g149(.A1(G651), .A2(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n569), .A2(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n506), .A2(G61), .A3(new_n507), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n498), .A2(KEYINPUT74), .A3(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(new_n585), .A3(G651), .ZN(new_n586));
  OAI211_X1 g161(.A(G48), .B(G543), .C1(new_n556), .C2(new_n557), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n504), .A2(new_n589), .A3(G48), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n568), .A2(G86), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n584), .A2(new_n586), .A3(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n500), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n513), .A2(G85), .B1(G47), .B2(new_n504), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n504), .A2(G54), .ZN(new_n598));
  OAI211_X1 g173(.A(G66), .B(new_n507), .C1(new_n551), .C2(new_n552), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n599), .A2(KEYINPUT77), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  AOI21_X1  g177(.A(KEYINPUT77), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n544), .A2(G92), .A3(new_n545), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .A4(new_n545), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G284));
  OAI21_X1  g185(.A(new_n597), .B1(new_n609), .B2(G868), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n609), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n607), .A2(new_n608), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n498), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n500), .B1(new_n619), .B2(KEYINPUT77), .ZN(new_n620));
  INV_X1    g195(.A(new_n603), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n620), .A2(new_n621), .B1(G54), .B2(new_n504), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n618), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g201(.A1(new_n461), .A2(new_n463), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n488), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(G2100), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n474), .A2(G135), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT78), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(G2105), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n476), .B2(G123), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(G14), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n653), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT80), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n664), .B1(new_n661), .B2(new_n663), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n663), .ZN(new_n667));
  INV_X1    g242(.A(new_n663), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n664), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n676), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n676), .B2(new_n682), .ZN(new_n684));
  AND2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n488), .A2(G127), .ZN(new_n693));
  AND2_X1   g268(.A1(G115), .A2(G2104), .ZN(new_n694));
  OAI21_X1  g269(.A(G2105), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT25), .ZN(new_n696));
  NAND2_X1  g271(.A1(G103), .A2(G2104), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G2105), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n460), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n474), .A2(G139), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n692), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n692), .B2(G33), .ZN(new_n702));
  INV_X1    g277(.A(G2072), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n627), .A2(G105), .B1(new_n474), .B2(G141), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT26), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G129), .B2(new_n476), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n692), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n692), .B2(G32), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n704), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G2084), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n692), .B1(KEYINPUT24), .B2(G34), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(KEYINPUT24), .B2(G34), .ZN(new_n717));
  INV_X1    g292(.A(G160), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G29), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT88), .Z(new_n720));
  OAI221_X1 g295(.A(new_n714), .B1(new_n703), .B2(new_n702), .C1(new_n715), .C2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT89), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NOR2_X1   g298(.A1(G171), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G5), .B2(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(G1961), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n692), .A2(G35), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT91), .Z(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n692), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT29), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n727), .B1(new_n732), .B2(G2090), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n720), .A2(new_n715), .ZN(new_n734));
  INV_X1    g309(.A(G2090), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n731), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n692), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n692), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2078), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n692), .A2(G26), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT28), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n474), .A2(G140), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n476), .A2(G128), .ZN(new_n743));
  OR2_X1    g318(.A1(G104), .A2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n744), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n741), .B1(new_n746), .B2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT87), .B(G2067), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n739), .B(new_n749), .C1(new_n712), .C2(new_n713), .ZN(new_n750));
  NOR3_X1   g325(.A1(new_n733), .A2(new_n736), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n722), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G4), .A2(G16), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n609), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT85), .B(G1348), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n723), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n537), .B2(new_n723), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT86), .B(G1341), .Z(new_n759));
  XOR2_X1   g334(.A(new_n758), .B(new_n759), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n640), .A2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G11), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT30), .B(G28), .Z(new_n763));
  OAI211_X1 g338(.A(new_n761), .B(new_n762), .C1(G29), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n723), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n723), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n764), .B1(G1966), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G1966), .B2(new_n766), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n725), .A2(new_n726), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n756), .B(new_n760), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n723), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n613), .B2(new_n723), .ZN(new_n775));
  INV_X1    g350(.A(G1956), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n768), .A2(new_n771), .A3(new_n769), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n754), .B2(new_n755), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n752), .A2(new_n772), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  MUX2_X1   g355(.A(G6), .B(G305), .S(G16), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT84), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT32), .B(G1981), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT34), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  INV_X1    g361(.A(G288), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n787), .A2(new_n723), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n723), .B2(G23), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n789), .A2(new_n791), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n723), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G166), .B2(new_n723), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G1971), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n795), .A2(G1971), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n792), .A2(new_n793), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT81), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n474), .A2(G131), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n476), .A2(G119), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G25), .B(new_n805), .S(G29), .Z(new_n806));
  XOR2_X1   g381(.A(KEYINPUT35), .B(G1991), .Z(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT82), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n723), .A2(G24), .ZN(new_n810));
  INV_X1    g385(.A(G290), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n723), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT83), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n809), .B1(new_n813), .B2(G1986), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G1986), .B2(new_n813), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n799), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n784), .A2(new_n786), .A3(new_n798), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT36), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n816), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n780), .B1(new_n820), .B2(new_n822), .ZN(G311));
  INV_X1    g398(.A(new_n780), .ZN(new_n824));
  INV_X1    g399(.A(new_n822), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n821), .B1(new_n816), .B2(new_n818), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(G150));
  NAND2_X1  g402(.A1(new_n498), .A2(G67), .ZN(new_n828));
  NAND2_X1  g403(.A1(G80), .A2(G543), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G651), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT92), .B(G93), .Z(new_n832));
  NAND3_X1  g407(.A1(new_n498), .A2(new_n508), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n504), .A2(G55), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT93), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT93), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n833), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n528), .A2(new_n529), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G651), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n531), .A2(new_n532), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT70), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n831), .A2(new_n839), .B1(new_n843), .B2(new_n534), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n833), .A2(new_n837), .A3(new_n834), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n837), .B1(new_n833), .B2(new_n834), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n831), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n841), .A2(new_n842), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n609), .A2(G559), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n855));
  XNOR2_X1  g430(.A(KEYINPUT94), .B(G860), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n839), .B2(new_n831), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n629), .B(new_n805), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n695), .A2(KEYINPUT95), .A3(new_n700), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n709), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n861), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n490), .A2(new_n487), .ZN(new_n869));
  INV_X1    g444(.A(new_n485), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n746), .ZN(new_n872));
  AOI22_X1  g447(.A1(G130), .A2(new_n476), .B1(new_n474), .B2(G142), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n460), .A2(KEYINPUT96), .A3(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT96), .B1(new_n460), .B2(G118), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n480), .B(G160), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n640), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n865), .A2(new_n867), .A3(new_n878), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT97), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n882), .B1(new_n880), .B2(new_n883), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(G37), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT98), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(KEYINPUT98), .A3(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT40), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(new_n888), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n891), .A2(new_n894), .ZN(G395));
  INV_X1    g470(.A(G868), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n609), .B(new_n616), .C1(new_n844), .C2(new_n849), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n847), .B1(new_n535), .B2(new_n536), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n839), .A2(new_n841), .A3(new_n842), .A4(new_n831), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n623), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n618), .A2(new_n622), .ZN(new_n902));
  NAND2_X1  g477(.A1(G299), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n550), .A2(new_n618), .A3(new_n562), .A4(new_n622), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT99), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  AND4_X1   g481(.A1(new_n550), .A2(new_n618), .A3(new_n562), .A4(new_n622), .ZN(new_n907));
  AOI22_X1  g482(.A1(new_n550), .A2(new_n562), .B1(new_n618), .B2(new_n622), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT99), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n909), .A2(new_n910), .A3(new_n900), .A4(new_n897), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n907), .B2(new_n908), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n901), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT100), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n901), .A2(new_n914), .A3(new_n918), .A4(new_n915), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n912), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT42), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n912), .A2(new_n917), .A3(new_n922), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n811), .A2(new_n569), .A3(new_n575), .ZN(new_n926));
  NAND2_X1  g501(.A1(G288), .A2(G290), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G305), .A2(G166), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(G305), .A2(G166), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n926), .A2(new_n927), .A3(new_n925), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n934), .B(new_n930), .C1(new_n935), .C2(new_n928), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n924), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n921), .A2(new_n937), .A3(new_n923), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n896), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n847), .A2(new_n896), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT102), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n940), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n937), .B1(new_n921), .B2(new_n923), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n948), .A3(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n944), .A2(new_n949), .ZN(G295));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n942), .ZN(G331));
  XNOR2_X1  g526(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n952));
  NAND2_X1  g527(.A1(G168), .A2(G171), .ZN(new_n953));
  NAND2_X1  g528(.A1(G301), .A2(G286), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n844), .B2(new_n849), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n898), .A2(new_n899), .B1(new_n953), .B2(new_n954), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n898), .A2(new_n953), .A3(new_n899), .A4(new_n954), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n957), .A2(new_n960), .A3(new_n909), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND4_X1   g539(.A1(new_n898), .A2(new_n953), .A3(new_n899), .A4(new_n954), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n965), .B1(KEYINPUT105), .B2(new_n956), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n966), .A2(KEYINPUT106), .A3(new_n909), .A4(new_n960), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n965), .B1(new_n958), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n956), .A2(KEYINPUT104), .A3(new_n961), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n970), .A3(new_n914), .A4(new_n915), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n964), .A2(new_n967), .A3(new_n937), .A4(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G37), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n937), .A2(KEYINPUT108), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n933), .A2(new_n936), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n966), .A2(new_n960), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n914), .A2(new_n915), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n969), .A2(new_n970), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n979), .A2(new_n980), .B1(new_n981), .B2(new_n909), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT109), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n933), .A2(new_n936), .A3(new_n976), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n976), .B1(new_n933), .B2(new_n936), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n980), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n909), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI211_X1 g566(.A(KEYINPUT43), .B(new_n974), .C1(new_n983), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n964), .A2(new_n971), .A3(new_n967), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT107), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n964), .A2(new_n967), .A3(new_n996), .A4(new_n971), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n997), .A3(new_n986), .ZN(new_n998));
  INV_X1    g573(.A(new_n974), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n952), .B1(new_n992), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n998), .A2(new_n993), .A3(new_n999), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n974), .B1(new_n983), .B2(new_n991), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1002), .B(KEYINPUT44), .C1(new_n1003), .C2(new_n993), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1001), .A2(new_n1004), .ZN(G397));
  INV_X1    g580(.A(G1384), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n871), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(KEYINPUT110), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(KEYINPUT110), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n471), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(G40), .A3(new_n464), .A4(new_n467), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT112), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G160), .A2(new_n1015), .A3(G40), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1996), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n709), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G2067), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n746), .B(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n807), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n805), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n805), .A2(new_n1025), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g604(.A(G290), .B(G1986), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1019), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1007), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1033));
  INV_X1    g608(.A(G8), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n787), .A2(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1037), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(G166), .A2(new_n1034), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(KEYINPUT55), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G164), .A2(G1384), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT45), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1017), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1971), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1045), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1017), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G2090), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1043), .B(G8), .C1(new_n1050), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n590), .A2(new_n588), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n498), .A2(G86), .A3(new_n508), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1058), .A2(KEYINPUT113), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT113), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n584), .A2(new_n1062), .A3(new_n586), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G1981), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n584), .A2(new_n1065), .A3(new_n586), .A4(new_n591), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1057), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT49), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1035), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1057), .B(KEYINPUT49), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1041), .B(new_n1056), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1015), .B1(G160), .B2(G40), .ZN(new_n1072));
  INV_X1    g647(.A(G40), .ZN(new_n1073));
  NOR4_X1   g648(.A1(new_n468), .A2(new_n471), .A3(KEYINPUT112), .A4(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1053), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT115), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT115), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1053), .B(new_n1077), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1076), .A2(new_n735), .A3(new_n1078), .A4(new_n1052), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1049), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1034), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1079), .A2(KEYINPUT116), .A3(new_n1049), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1043), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1071), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G168), .A2(new_n1034), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT51), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1054), .ZN(new_n1091));
  INV_X1    g666(.A(G1966), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT45), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1007), .A2(new_n1093), .ZN(new_n1094));
  OR3_X1    g669(.A1(G164), .A2(G1384), .A3(new_n1009), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1017), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1091), .A2(new_n715), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1090), .B(new_n1087), .C1(new_n1097), .C2(new_n1034), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1092), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(G2084), .B2(new_n1054), .ZN(new_n1100));
  OAI211_X1 g675(.A(G8), .B(new_n1089), .C1(new_n1100), .C2(G286), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1086), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(G301), .B(KEYINPUT54), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1011), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n469), .A2(new_n470), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n460), .B1(new_n1107), .B2(KEYINPUT123), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(KEYINPUT123), .B2(new_n1107), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(G2078), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n468), .A2(new_n1073), .A3(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1046), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1104), .B1(new_n1105), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1110), .B1(new_n1047), .B2(G2078), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1054), .A2(new_n726), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1116), .B(new_n1117), .C1(new_n1096), .C2(new_n1112), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n1104), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1085), .A2(new_n1103), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1122));
  AOI21_X1  g697(.A(new_n560), .B1(new_n504), .B2(G53), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n558), .A2(KEYINPUT9), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT117), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n555), .A2(G651), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n561), .A2(new_n559), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n547), .B2(new_n549), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT118), .B1(new_n1130), .B2(KEYINPUT57), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n548), .B1(new_n568), .B2(G91), .ZN(new_n1133));
  INV_X1    g708(.A(new_n549), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n550), .A2(KEYINPUT57), .A3(new_n562), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1131), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1078), .A2(new_n1052), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1077), .B1(new_n1017), .B2(new_n1053), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n776), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1047), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT119), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1140), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1140), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1122), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1140), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1140), .A2(new_n1143), .A3(new_n1147), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(KEYINPUT61), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1047), .A2(G1996), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT58), .B(G1341), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1033), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n537), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT59), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1150), .A2(new_n1155), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT121), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1150), .A2(new_n1160), .A3(new_n1155), .A4(KEYINPUT121), .ZN(new_n1164));
  INV_X1    g739(.A(G1348), .ZN(new_n1165));
  AOI22_X1  g740(.A1(new_n1054), .A2(new_n1165), .B1(new_n1033), .B2(new_n1022), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT60), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(new_n609), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(KEYINPUT60), .B2(new_n1166), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n1164), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1166), .A2(new_n902), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1154), .B1(new_n1149), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1121), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1119), .A2(G171), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1103), .B2(KEYINPUT62), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1098), .A2(new_n1101), .A3(new_n1176), .A4(new_n1102), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1085), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1041), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1179), .A2(new_n1180), .A3(new_n1056), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n787), .A2(new_n1039), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1066), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1181), .B1(new_n1035), .B2(new_n1183), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1097), .A2(new_n1034), .A3(G286), .ZN(new_n1185));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n1085), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1055), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1034), .B1(new_n1187), .B2(new_n1049), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1185), .B(KEYINPUT63), .C1(new_n1188), .C2(new_n1043), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n1071), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1178), .B(new_n1184), .C1(new_n1186), .C2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1031), .B1(new_n1173), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1026), .B1(new_n1018), .B2(new_n1024), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n746), .A2(G2067), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1195), .A2(KEYINPUT124), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1019), .B1(new_n1195), .B2(KEYINPUT124), .ZN(new_n1197));
  OR3_X1    g772(.A1(new_n1196), .A2(new_n1197), .A3(KEYINPUT125), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1018), .B1(new_n710), .B2(new_n1023), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT46), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(new_n1018), .B2(G1996), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1019), .A2(KEYINPUT46), .A3(new_n1020), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1201), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(KEYINPUT47), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT47), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1201), .A2(new_n1207), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(KEYINPUT125), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1210));
  NOR3_X1   g785(.A1(new_n1018), .A2(G1986), .A3(G290), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1212));
  XNOR2_X1  g787(.A(new_n1211), .B(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT48), .ZN(new_n1214));
  OR2_X1    g789(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1019), .A2(new_n1029), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  AND4_X1   g793(.A1(new_n1198), .A2(new_n1209), .A3(new_n1210), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1192), .A2(new_n1219), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g795(.A1(new_n992), .A2(new_n1000), .ZN(new_n1222));
  INV_X1    g796(.A(G319), .ZN(new_n1223));
  OR2_X1    g797(.A1(G227), .A2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g798(.A1(G229), .A2(G401), .A3(new_n1224), .ZN(new_n1225));
  OAI21_X1  g799(.A(new_n1225), .B1(new_n892), .B2(new_n888), .ZN(new_n1226));
  NOR2_X1   g800(.A1(new_n1222), .A2(new_n1226), .ZN(G308));
  OAI221_X1 g801(.A(new_n1225), .B1(new_n892), .B2(new_n888), .C1(new_n992), .C2(new_n1000), .ZN(G225));
endmodule


