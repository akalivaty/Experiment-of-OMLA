//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  INV_X1    g0009(.A(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  XNOR2_X1  g0011(.A(KEYINPUT67), .B(G244), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT68), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n205), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n205), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT64), .Z(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT0), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n202), .A2(KEYINPUT66), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n222), .A2(G50), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT65), .Z(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR3_X1   g0027(.A1(new_n217), .A2(new_n221), .A3(new_n227), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XOR2_X1   g0035(.A(new_n232), .B(new_n235), .Z(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n211), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  INV_X1    g0041(.A(G107), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n240), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(G58), .B(G68), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  AOI22_X1  g0048(.A1(new_n247), .A2(G20), .B1(G159), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT7), .ZN(new_n251));
  NOR3_X1   g0051(.A1(new_n250), .A2(new_n251), .A3(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G20), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G33), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT77), .ZN(new_n258));
  AOI21_X1  g0058(.A(KEYINPUT77), .B1(new_n255), .B2(new_n257), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n252), .B1(new_n260), .B2(new_n251), .ZN(new_n261));
  OAI211_X1 g0061(.A(KEYINPUT16), .B(new_n249), .C1(new_n261), .C2(new_n209), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G1), .A2(G13), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT70), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n267), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n251), .B1(new_n250), .B2(G20), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n255), .A2(new_n257), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n253), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n209), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n249), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n271), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n262), .A2(new_n269), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT71), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n253), .B2(G1), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n266), .A2(new_n268), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n283), .A2(new_n253), .A3(G1), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n280), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(new_n282), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT79), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n287), .A2(KEYINPUT79), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n255), .A2(new_n257), .A3(G226), .A4(G1698), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n255), .A2(new_n257), .A3(G223), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G87), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n294), .B(new_n296), .C1(new_n254), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n264), .B1(G33), .B2(G41), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n281), .B1(G41), .B2(G45), .ZN(new_n302));
  INV_X1    g0102(.A(G274), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G41), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n306), .A2(G1), .A3(G13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(G232), .A3(new_n302), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n300), .A2(new_n301), .A3(new_n305), .A4(new_n308), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n300), .A2(new_n305), .A3(new_n308), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(G200), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n278), .A2(new_n293), .A3(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n312), .A2(KEYINPUT17), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(KEYINPUT81), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT81), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n278), .A2(new_n293), .A3(new_n311), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n313), .B1(new_n317), .B2(KEYINPUT17), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n278), .A2(new_n293), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n310), .A2(G179), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n310), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n319), .A2(KEYINPUT18), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT18), .B1(new_n319), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT80), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT18), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT80), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n319), .A2(KEYINPUT18), .A3(new_n322), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n318), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n250), .A2(G226), .A3(new_n295), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n250), .A2(G232), .A3(G1698), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G97), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n299), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n307), .A2(G238), .A3(new_n302), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n338), .A2(KEYINPUT74), .A3(new_n305), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT74), .B1(new_n305), .B2(new_n338), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT13), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT13), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n337), .B(new_n343), .C1(new_n339), .C2(new_n340), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT14), .B1(new_n346), .B2(new_n321), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(G179), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n349), .A3(G169), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n285), .A2(new_n286), .ZN(new_n352));
  OR2_X1    g0152(.A1(new_n352), .A2(new_n209), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n253), .A2(G33), .ZN(new_n354));
  OAI22_X1  g0154(.A1(new_n354), .A2(new_n211), .B1(new_n253), .B2(G68), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT75), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n357), .B1(new_n253), .B2(G68), .C1(new_n354), .C2(new_n211), .ZN(new_n358));
  INV_X1    g0158(.A(G50), .ZN(new_n359));
  INV_X1    g0159(.A(new_n248), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n356), .B(new_n358), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(KEYINPUT11), .A3(new_n269), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n269), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT11), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n282), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n209), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT12), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n353), .A2(new_n362), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n351), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n250), .A2(G232), .A3(new_n295), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n250), .A2(G1698), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n372), .B1(new_n242), .B2(new_n250), .C1(new_n373), .C2(new_n210), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n304), .B1(new_n374), .B2(new_n299), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n307), .A2(new_n302), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(new_n212), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G179), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n366), .A2(new_n211), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n279), .A2(new_n360), .B1(new_n253), .B2(new_n211), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT15), .B(G87), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n354), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n269), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n381), .B(new_n385), .C1(new_n352), .C2(new_n211), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n380), .B(new_n386), .C1(G169), .C2(new_n378), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n371), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n369), .B1(new_n345), .B2(G200), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n346), .A2(G190), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT76), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  AND4_X1   g0195(.A1(new_n332), .A2(new_n389), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n354), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n280), .A2(new_n397), .B1(G150), .B2(new_n248), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n253), .B1(new_n201), .B2(new_n359), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n398), .A2(new_n400), .B1(new_n266), .B2(new_n268), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n352), .A2(G50), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(G50), .B2(new_n366), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n404), .A2(KEYINPUT72), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(KEYINPUT72), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n250), .A2(G222), .A3(new_n295), .ZN(new_n408));
  INV_X1    g0208(.A(G223), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n408), .B1(new_n211), .B2(new_n250), .C1(new_n373), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n304), .B1(new_n410), .B2(new_n299), .ZN(new_n411));
  INV_X1    g0211(.A(G226), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n376), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n321), .ZN(new_n414));
  OR2_X1    g0214(.A1(new_n413), .A2(G179), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n407), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n375), .B2(new_n377), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT73), .ZN(new_n419));
  OR3_X1    g0219(.A1(new_n418), .A2(new_n419), .A3(new_n386), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n378), .A2(G190), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n418), .B2(new_n386), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT9), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n407), .A2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(KEYINPUT9), .B(new_n402), .C1(new_n405), .C2(new_n406), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n413), .A2(new_n301), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n413), .A2(G200), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT10), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n427), .A2(new_n429), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT10), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n428), .A4(new_n426), .ZN(new_n434));
  AOI211_X1 g0234(.A(new_n416), .B(new_n424), .C1(new_n431), .C2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n396), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n273), .A2(G20), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n438), .A2(KEYINPUT90), .A3(KEYINPUT22), .A4(G87), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n397), .A2(G116), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT22), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT90), .A4(new_n253), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n297), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n242), .A2(G20), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT23), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n439), .A2(new_n440), .A3(new_n443), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT24), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n442), .A2(new_n297), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n445), .B1(new_n450), .B2(KEYINPUT22), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT24), .A3(new_n440), .A4(new_n443), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n269), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT25), .B1(new_n366), .B2(new_n242), .ZN(new_n454));
  XOR2_X1   g0254(.A(new_n454), .B(KEYINPUT92), .Z(new_n455));
  NAND3_X1  g0255(.A1(new_n366), .A2(KEYINPUT25), .A3(new_n242), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT91), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  INV_X1    g0260(.A(G45), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n461), .A2(G1), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n299), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G264), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT93), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT93), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n466), .A3(G264), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n250), .A2(G257), .A3(G1698), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n250), .A2(G250), .A3(new_n295), .ZN(new_n469));
  INV_X1    g0269(.A(G294), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n468), .B(new_n469), .C1(new_n254), .C2(new_n470), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n465), .A2(new_n467), .B1(new_n299), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n460), .A2(new_n462), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G274), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G200), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(G190), .A3(new_n474), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n266), .A2(new_n268), .A3(new_n282), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n281), .A2(G33), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(G107), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n459), .A2(new_n476), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n255), .A2(new_n257), .A3(G244), .A4(new_n295), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n250), .A2(KEYINPUT4), .A3(G244), .A4(new_n295), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n250), .A2(G250), .A3(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n299), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n463), .A2(G257), .B1(new_n473), .B2(G274), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT82), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G190), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(G200), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n266), .A2(new_n268), .A3(new_n282), .A4(new_n479), .ZN(new_n499));
  INV_X1    g0299(.A(G97), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT7), .B1(new_n273), .B2(new_n253), .ZN(new_n502));
  OAI21_X1  g0302(.A(G107), .B1(new_n252), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n242), .A2(KEYINPUT6), .A3(G97), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n500), .A2(new_n242), .ZN(new_n505));
  NOR2_X1   g0305(.A1(G97), .A2(G107), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n248), .A2(G77), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n501), .B1(new_n511), .B2(new_n269), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n282), .A2(G97), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n497), .A2(new_n498), .A3(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n255), .A2(new_n257), .A3(G238), .A4(new_n295), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT84), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n250), .A2(new_n520), .A3(G238), .A4(new_n295), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n250), .A2(G244), .A3(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G116), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n519), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n299), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n281), .A2(G45), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT83), .B1(new_n526), .B2(new_n303), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n462), .A2(new_n528), .A3(G274), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n307), .A2(G250), .A3(new_n526), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(G200), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  AOI211_X1 g0334(.A(G190), .B(new_n532), .C1(new_n524), .C2(new_n299), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n253), .B1(new_n335), .B2(new_n537), .ZN(new_n538));
  NOR4_X1   g0338(.A1(KEYINPUT85), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT85), .ZN(new_n540));
  NOR2_X1   g0340(.A1(G87), .A2(G97), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n242), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n538), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n250), .A2(new_n253), .A3(G68), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n537), .B1(new_n354), .B2(new_n500), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT86), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n543), .A2(new_n548), .A3(new_n544), .A4(new_n545), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n269), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n383), .A2(new_n366), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n478), .A2(G87), .A3(new_n479), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n532), .B1(new_n524), .B2(new_n299), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G169), .ZN(new_n556));
  AOI211_X1 g0356(.A(G179), .B(new_n532), .C1(new_n524), .C2(new_n299), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g0358(.A1(new_n499), .A2(new_n383), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n550), .A2(new_n559), .A3(new_n551), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n536), .A2(new_n554), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n493), .A2(new_n321), .A3(new_n495), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n490), .A2(new_n379), .A3(new_n491), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n515), .A3(new_n563), .ZN(new_n564));
  AND4_X1   g0364(.A1(new_n481), .A2(new_n517), .A3(new_n561), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n453), .A2(new_n480), .A3(new_n458), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n475), .A2(new_n321), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n472), .A2(new_n379), .A3(new_n474), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n488), .B(new_n253), .C1(G33), .C2(new_n500), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n244), .A2(G20), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n265), .A2(KEYINPUT88), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT88), .B1(new_n265), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n570), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(KEYINPUT20), .B(new_n570), .C1(new_n572), .C2(new_n573), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n478), .A2(KEYINPUT87), .A3(G116), .A4(new_n479), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT87), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n499), .B2(new_n244), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n366), .A2(new_n244), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n255), .A2(new_n257), .A3(G257), .A4(new_n295), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n255), .A2(new_n257), .A3(G264), .A4(G1698), .ZN(new_n586));
  INV_X1    g0386(.A(G303), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n250), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n299), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n463), .A2(G270), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n474), .A3(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n591), .A2(G169), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n589), .A2(G179), .A3(new_n474), .A4(new_n590), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n593), .A2(new_n594), .B1(new_n596), .B2(new_n584), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT89), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n591), .A2(G169), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n576), .A2(new_n577), .B1(new_n244), .B2(new_n366), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n599), .B1(new_n600), .B2(new_n582), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n601), .B2(KEYINPUT21), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n598), .A2(new_n584), .A3(KEYINPUT21), .A4(new_n592), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n569), .B(new_n597), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n584), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n591), .A2(G200), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n607), .C1(new_n301), .C2(new_n591), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n437), .A2(new_n565), .A3(new_n605), .A4(new_n608), .ZN(G372));
  NAND2_X1  g0409(.A1(new_n565), .A2(new_n604), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n550), .A2(new_n559), .A3(new_n551), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n555), .A2(new_n379), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(G169), .B2(new_n555), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n564), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(new_n561), .A3(KEYINPUT26), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n534), .A2(new_n535), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n611), .A2(new_n613), .B1(new_n618), .B2(new_n553), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n619), .B2(new_n564), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n614), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n437), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n323), .A2(new_n324), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n392), .B1(new_n371), .B2(new_n388), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n625), .B1(new_n626), .B2(new_n318), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n431), .A2(new_n434), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n416), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n623), .A2(new_n629), .ZN(G369));
  INV_X1    g0430(.A(G13), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n281), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n566), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT95), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n481), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n569), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n569), .A2(new_n638), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT94), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT89), .B1(new_n593), .B2(new_n594), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n601), .A2(new_n598), .A3(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n597), .ZN(new_n652));
  INV_X1    g0452(.A(new_n638), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n606), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n652), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n608), .ZN(new_n656));
  INV_X1    g0456(.A(G330), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n656), .A2(new_n648), .A3(new_n657), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n647), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n652), .A2(new_n653), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n644), .B1(new_n643), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n661), .A2(new_n664), .ZN(G399));
  OR3_X1    g0465(.A1(new_n539), .A2(new_n542), .A3(G116), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n218), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n667), .A2(G1), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n224), .B2(new_n670), .ZN(new_n672));
  XOR2_X1   g0472(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n673));
  XNOR2_X1  g0473(.A(new_n672), .B(new_n673), .ZN(new_n674));
  AOI211_X1 g0474(.A(KEYINPUT29), .B(new_n638), .C1(new_n610), .C2(new_n621), .ZN(new_n675));
  INV_X1    g0475(.A(new_n614), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT26), .B1(new_n615), .B2(new_n561), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n619), .A2(new_n564), .A3(new_n617), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(KEYINPUT99), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT99), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n621), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n604), .A2(KEYINPUT100), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT100), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n651), .A2(new_n684), .A3(new_n597), .A4(new_n569), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n683), .A2(new_n565), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n680), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n653), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n675), .B1(new_n688), .B2(KEYINPUT29), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT97), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n595), .B(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n472), .A2(new_n555), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n496), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n555), .B1(new_n472), .B2(new_n474), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n379), .A3(new_n492), .A4(new_n591), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n691), .A2(new_n496), .A3(new_n692), .A4(KEYINPUT30), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n699), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT31), .B1(new_n699), .B2(new_n638), .ZN(new_n702));
  OAI21_X1  g0502(.A(KEYINPUT98), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n702), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT98), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n700), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n565), .A2(new_n605), .A3(new_n608), .A4(new_n653), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n689), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n674), .B1(new_n711), .B2(G1), .ZN(G364));
  AOI21_X1  g0512(.A(new_n281), .B1(new_n632), .B2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n669), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n264), .B1(G20), .B2(new_n321), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT102), .B(G159), .Z(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n253), .A2(G190), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G179), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT32), .ZN(new_n724));
  NAND3_X1  g0524(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(new_n301), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n253), .B1(new_n721), .B2(G190), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n724), .B1(new_n359), .B2(new_n727), .C1(new_n500), .C2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n253), .A2(new_n301), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n417), .A2(G179), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n297), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n379), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n720), .A2(new_n734), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g0538(.A1(G58), .A2(new_n736), .B1(new_n738), .B2(G77), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n720), .A2(new_n731), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n725), .A2(G190), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI221_X1 g0542(.A(new_n739), .B1(new_n242), .B2(new_n740), .C1(new_n209), .C2(new_n742), .ZN(new_n743));
  NOR4_X1   g0543(.A1(new_n729), .A2(new_n273), .A3(new_n733), .A4(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n250), .B1(new_n726), .B2(G326), .ZN(new_n745));
  INV_X1    g0545(.A(G317), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT33), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n741), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n745), .B(new_n749), .C1(new_n750), .C2(new_n737), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n736), .A2(G322), .ZN(new_n752));
  INV_X1    g0552(.A(new_n722), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G329), .ZN(new_n754));
  AND2_X1   g0554(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n755), .B1(new_n756), .B2(new_n740), .C1(new_n587), .C2(new_n732), .ZN(new_n757));
  INV_X1    g0557(.A(new_n728), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n751), .B(new_n757), .C1(G294), .C2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n717), .B1(new_n744), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n240), .A2(G45), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n258), .A2(new_n259), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n668), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n224), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT101), .Z(new_n765));
  AOI22_X1  g0565(.A1(new_n761), .A2(new_n765), .B1(new_n244), .B2(new_n668), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n250), .A2(G355), .A3(new_n218), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n717), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n760), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n716), .B(new_n774), .C1(new_n656), .C2(new_n771), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n659), .A2(new_n660), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n715), .B1(new_n656), .B2(new_n657), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(G396));
  AOI21_X1  g0579(.A(new_n638), .B1(new_n610), .B2(new_n621), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n387), .A2(new_n638), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n386), .A2(new_n638), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n423), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n781), .B1(new_n783), .B2(new_n387), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n780), .B(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n709), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n716), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n717), .A2(new_n769), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n716), .B1(new_n211), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT103), .Z(new_n791));
  INV_X1    g0591(.A(new_n717), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n738), .A2(new_n718), .B1(G137), .B2(new_n726), .ZN(new_n793));
  INV_X1    g0593(.A(G150), .ZN(new_n794));
  XOR2_X1   g0594(.A(KEYINPUT104), .B(G143), .Z(new_n795));
  OAI221_X1 g0595(.A(new_n793), .B1(new_n794), .B2(new_n742), .C1(new_n735), .C2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT105), .B(KEYINPUT34), .Z(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n740), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G68), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n796), .A2(new_n797), .ZN(new_n801));
  INV_X1    g0601(.A(G132), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n732), .A2(new_n359), .B1(new_n722), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n762), .ZN(new_n804));
  AOI211_X1 g0604(.A(new_n803), .B(new_n804), .C1(G58), .C2(new_n758), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n798), .A2(new_n800), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n742), .A2(new_n756), .B1(new_n727), .B2(new_n587), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n250), .B(new_n807), .C1(G87), .C2(new_n799), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n737), .A2(new_n244), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n735), .A2(new_n470), .B1(new_n722), .B2(new_n750), .ZN(new_n810));
  INV_X1    g0610(.A(new_n732), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n809), .B(new_n810), .C1(G107), .C2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n808), .B(new_n812), .C1(new_n500), .C2(new_n728), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n791), .B1(new_n792), .B2(new_n814), .C1(new_n784), .C2(new_n770), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n788), .A2(new_n815), .ZN(G384));
  INV_X1    g0616(.A(new_n636), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n319), .B(new_n817), .C1(new_n318), .C2(new_n624), .ZN(new_n818));
  XOR2_X1   g0618(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n314), .B2(new_n316), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n319), .B1(new_n322), .B2(new_n817), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n312), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n819), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n261), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n276), .B1(new_n829), .B2(G68), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n269), .B(new_n262), .C1(new_n830), .C2(new_n270), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n289), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n817), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n322), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n317), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n822), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n837), .B(KEYINPUT38), .C1(new_n332), .C2(new_n833), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n828), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n704), .A2(new_n707), .A3(new_n700), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n369), .A2(new_n638), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n393), .A2(new_n395), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n351), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT107), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n841), .B(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n370), .A2(new_n392), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n785), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n839), .A2(KEYINPUT40), .A3(new_n840), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n840), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n325), .A2(new_n331), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n317), .A2(KEYINPUT17), .ZN(new_n852));
  INV_X1    g0652(.A(new_n313), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n833), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n835), .A2(KEYINPUT37), .B1(new_n821), .B2(new_n820), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n827), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n850), .B1(new_n838), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n849), .B1(new_n858), .B2(KEYINPUT40), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT109), .ZN(new_n860));
  INV_X1    g0660(.A(new_n840), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n436), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n860), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(G330), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n370), .A2(new_n638), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n855), .A2(new_n827), .A3(new_n856), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n818), .B2(new_n825), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n866), .A2(KEYINPUT39), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n857), .B2(new_n838), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n865), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n857), .A2(new_n838), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n481), .A2(new_n517), .A3(new_n561), .A4(new_n564), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n605), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n653), .B(new_n784), .C1(new_n874), .C2(new_n679), .ZN(new_n875));
  INV_X1    g0675(.A(new_n781), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n844), .A2(new_n847), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n872), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n625), .A2(new_n817), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n871), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n629), .B1(new_n689), .B2(new_n436), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n882), .B(new_n883), .Z(new_n884));
  XNOR2_X1  g0684(.A(new_n864), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n281), .B2(new_n632), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n244), .B1(new_n508), .B2(KEYINPUT35), .ZN(new_n887));
  INV_X1    g0687(.A(new_n226), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n887), .B(new_n888), .C1(KEYINPUT35), .C2(new_n508), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT36), .ZN(new_n890));
  INV_X1    g0690(.A(G58), .ZN(new_n891));
  OAI21_X1  g0691(.A(G77), .B1(new_n891), .B2(new_n209), .ZN(new_n892));
  OAI22_X1  g0692(.A1(new_n224), .A2(new_n892), .B1(G50), .B2(new_n209), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(G1), .A3(new_n631), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT106), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n886), .A2(new_n890), .A3(new_n895), .ZN(G367));
  OAI221_X1 g0696(.A(new_n804), .B1(new_n242), .B2(new_n728), .C1(new_n470), .C2(new_n742), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(G311), .B2(new_n726), .ZN(new_n898));
  AOI22_X1  g0698(.A1(G303), .A2(new_n736), .B1(new_n738), .B2(G283), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n746), .B2(new_n722), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT46), .B1(new_n732), .B2(new_n244), .ZN(new_n901));
  OR3_X1    g0701(.A1(new_n732), .A2(KEYINPUT46), .A3(new_n244), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n898), .B(new_n903), .C1(new_n500), .C2(new_n740), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n799), .A2(G77), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n753), .A2(G137), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(new_n359), .C2(new_n737), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n273), .B(new_n907), .C1(new_n741), .C2(new_n718), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n758), .A2(G68), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n909), .B1(new_n794), .B2(new_n735), .C1(new_n727), .C2(new_n795), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT111), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(KEYINPUT111), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n732), .A2(new_n891), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT47), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n716), .B1(new_n916), .B2(new_n717), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n554), .A2(new_n653), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n614), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n619), .B2(new_n918), .ZN(new_n920));
  INV_X1    g0720(.A(new_n771), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n763), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n772), .B1(new_n218), .B2(new_n383), .C1(new_n235), .C2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n660), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n646), .B1(new_n926), .B2(new_n658), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n564), .A2(new_n638), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n515), .A2(new_n638), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n517), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n928), .B1(new_n930), .B2(new_n564), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n647), .A2(new_n663), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n928), .B1(new_n932), .B2(KEYINPUT42), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n644), .A2(new_n517), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n933), .B(new_n934), .C1(KEYINPUT42), .C2(new_n932), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n920), .B(KEYINPUT43), .Z(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n936), .B2(new_n937), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n927), .B(new_n931), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n927), .A2(new_n931), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n944), .B(new_n945), .C1(new_n939), .C2(new_n938), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n926), .A2(new_n658), .A3(new_n646), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n661), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n663), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n661), .A2(new_n948), .A3(new_n662), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n710), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n664), .A2(new_n931), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT45), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n664), .A2(new_n956), .A3(new_n931), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n956), .B1(new_n664), .B2(new_n931), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n955), .A2(new_n661), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n955), .A2(new_n959), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n927), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n952), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n711), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n669), .B(KEYINPUT41), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n714), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n925), .B1(new_n947), .B2(new_n966), .ZN(G387));
  NAND2_X1  g0767(.A1(new_n950), .A2(new_n951), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n714), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT112), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n968), .A2(KEYINPUT112), .A3(new_n714), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n968), .A2(new_n711), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n950), .A2(new_n710), .A3(new_n951), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n669), .B(KEYINPUT115), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(G68), .A2(G77), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT50), .B1(new_n279), .B2(G50), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n279), .A2(KEYINPUT50), .A3(G50), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n980), .A2(G45), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n667), .A2(new_n978), .A3(new_n979), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n923), .B1(new_n232), .B2(G45), .ZN(new_n983));
  NOR3_X1   g0783(.A1(new_n667), .A2(new_n668), .A3(new_n273), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n668), .A2(new_n242), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n773), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n753), .A2(G326), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n735), .A2(new_n746), .B1(new_n737), .B2(new_n587), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n989), .A2(KEYINPUT114), .B1(G311), .B2(new_n741), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(KEYINPUT114), .B2(new_n989), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G322), .B2(new_n726), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT48), .Z(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n756), .B2(new_n728), .C1(new_n470), .C2(new_n732), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT49), .ZN(new_n995));
  AOI211_X1 g0795(.A(new_n762), .B(new_n988), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n995), .B2(new_n994), .C1(new_n244), .C2(new_n740), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n732), .A2(new_n211), .B1(new_n740), .B2(new_n500), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n998), .B(new_n804), .C1(G150), .C2(new_n753), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT113), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n728), .A2(new_n383), .ZN(new_n1001));
  INV_X1    g0801(.A(G159), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n1002), .A2(new_n727), .B1(new_n742), .B2(new_n279), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(G50), .C2(new_n736), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1000), .B(new_n1004), .C1(new_n209), .C2(new_n737), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n997), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n987), .B1(new_n1006), .B2(new_n717), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1007), .B(new_n715), .C1(new_n647), .C2(new_n921), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n973), .A2(new_n977), .A3(new_n1008), .ZN(G393));
  NAND3_X1  g0809(.A1(new_n962), .A2(KEYINPUT116), .A3(new_n960), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n960), .A2(KEYINPUT116), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT117), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1010), .A2(new_n1011), .A3(KEYINPUT117), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n714), .A3(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n245), .A2(new_n763), .B1(G97), .B2(new_n668), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n772), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n727), .A2(new_n794), .B1(new_n735), .B2(new_n1002), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT51), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n795), .A2(new_n722), .B1(new_n740), .B2(new_n297), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n742), .A2(new_n359), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n732), .A2(new_n209), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n737), .A2(new_n279), .ZN(new_n1024));
  NOR4_X1   g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n758), .A2(G77), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1020), .A2(new_n1025), .A3(new_n762), .A4(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n727), .A2(new_n746), .B1(new_n735), .B2(new_n750), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT52), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G283), .A2(new_n811), .B1(new_n753), .B2(G322), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n250), .B1(new_n758), .B2(G116), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n799), .A2(G107), .B1(G303), .B2(new_n741), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n737), .A2(new_n470), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1027), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n716), .B1(new_n1035), .B2(new_n717), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1018), .B(new_n1036), .C1(new_n931), .C2(new_n921), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n963), .B(new_n976), .C1(new_n1012), .C2(new_n952), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1016), .A2(new_n1037), .A3(new_n1038), .ZN(G390));
  NAND4_X1  g0839(.A1(new_n396), .A2(G330), .A3(new_n435), .A4(new_n840), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n629), .C1(new_n689), .C2(new_n436), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n785), .A2(new_n657), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n878), .B1(new_n708), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n878), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1042), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n861), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n877), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n616), .A2(new_n620), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n681), .B1(new_n1048), .B2(new_n676), .ZN(new_n1049));
  AOI211_X1 g0849(.A(KEYINPUT99), .B(new_n614), .C1(new_n616), .C2(new_n620), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n638), .B1(new_n1051), .B2(new_n686), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n783), .A2(new_n387), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n781), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n708), .A2(new_n878), .A3(new_n1042), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1044), .B1(new_n861), .B2(new_n1045), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1041), .B1(new_n1047), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1046), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n865), .B1(new_n877), .B2(new_n878), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n868), .A2(new_n1060), .A3(new_n870), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n687), .A2(new_n653), .A3(new_n1053), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1044), .B1(new_n1062), .B2(new_n876), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n865), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n866), .B2(new_n867), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1059), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n865), .B1(new_n828), .B2(new_n838), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1054), .B2(new_n1044), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1055), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n872), .A2(KEYINPUT39), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n781), .B1(new_n780), .B2(new_n784), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1064), .B1(new_n1072), .B2(new_n1044), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n828), .A2(new_n838), .A3(new_n869), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1069), .A2(new_n1070), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1067), .A2(new_n1076), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n1061), .A2(new_n1066), .A3(new_n1055), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1046), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1079));
  OAI211_X1 g0879(.A(KEYINPUT118), .B(new_n1058), .C1(new_n1078), .C2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT118), .B1(new_n1077), .B2(new_n1058), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n976), .B1(new_n1058), .B2(new_n1077), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1071), .A2(new_n769), .A3(new_n1074), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n800), .B1(new_n244), .B2(new_n735), .C1(new_n470), .C2(new_n722), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n733), .B(new_n1085), .C1(G97), .C2(new_n738), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n741), .A2(G107), .B1(new_n726), .B2(G283), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1086), .A2(new_n273), .A3(new_n1026), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(G125), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n250), .B1(new_n722), .B2(new_n1089), .C1(new_n359), .C2(new_n740), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n732), .A2(new_n794), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT53), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n727), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1090), .B(new_n1094), .C1(G132), .C2(new_n736), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n758), .A2(G159), .B1(G137), .B2(new_n741), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT54), .B(G143), .Z(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n737), .B2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT119), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(KEYINPUT119), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1095), .A2(new_n1096), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n792), .B1(new_n1088), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n279), .B2(new_n789), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1084), .A2(new_n715), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1106), .A2(KEYINPUT120), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n1077), .B2(new_n714), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1083), .A2(new_n1107), .A3(new_n1109), .ZN(G378));
  INV_X1    g0910(.A(KEYINPUT57), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1058), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1041), .B1(new_n1114), .B2(new_n1080), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n849), .B(G330), .C1(new_n858), .C2(KEYINPUT40), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n882), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n416), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n407), .A2(new_n817), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n628), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n628), .B2(new_n1119), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT55), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1123), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT55), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1125), .A2(new_n1126), .A3(new_n1121), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1124), .A2(new_n1127), .A3(KEYINPUT56), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT56), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1116), .A2(new_n881), .A3(new_n871), .A4(new_n879), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1118), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1130), .B1(new_n1118), .B2(new_n1131), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1111), .B1(new_n1115), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1041), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1133), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1118), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1140), .A3(KEYINPUT57), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1135), .A2(new_n1141), .A3(new_n976), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1130), .A2(new_n769), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n789), .A2(new_n359), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G41), .B1(new_n762), .B2(G33), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1145), .A2(G50), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n738), .A2(G137), .B1(G132), .B2(new_n741), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT121), .Z(new_n1148));
  NOR2_X1   g0948(.A1(new_n1099), .A2(new_n732), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT122), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n758), .A2(G150), .B1(G125), .B2(new_n726), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT123), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n736), .A2(G128), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1148), .A2(new_n1150), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G33), .B(new_n1155), .C1(new_n799), .C2(new_n718), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G41), .B1(new_n753), .B2(G124), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1146), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n740), .A2(new_n891), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n737), .A2(new_n383), .B1(new_n722), .B2(new_n756), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(G107), .C2(new_n736), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n211), .B2(new_n732), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n909), .B1(new_n727), .B2(new_n244), .C1(new_n500), .C2(new_n742), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1162), .A2(new_n1163), .A3(G41), .A4(new_n762), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n1164), .B(KEYINPUT58), .Z(new_n1165));
  AOI21_X1  g0965(.A(new_n792), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1144), .B1(new_n1166), .B2(KEYINPUT124), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(KEYINPUT124), .B2(new_n1166), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1143), .A2(new_n715), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n1140), .B2(new_n714), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1142), .A2(new_n1170), .ZN(G375));
  NAND2_X1  g0971(.A1(new_n1044), .A2(new_n769), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n737), .A2(new_n242), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n500), .A2(new_n732), .B1(new_n735), .B2(new_n756), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G303), .C2(new_n753), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n742), .A2(new_n244), .B1(new_n727), .B2(new_n470), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1176), .A2(new_n250), .A3(new_n1001), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n905), .A3(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n737), .A2(new_n794), .B1(new_n722), .B2(new_n1093), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1159), .B(new_n1179), .C1(G137), .C2(new_n736), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n758), .A2(G50), .B1(new_n1098), .B2(new_n741), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n804), .B1(G159), .B2(new_n811), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n727), .A2(new_n802), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1178), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1185), .A2(new_n717), .B1(new_n209), .B2(new_n789), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1172), .A2(new_n715), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1047), .A2(new_n1057), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n714), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1047), .A2(new_n1041), .A3(new_n1057), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(new_n965), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1191), .B2(new_n1058), .ZN(G381));
  XOR2_X1   g0992(.A(G375), .B(KEYINPUT125), .Z(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(G378), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n925), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n943), .A2(new_n946), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n966), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n973), .A2(new_n778), .A3(new_n977), .A4(new_n1008), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(G390), .A2(new_n1199), .A3(G384), .A4(G381), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1194), .A2(new_n1198), .A3(new_n1200), .ZN(G407));
  INV_X1    g1001(.A(G213), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1194), .B2(new_n637), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(G407), .ZN(G409));
  NOR2_X1   g1004(.A1(new_n1202), .A2(G343), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1142), .A2(G378), .A3(new_n1170), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1083), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1137), .A2(new_n1140), .A3(new_n965), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1170), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1205), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT60), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1190), .B1(new_n1058), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT126), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT126), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n1190), .C1(new_n1058), .C2(new_n1212), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1190), .A2(new_n1212), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1216), .A3(new_n976), .A4(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G384), .B1(new_n1218), .B2(new_n1189), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(G384), .A3(new_n1189), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1205), .A2(G2897), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT63), .B1(new_n1211), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1222), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1211), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT112), .B1(new_n968), .B2(new_n714), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n970), .B(new_n713), .C1(new_n950), .C2(new_n951), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1008), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n1235));
  OAI21_X1  g1035(.A(G396), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(G390), .A2(new_n1199), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(G390), .B1(new_n1199), .B2(new_n1236), .ZN(new_n1239));
  OAI21_X1  g1039(.A(G387), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G390), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1236), .A2(new_n1199), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1198), .A2(new_n1243), .A3(new_n1237), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1240), .A2(new_n1244), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1205), .B(new_n1222), .C1(new_n1206), .C2(new_n1210), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(KEYINPUT63), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1231), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT62), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1211), .A2(new_n1250), .A3(new_n1229), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1248), .B1(new_n1211), .B2(new_n1227), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n1211), .B2(new_n1229), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1245), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1249), .B1(new_n1254), .B2(new_n1255), .ZN(G405));
  NAND2_X1  g1056(.A1(G375), .A2(new_n1207), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1222), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1206), .A2(KEYINPUT127), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1229), .A2(new_n1207), .A3(G375), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1259), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1245), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1263), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(new_n1255), .A3(new_n1261), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(G402));
endmodule


