//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  AND2_X1   g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n464), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(new_n469), .B2(G112), .ZN(new_n473));
  OR3_X1    g048(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n474));
  OAI21_X1  g049(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n467), .A2(new_n469), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  AOI211_X1 g054(.A(new_n476), .B(new_n479), .C1(G136), .C2(new_n468), .ZN(G162));
  OAI211_X1 g055(.A(G138), .B(new_n469), .C1(new_n465), .C2(new_n466), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT68), .B(G114), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n469), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .A4(new_n469), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n483), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G164));
  NAND2_X1  g066(.A1(G75), .A2(G543), .ZN(new_n492));
  INV_X1    g067(.A(G543), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n493), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n496));
  AOI21_X1  g071(.A(KEYINPUT69), .B1(new_n493), .B2(KEYINPUT5), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G62), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n493), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(G88), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI21_X1  g085(.A(G543), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n508), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n508), .B2(new_n513), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n501), .B1(new_n516), .B2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  AOI211_X1 g094(.A(KEYINPUT71), .B(new_n494), .C1(new_n504), .C2(new_n505), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n504), .A2(new_n505), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(new_n495), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n506), .A2(new_n507), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n511), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g105(.A(KEYINPUT72), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n528), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n525), .A2(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n527), .A2(G90), .B1(new_n532), .B2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n524), .B2(G64), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  OAI211_X1 g117(.A(KEYINPUT73), .B(new_n538), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n498), .A2(KEYINPUT71), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n506), .A2(new_n521), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G64), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n542), .B1(new_n547), .B2(new_n539), .ZN(new_n548));
  AOI21_X1  g123(.A(KEYINPUT72), .B1(new_n507), .B2(G543), .ZN(new_n549));
  INV_X1    g124(.A(new_n531), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n551), .A2(new_n552), .B1(new_n553), .B2(new_n526), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n544), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n543), .A2(new_n555), .ZN(G171));
  AND3_X1   g131(.A1(new_n545), .A2(G56), .A3(new_n546), .ZN(new_n557));
  AND2_X1   g132(.A1(G68), .A2(G543), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n527), .A2(G81), .B1(new_n532), .B2(G43), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  OAI211_X1 g143(.A(G53), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(KEYINPUT74), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n507), .A2(new_n572), .A3(G53), .A4(G543), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT75), .B1(new_n569), .B2(KEYINPUT9), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n573), .B2(new_n570), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT76), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n570), .A2(new_n573), .ZN(new_n579));
  INV_X1    g154(.A(new_n576), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n581), .A2(new_n582), .A3(new_n574), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G91), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n585), .A2(new_n542), .B1(new_n586), .B2(new_n526), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G299));
  AND2_X1   g164(.A1(new_n543), .A2(new_n555), .ZN(G301));
  INV_X1    g165(.A(G168), .ZN(G286));
  NAND3_X1  g166(.A1(new_n506), .A2(G87), .A3(new_n507), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n512), .A2(G49), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(G74), .B1(new_n545), .B2(new_n546), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n542), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g173(.A(KEYINPUT77), .B(new_n594), .C1(new_n595), .C2(new_n542), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(G288));
  AOI22_X1  g176(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n542), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n512), .A2(G48), .ZN(new_n604));
  INV_X1    g179(.A(G86), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n526), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G305));
  AOI22_X1  g183(.A1(new_n527), .A2(G85), .B1(new_n532), .B2(G47), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n542), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(G290));
  NAND4_X1  g190(.A1(new_n522), .A2(G92), .A3(new_n495), .A4(new_n507), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(KEYINPUT79), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n506), .A2(new_n618), .A3(G92), .A4(new_n507), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(G54), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n622));
  OAI22_X1  g197(.A1(new_n551), .A2(new_n621), .B1(new_n622), .B2(new_n542), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT10), .B1(new_n617), .B2(new_n619), .ZN(new_n624));
  NOR3_X1   g199(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g203(.A(new_n627), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n587), .B1(new_n578), .B2(new_n583), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n625), .B1(new_n634), .B2(G860), .ZN(G148));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n561), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n626), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n636), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n461), .A2(new_n470), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT80), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n468), .A2(G135), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n477), .A2(G123), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n469), .A2(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT81), .B(G2096), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n645), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G2451), .B(G2454), .Z(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  NOR2_X1   g248(.A1(G2072), .A2(G2078), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n444), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n671), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(KEYINPUT17), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n676), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n671), .B(new_n672), .C1(new_n444), .C2(new_n674), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n673), .A3(new_n671), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT85), .B(G2096), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(G1971), .B(G1976), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1956), .B(G2474), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n688), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n688), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G21), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G168), .B2(new_n705), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G1966), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(G1966), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT31), .B(G11), .Z(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT30), .B(G28), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n709), .B(new_n713), .C1(new_n711), .C2(new_n650), .ZN(new_n714));
  NOR2_X1   g289(.A1(G5), .A2(G16), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT94), .Z(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G171), .B2(G16), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n708), .B(new_n714), .C1(G1961), .C2(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n711), .A2(G35), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n711), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT29), .ZN(new_n722));
  INV_X1    g297(.A(G2090), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G34), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT24), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(KEYINPUT24), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n711), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G160), .B2(new_n711), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT91), .Z(new_n730));
  INV_X1    g305(.A(G2084), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT92), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n711), .A2(G32), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT26), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G129), .B2(new_n477), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n468), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g316(.A1(new_n730), .A2(new_n731), .B1(new_n733), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n711), .A2(G27), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT96), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G164), .B2(new_n711), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(new_n443), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n724), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n717), .A2(G1961), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n730), .A2(new_n731), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT25), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n468), .A2(KEYINPUT90), .A3(G139), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT90), .B1(new_n468), .B2(G139), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n752), .B1(new_n469), .B2(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G33), .B(new_n756), .S(G29), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2072), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n741), .A2(new_n733), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n749), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n747), .A2(new_n748), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n705), .A2(G20), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT23), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n631), .B2(new_n705), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  NOR2_X1   g343(.A1(G4), .A2(G16), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT88), .Z(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n626), .B2(new_n705), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1348), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n705), .A2(G19), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n562), .B2(new_n705), .ZN(new_n774));
  INV_X1    g349(.A(G1341), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n468), .A2(G140), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n477), .A2(G128), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n469), .A2(G116), .ZN(new_n779));
  OAI21_X1  g354(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n711), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT28), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n772), .A2(new_n776), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT89), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n719), .A2(new_n764), .A3(new_n768), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n705), .A2(G24), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G290), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT87), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(G1986), .ZN(new_n795));
  NOR2_X1   g370(.A1(G6), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n607), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT32), .ZN(new_n798));
  INV_X1    g373(.A(G1981), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n705), .A2(G22), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G166), .B2(new_n705), .ZN(new_n802));
  INV_X1    g377(.A(G1971), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  MUX2_X1   g379(.A(G23), .B(new_n596), .S(G16), .Z(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n800), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n794), .A2(G1986), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n795), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n468), .A2(G131), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n477), .A2(G119), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G29), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n711), .A2(G25), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT86), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT35), .B(G1991), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n808), .B2(KEYINPUT34), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n811), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n825), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n791), .B1(new_n827), .B2(new_n828), .ZN(G311));
  INV_X1    g404(.A(new_n828), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n790), .B1(new_n830), .B2(new_n826), .ZN(G150));
  XOR2_X1   g406(.A(KEYINPUT100), .B(G860), .Z(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n530), .B2(new_n531), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n506), .A2(G93), .A3(new_n507), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(G55), .B1(new_n549), .B2(new_n550), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n506), .A2(G93), .A3(new_n507), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(KEYINPUT98), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G67), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n520), .A2(new_n523), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g418(.A1(G80), .A2(G543), .ZN(new_n844));
  OAI21_X1  g419(.A(G651), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n832), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n625), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n849), .B(new_n851), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n559), .A2(new_n841), .A3(new_n845), .A4(new_n560), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n845), .A2(new_n841), .B1(new_n559), .B2(new_n560), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n852), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT39), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n857), .A2(KEYINPUT101), .A3(new_n832), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT101), .B1(new_n857), .B2(new_n832), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n848), .B1(new_n858), .B2(new_n859), .ZN(G145));
  INV_X1    g435(.A(KEYINPUT105), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n816), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n642), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n756), .B(new_n739), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(G164), .B(new_n781), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n477), .A2(G130), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n469), .A2(KEYINPUT103), .A3(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT103), .B1(new_n469), .B2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n869), .B(new_n870), .C1(KEYINPUT104), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(KEYINPUT104), .B2(new_n871), .ZN(new_n873));
  AOI211_X1 g448(.A(new_n868), .B(new_n873), .C1(G142), .C2(new_n468), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n866), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n865), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G160), .B(new_n650), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n876), .A2(new_n878), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n883), .B(KEYINPUT40), .Z(G395));
  INV_X1    g459(.A(new_n638), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n855), .ZN(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n626), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n631), .A2(new_n625), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(KEYINPUT106), .Z(new_n891));
  INV_X1    g466(.A(KEYINPUT107), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n584), .A2(new_n625), .A3(new_n588), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n631), .A2(new_n625), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT41), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n887), .A2(new_n896), .A3(new_n888), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n892), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT107), .B1(new_n889), .B2(KEYINPUT41), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n886), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G305), .B(new_n596), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n613), .A2(G303), .A3(new_n614), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G303), .B1(new_n613), .B2(new_n614), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n901), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT42), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n891), .A2(new_n900), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n910), .B1(new_n891), .B2(new_n900), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n841), .A2(new_n845), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n636), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(G295));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n915), .ZN(G331));
  OAI21_X1  g492(.A(G301), .B1(new_n854), .B2(new_n853), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(new_n561), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n559), .A2(new_n841), .A3(new_n845), .A4(new_n560), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(G171), .A3(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n918), .A2(G168), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G168), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n898), .A2(new_n899), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n918), .A2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(G286), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(G168), .A3(new_n921), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n887), .A3(new_n927), .A4(new_n888), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n909), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(new_n928), .ZN(new_n931));
  INV_X1    g506(.A(new_n909), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n909), .B1(new_n924), .B2(new_n928), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT108), .B1(new_n936), .B2(G37), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT43), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n926), .A2(new_n927), .B1(new_n895), .B2(new_n897), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n909), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n941), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  AND4_X1   g518(.A1(KEYINPUT43), .A2(new_n943), .A3(new_n880), .A4(new_n929), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n935), .B2(new_n937), .ZN(new_n948));
  AND4_X1   g523(.A1(new_n947), .A2(new_n943), .A3(new_n880), .A4(new_n929), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n945), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n490), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n464), .A2(new_n471), .A3(G40), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n958), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT46), .B1(new_n958), .B2(G1996), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n781), .B(new_n786), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n738), .A3(new_n737), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n959), .A2(new_n960), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n957), .A2(G1996), .A3(new_n739), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT110), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n961), .B1(G1996), .B2(new_n739), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n957), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n816), .B(new_n821), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n958), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g545(.A1(G290), .A2(G1986), .A3(new_n958), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n821), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n816), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n968), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(G2067), .B2(new_n781), .ZN(new_n979));
  AOI211_X1 g554(.A(new_n964), .B(new_n975), .C1(new_n957), .C2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n490), .A2(new_n981), .A3(new_n952), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT111), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n490), .A2(new_n984), .A3(new_n981), .A4(new_n952), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n981), .B1(new_n490), .B2(new_n952), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(new_n956), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1961), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n991));
  INV_X1    g566(.A(new_n956), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n490), .A2(KEYINPUT45), .A3(new_n952), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n955), .A2(new_n992), .A3(new_n443), .A4(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n989), .A2(new_n990), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n994), .A2(new_n991), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G171), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n989), .A2(new_n990), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT122), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1961), .B1(new_n986), .B2(new_n988), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n955), .A2(new_n992), .A3(KEYINPUT123), .A4(new_n993), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT53), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n994), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n955), .A2(new_n992), .A3(new_n993), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1008), .A2(KEYINPUT53), .A3(new_n1004), .A4(new_n443), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1000), .A2(new_n1003), .A3(new_n1006), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n998), .B1(new_n1010), .B2(G171), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT124), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(KEYINPUT124), .A3(new_n1012), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n953), .A2(KEYINPUT50), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1018), .A2(new_n956), .A3(new_n987), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT56), .B(G2072), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OAI22_X1  g596(.A1(new_n1019), .A2(G1956), .B1(new_n1007), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n584), .A2(KEYINPUT57), .A3(new_n588), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n581), .A2(new_n574), .ZN(new_n1025));
  OAI211_X1 g600(.A(KEYINPUT117), .B(new_n1024), .C1(new_n1025), .C2(new_n587), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n587), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1022), .A2(new_n1023), .A3(new_n1026), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1348), .B1(new_n986), .B2(new_n988), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n953), .A2(new_n956), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2067), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1030), .B1(new_n626), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1023), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n988), .A2(new_n982), .ZN(new_n1037));
  INV_X1    g612(.A(G1956), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n1008), .A2(new_n1020), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1034), .A2(KEYINPUT60), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT60), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1031), .A2(new_n1043), .A3(new_n1033), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n625), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1348), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n989), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1033), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(KEYINPUT60), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT120), .A3(new_n626), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT118), .B(G1996), .Z(new_n1055));
  NOR2_X1   g630(.A1(new_n956), .A2(new_n953), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(new_n775), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1007), .A2(new_n1055), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n562), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT59), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT61), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1030), .A2(new_n1040), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1030), .B2(new_n1040), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1041), .B1(new_n1054), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n594), .B(G1976), .C1(new_n595), .C2(new_n542), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT113), .B(G8), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n956), .B2(new_n953), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1072), .B(new_n1073), .C1(new_n600), .C2(G1976), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT114), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1032), .A2(new_n1076), .A3(new_n1070), .A4(new_n1067), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1077), .A3(KEYINPUT52), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  OAI21_X1  g654(.A(G1981), .B1(new_n603), .B2(new_n606), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n603), .A2(new_n606), .A3(G1981), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1082), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1071), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1074), .A2(new_n1078), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT112), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1091), .B1(G166), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT112), .ZN(new_n1094));
  NAND4_X1  g669(.A1(G303), .A2(new_n1094), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n986), .A2(new_n723), .A3(new_n988), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1007), .A2(new_n803), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1092), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1088), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1096), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(G2090), .B2(new_n1037), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1070), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1001), .B(KEYINPUT122), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1106));
  AOI21_X1  g681(.A(G301), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n997), .B2(G171), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1100), .B(new_n1104), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n986), .A2(new_n731), .A3(new_n988), .ZN(new_n1110));
  INV_X1    g685(.A(G1966), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1007), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1070), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(G168), .B2(new_n1069), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1114), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1092), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1120));
  NOR2_X1   g695(.A1(G168), .A2(new_n1069), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT51), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1069), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n1123), .B2(new_n1117), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1119), .A2(new_n1122), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1109), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1017), .A2(new_n1066), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1130), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1088), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1134));
  AOI21_X1  g709(.A(G301), .B1(new_n995), .B2(new_n996), .ZN(new_n1135));
  AND4_X1   g710(.A1(new_n1104), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1125), .A2(new_n1131), .A3(new_n1126), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1132), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(G288), .A2(G1976), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1084), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(new_n1086), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1134), .B2(new_n1088), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1123), .A2(G168), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT115), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1148), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1150), .A2(KEYINPUT63), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1100), .A3(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT116), .B(KEYINPUT63), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(new_n1154), .B2(new_n1148), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1146), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1129), .A2(new_n1141), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n1158));
  XNOR2_X1  g733(.A(G290), .B(G1986), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n970), .B1(new_n957), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n980), .B1(new_n1161), .B2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g738(.A1(new_n685), .A2(G319), .A3(new_n669), .ZN(new_n1165));
  NOR3_X1   g739(.A1(new_n883), .A2(G229), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g740(.A(new_n1166), .B1(new_n948), .B2(new_n949), .ZN(G225));
  INV_X1    g741(.A(G225), .ZN(G308));
endmodule


