//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n202), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G58), .C2(G232), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G1), .B2(G20), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G1), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n223), .A2(new_n220), .A3(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NOR3_X1   g0026(.A1(new_n218), .A2(new_n222), .A3(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n209), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G58), .ZN(new_n238));
  INV_X1    g0038(.A(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G351));
  OAI21_X1  g0045(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n246));
  INV_X1    g0046(.A(G150), .ZN(new_n247));
  NOR2_X1   g0047(.A1(G20), .A2(G33), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n220), .A2(G33), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n246), .B1(new_n247), .B2(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n221), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT65), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n223), .A2(G13), .A3(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n254), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT66), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n259), .A2(new_n260), .A3(new_n258), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n223), .A2(G20), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n261), .B(new_n262), .C1(new_n260), .C2(new_n259), .ZN(new_n263));
  MUX2_X1   g0063(.A(new_n258), .B(new_n263), .S(G50), .Z(new_n264));
  AOI21_X1  g0064(.A(KEYINPUT67), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n257), .A2(KEYINPUT67), .A3(new_n264), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G1698), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(G222), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G223), .ZN(new_n277));
  OAI221_X1 g0077(.A(new_n275), .B1(new_n239), .B2(new_n273), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n269), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n223), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G226), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n268), .A2(KEYINPUT9), .B1(G200), .B2(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n282), .A2(G190), .A3(new_n286), .A4(new_n289), .ZN(new_n292));
  XOR2_X1   g0092(.A(new_n292), .B(KEYINPUT68), .Z(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n266), .A2(new_n294), .A3(new_n267), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n291), .A2(KEYINPUT10), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n267), .ZN(new_n297));
  OAI21_X1  g0097(.A(KEYINPUT9), .B1(new_n297), .B2(new_n265), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n290), .A2(G200), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n298), .A2(new_n295), .A3(new_n293), .A4(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n290), .A2(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n257), .A2(new_n264), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n290), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n250), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n308), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT15), .B(G87), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n309), .B1(new_n251), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n258), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n311), .A2(new_n254), .B1(new_n239), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n259), .A2(G77), .A3(new_n262), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G107), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n276), .A2(new_n212), .B1(new_n316), .B2(new_n273), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n270), .A2(new_n272), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n318), .A2(new_n229), .A3(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n281), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G244), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n289), .C1(new_n321), .C2(new_n284), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n315), .B1(new_n322), .B2(G200), .ZN(new_n323));
  INV_X1    g0123(.A(G190), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n296), .A2(new_n302), .A3(new_n307), .A4(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT75), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n308), .A2(new_n312), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n263), .B2(new_n308), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G58), .A2(G68), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT72), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n331), .B(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n203), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n334), .A2(G20), .B1(G159), .B2(new_n248), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT7), .B1(new_n318), .B2(new_n220), .ZN(new_n336));
  OR2_X1    g0136(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n337));
  NAND2_X1  g0137(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(new_n269), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n272), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n336), .B1(new_n340), .B2(KEYINPUT7), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n335), .B1(new_n341), .B2(new_n202), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT16), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n259), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT70), .A2(KEYINPUT3), .ZN(new_n346));
  OAI21_X1  g0146(.A(G33), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT71), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT71), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n351), .B(G33), .C1(new_n345), .C2(new_n346), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g0155(.A(KEYINPUT7), .B(G20), .C1(new_n350), .C2(new_n352), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT16), .B(new_n335), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n330), .B1(new_n344), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n277), .A2(new_n274), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n269), .B1(new_n337), .B2(new_n338), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n352), .B(new_n359), .C1(new_n360), .C2(new_n348), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n274), .A2(G226), .ZN(new_n362));
  INV_X1    g0162(.A(G87), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n361), .A2(new_n362), .B1(new_n269), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n281), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n284), .A2(new_n229), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n365), .A2(new_n324), .A3(new_n289), .A4(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n288), .B(new_n366), .C1(new_n364), .C2(new_n281), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(G200), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n358), .A2(new_n370), .A3(KEYINPUT74), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n358), .A2(new_n370), .A3(KEYINPUT74), .A4(KEYINPUT17), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n369), .A2(G179), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n365), .A2(new_n289), .A3(new_n367), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G169), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n344), .A2(new_n357), .ZN(new_n381));
  INV_X1    g0181(.A(new_n330), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI211_X1 g0183(.A(KEYINPUT73), .B(new_n330), .C1(new_n344), .C2(new_n357), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT18), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT18), .B(new_n379), .C1(new_n383), .C2(new_n384), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n375), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n273), .A2(G226), .A3(new_n274), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n273), .A2(G232), .A3(G1698), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G33), .A2(G97), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n288), .B1(new_n393), .B2(new_n281), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n285), .A2(G238), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n394), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT14), .B1(new_n399), .B2(new_n305), .ZN(new_n400));
  INV_X1    g0200(.A(new_n398), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT14), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(G169), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n399), .A2(G179), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n400), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G50), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n249), .A2(new_n408), .B1(new_n251), .B2(new_n239), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n220), .A2(G68), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n254), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT11), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n259), .A2(G68), .A3(new_n262), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n258), .A2(G68), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n413), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n407), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n399), .A2(G190), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT69), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n403), .B2(G200), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n399), .A2(KEYINPUT69), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n418), .B(new_n421), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n322), .A2(new_n305), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n315), .C1(G179), .C2(new_n322), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n420), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n327), .A2(new_n328), .A3(new_n389), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n389), .ZN(new_n431));
  OAI21_X1  g0231(.A(KEYINPUT75), .B1(new_n431), .B2(new_n326), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n258), .A2(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n223), .A2(G33), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n258), .A2(new_n435), .A3(new_n221), .A4(new_n253), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(new_n213), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n248), .A2(G77), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT6), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n213), .A2(new_n316), .ZN(new_n440));
  NOR2_X1   g0240(.A1(G97), .A2(G107), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n316), .A2(KEYINPUT6), .A3(G97), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI221_X1 g0244(.A(new_n438), .B1(new_n220), .B2(new_n444), .C1(new_n341), .C2(new_n316), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n434), .B(new_n437), .C1(new_n445), .C2(new_n254), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G257), .A3(new_n280), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT76), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n451), .A2(new_n287), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n451), .A2(KEYINPUT76), .A3(G257), .A4(new_n280), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n454), .A2(KEYINPUT77), .A3(new_n455), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n321), .A2(G1698), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n350), .A2(new_n352), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT4), .ZN(new_n464));
  AND2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  INV_X1    g0267(.A(G250), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n466), .B(new_n467), .C1(new_n276), .C2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n281), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n461), .A2(G190), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT78), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n461), .A2(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G200), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n461), .A2(new_n470), .A3(KEYINPUT78), .A4(G190), .ZN(new_n476));
  AND4_X1   g0276(.A1(new_n446), .A2(new_n473), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G179), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n461), .A2(new_n478), .A3(new_n470), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(new_n305), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n445), .A2(new_n254), .ZN(new_n482));
  INV_X1    g0282(.A(new_n434), .ZN(new_n483));
  INV_X1    g0283(.A(new_n437), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT79), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n461), .A2(new_n470), .A3(new_n486), .A4(new_n478), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n480), .A2(new_n481), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT80), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n434), .B1(new_n445), .B2(new_n254), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n491), .A2(new_n484), .B1(new_n474), .B2(new_n305), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(KEYINPUT80), .A3(new_n480), .A4(new_n487), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n477), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n350), .A2(new_n220), .A3(G87), .A4(new_n352), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n363), .A2(G20), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n273), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT86), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n273), .A2(new_n500), .A3(new_n496), .A4(new_n497), .ZN(new_n501));
  AOI22_X1  g0301(.A1(KEYINPUT22), .A2(new_n495), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n316), .A2(KEYINPUT23), .A3(G20), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT23), .B1(new_n316), .B2(G20), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G116), .ZN(new_n506));
  OAI22_X1  g0306(.A1(new_n504), .A2(new_n505), .B1(G20), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT24), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n495), .A2(KEYINPUT22), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n499), .A2(new_n501), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT24), .ZN(new_n512));
  INV_X1    g0312(.A(new_n507), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n259), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT25), .B1(new_n312), .B2(new_n316), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n312), .A2(KEYINPUT25), .A3(new_n316), .ZN(new_n518));
  INV_X1    g0318(.A(new_n436), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n517), .A2(new_n518), .B1(G107), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G257), .A2(G1698), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n468), .B2(G1698), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n350), .A2(new_n352), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G294), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n280), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n451), .A2(G264), .A3(new_n280), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n324), .A3(new_n455), .ZN(new_n531));
  INV_X1    g0331(.A(new_n455), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n525), .A2(new_n526), .ZN(new_n533));
  OAI211_X1 g0333(.A(KEYINPUT87), .B(new_n528), .C1(new_n533), .C2(new_n280), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT87), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n527), .B2(new_n529), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n531), .B1(new_n537), .B2(G200), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n522), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n478), .B(new_n532), .C1(new_n534), .C2(new_n536), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n305), .B1(new_n530), .B2(new_n455), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n540), .A2(new_n541), .B1(new_n515), .B2(new_n521), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G238), .A2(G1698), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n321), .B2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n352), .B(new_n545), .C1(new_n360), .C2(new_n348), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n506), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n281), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n447), .A2(new_n287), .A3(G1), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n280), .B(G250), .C1(G1), .C2(new_n447), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT81), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n280), .B1(new_n546), .B2(new_n506), .ZN(new_n554));
  INV_X1    g0354(.A(new_n551), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n554), .A2(new_n549), .A3(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT81), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n553), .A2(new_n558), .A3(new_n305), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n555), .B1(new_n547), .B2(new_n281), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n557), .B1(new_n560), .B2(new_n550), .ZN(new_n561));
  NOR4_X1   g0361(.A1(new_n554), .A2(KEYINPUT81), .A3(new_n549), .A4(new_n555), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n478), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n220), .B1(new_n392), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT82), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n363), .A2(new_n213), .A3(new_n316), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n220), .C1(new_n392), .C2(new_n564), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n564), .B1(new_n251), .B2(new_n213), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n350), .A2(new_n220), .A3(new_n352), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n202), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n254), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n310), .A2(new_n312), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n310), .C2(new_n436), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n559), .A2(new_n563), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n553), .A2(new_n558), .A3(G200), .ZN(new_n578));
  OAI21_X1  g0378(.A(G190), .B1(new_n561), .B2(new_n562), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n519), .A2(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n574), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n467), .B(new_n220), .C1(G33), .C2(new_n213), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n208), .A2(G20), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n254), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT20), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n585), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n586), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n589), .A2(new_n590), .B1(new_n208), .B2(new_n312), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n519), .A2(KEYINPUT84), .A3(G116), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT84), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n436), .B2(new_n208), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT85), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT85), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n591), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT83), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n451), .A2(G270), .A3(new_n280), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n455), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n602), .B1(new_n455), .B2(new_n603), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n274), .A2(G264), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n214), .A2(new_n274), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n350), .A2(new_n352), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n318), .A2(G303), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n280), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G200), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n612), .A2(new_n604), .A3(new_n605), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G190), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n601), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n591), .A2(new_n595), .A3(new_n598), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n598), .B1(new_n591), .B2(new_n595), .ZN(new_n621));
  OAI21_X1  g0421(.A(G169), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n619), .B1(new_n622), .B2(new_n616), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n614), .A2(new_n478), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n600), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n600), .A2(new_n614), .A3(KEYINPUT21), .A4(G169), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n618), .A2(new_n623), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NOR3_X1   g0427(.A1(new_n543), .A2(new_n584), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n433), .A2(new_n494), .A3(new_n628), .ZN(G372));
  INV_X1    g0429(.A(KEYINPUT89), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n581), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n574), .A2(KEYINPUT89), .A3(new_n575), .A4(new_n580), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n552), .A2(G200), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n579), .A2(new_n631), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT88), .B1(new_n556), .B2(G169), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n552), .A2(new_n636), .A3(new_n305), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n638), .A2(new_n563), .A3(new_n576), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n542), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n494), .A2(new_n642), .A3(new_n539), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n577), .A2(new_n583), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n644), .A2(new_n490), .A3(new_n493), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n640), .A2(new_n488), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n643), .A2(new_n639), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n433), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n296), .A2(new_n302), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n420), .A2(new_n428), .ZN(new_n653));
  INV_X1    g0453(.A(new_n375), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n426), .ZN(new_n655));
  INV_X1    g0455(.A(new_n379), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(new_n358), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(new_n386), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n652), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n307), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n651), .A2(new_n661), .ZN(G369));
  INV_X1    g0462(.A(new_n543), .ZN(new_n663));
  INV_X1    g0463(.A(G13), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n223), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n663), .B1(new_n522), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n542), .B2(new_n672), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n601), .A2(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n627), .B2(new_n676), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(G330), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n641), .A2(new_n671), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n663), .A2(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n679), .B(new_n681), .C1(new_n542), .C2(new_n671), .ZN(G399));
  NAND2_X1  g0482(.A1(new_n224), .A2(new_n279), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n567), .A2(G116), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G1), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n219), .B2(new_n683), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n641), .A2(new_n689), .A3(new_n542), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n508), .A2(new_n514), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n254), .ZN(new_n692));
  INV_X1    g0492(.A(new_n536), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n527), .A2(new_n535), .A3(new_n529), .ZN(new_n694));
  OAI211_X1 g0494(.A(G179), .B(new_n455), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n541), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n692), .A2(new_n520), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT90), .B1(new_n697), .B2(new_n675), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n690), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n640), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n494), .A4(new_n539), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT26), .B1(new_n640), .B2(new_n488), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n645), .A2(KEYINPUT26), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n701), .A2(new_n639), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n688), .B1(new_n704), .B2(new_n672), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n650), .A2(new_n688), .A3(new_n672), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n628), .A2(new_n494), .A3(new_n672), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n478), .B(new_n614), .C1(new_n536), .C2(new_n534), .ZN(new_n710));
  INV_X1    g0510(.A(new_n474), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n553), .A2(new_n558), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR4_X1   g0515(.A1(new_n537), .A2(G179), .A3(new_n616), .A4(new_n556), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n474), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n711), .A4(new_n712), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n671), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n709), .A2(KEYINPUT31), .A3(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT31), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(new_n722), .A3(new_n671), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n708), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n687), .B1(new_n727), .B2(G1), .ZN(G364));
  OR2_X1    g0528(.A1(new_n678), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n678), .A2(G330), .ZN(new_n730));
  INV_X1    g0530(.A(new_n683), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n665), .A2(G45), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G1), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT91), .Z(new_n735));
  NAND3_X1  g0535(.A1(new_n729), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n350), .A2(new_n352), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n224), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT92), .ZN(new_n739));
  INV_X1    g0539(.A(new_n219), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n447), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n739), .B(new_n741), .C1(new_n447), .C2(new_n240), .ZN(new_n742));
  NAND3_X1  g0542(.A1(G355), .A2(new_n224), .A3(new_n273), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n742), .B(new_n743), .C1(G116), .C2(new_n224), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n664), .A2(new_n269), .A3(KEYINPUT93), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT93), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G13), .B2(G33), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n221), .B1(G20), .B2(new_n305), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n735), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n751), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n220), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(new_n324), .A3(G200), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(G303), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n755), .A2(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G329), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n220), .A2(new_n478), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n766), .A2(new_n324), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G322), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n318), .B(new_n764), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n765), .A2(new_n761), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI211_X1 g0572(.A(new_n760), .B(new_n770), .C1(G311), .C2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n324), .A2(G179), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n220), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G294), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n765), .A2(G200), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT94), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n324), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G326), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n780), .A2(G190), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT95), .B(G317), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT33), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n773), .A2(new_n777), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n758), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G87), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n213), .B2(new_n775), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n318), .B(new_n790), .C1(G58), .C2(new_n767), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n763), .A2(G159), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  INV_X1    g0593(.A(new_n757), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n793), .B1(G107), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G50), .A2(new_n781), .B1(new_n783), .B2(G68), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n772), .A2(G77), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n791), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n787), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n750), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n753), .B1(new_n754), .B2(new_n799), .C1(new_n678), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n736), .A2(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n315), .A2(new_n671), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n325), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n428), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n428), .A2(new_n671), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n650), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n808), .B2(new_n671), .ZN(new_n809));
  INV_X1    g0609(.A(new_n807), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n646), .A2(new_n639), .A3(new_n649), .ZN(new_n811));
  AND3_X1   g0611(.A1(new_n494), .A2(new_n642), .A3(new_n539), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n672), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n726), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n735), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n318), .B1(new_n208), .B2(new_n771), .C1(new_n768), .C2(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n775), .A2(new_n213), .B1(new_n758), .B2(new_n316), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n757), .A2(new_n363), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n762), .A2(new_n821), .ZN(new_n822));
  NOR4_X1   g0622(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n783), .ZN(new_n824));
  INV_X1    g0624(.A(new_n781), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n755), .B2(new_n824), .C1(new_n759), .C2(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n781), .A2(G137), .B1(G159), .B2(new_n772), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT96), .B(G143), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n247), .B2(new_n824), .C1(new_n768), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n794), .A2(G68), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n775), .A2(new_n201), .B1(new_n832), .B2(new_n762), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(G50), .B2(new_n788), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n830), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n826), .B1(new_n835), .B2(new_n737), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n735), .B1(new_n836), .B2(new_n751), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n748), .A2(new_n751), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n837), .B1(G77), .B2(new_n839), .C1(new_n749), .C2(new_n810), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n816), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(KEYINPUT35), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n220), .B(new_n221), .C1(new_n444), .C2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(G116), .C1(new_n842), .C2(new_n444), .ZN(new_n844));
  XNOR2_X1  g0644(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n333), .A2(new_n740), .A3(G77), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(G50), .B2(new_n202), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(G1), .A3(new_n664), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n844), .A2(new_n845), .B1(KEYINPUT98), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n845), .B2(new_n844), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(KEYINPUT98), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT99), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n420), .A2(new_n426), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n418), .A2(new_n672), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n420), .B(new_n426), .C1(new_n418), .C2(new_n672), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n807), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n721), .A2(new_n858), .A3(new_n723), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT102), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT40), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n721), .A2(new_n858), .A3(new_n723), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT102), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n358), .A2(new_n370), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n335), .B1(new_n355), .B2(new_n356), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n259), .B1(new_n866), .B2(new_n343), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT100), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n357), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n867), .B2(new_n868), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n330), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n865), .B1(new_n872), .B2(new_n669), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n656), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n669), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n383), .B2(new_n384), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n385), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT37), .B1(new_n358), .B2(new_n370), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n387), .A2(new_n388), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n654), .ZN(new_n883));
  OR2_X1    g0683(.A1(new_n872), .A2(new_n669), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT101), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT101), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n389), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n881), .C1(new_n886), .C2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n877), .B1(new_n658), .B2(new_n654), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n657), .A2(new_n865), .A3(new_n877), .ZN(new_n892));
  AOI22_X1  g0692(.A1(KEYINPUT37), .A2(new_n892), .B1(new_n878), .B2(new_n879), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n860), .A2(new_n864), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT103), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n859), .A2(KEYINPUT102), .B1(new_n889), .B2(new_n894), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT103), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(new_n899), .A3(new_n864), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n881), .B1(new_n886), .B2(new_n888), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n890), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n889), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n859), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n861), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n433), .A2(new_n725), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n907), .B(new_n908), .Z(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(G330), .ZN(new_n910));
  INV_X1    g0710(.A(new_n889), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n883), .A2(KEYINPUT101), .A3(new_n885), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n887), .B1(new_n389), .B2(new_n884), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n914), .B2(new_n881), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT39), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n889), .A2(new_n917), .A3(new_n894), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n420), .A2(new_n671), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n658), .A2(new_n876), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n856), .A2(new_n857), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n813), .A2(new_n806), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n904), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n433), .B1(new_n705), .B2(new_n707), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(new_n661), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n926), .B(new_n928), .Z(new_n929));
  XNOR2_X1  g0729(.A(new_n910), .B(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n665), .A2(new_n223), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n853), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT104), .ZN(G367));
  NOR2_X1   g0733(.A1(new_n488), .A2(new_n672), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n485), .A2(new_n671), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n934), .B1(new_n494), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n679), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n494), .A2(new_n663), .A3(new_n680), .A4(new_n935), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT42), .Z(new_n939));
  NAND2_X1  g0739(.A1(new_n490), .A2(new_n493), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n936), .B2(new_n542), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n672), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n631), .A2(new_n632), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n639), .A2(new_n944), .A3(new_n672), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n672), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n945), .B1(new_n640), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT105), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n943), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n937), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(KEYINPUT106), .Z(new_n954));
  OAI21_X1  g0754(.A(new_n681), .B1(new_n542), .B2(new_n671), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n936), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT44), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(new_n936), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(new_n679), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n681), .B1(new_n674), .B2(new_n680), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(new_n730), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n727), .B1(new_n961), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n683), .B(KEYINPUT41), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n733), .B(KEYINPUT107), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n950), .A2(new_n937), .A3(new_n952), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n954), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT108), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n954), .A2(KEYINPUT108), .A3(new_n969), .A4(new_n970), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n757), .A2(new_n239), .ZN(new_n976));
  INV_X1    g0776(.A(G137), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n273), .B1(new_n762), .B2(new_n977), .C1(new_n768), .C2(new_n247), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(G50), .C2(new_n772), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n776), .A2(G68), .B1(new_n788), .B2(G58), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(new_n825), .C2(new_n828), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G159), .B2(new_n783), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n776), .A2(G107), .B1(new_n794), .B2(G97), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G283), .A2(new_n772), .B1(new_n763), .B2(G317), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n767), .A2(G303), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n983), .A2(new_n984), .A3(new_n737), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT109), .B1(new_n758), .B2(new_n208), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n783), .A2(G294), .B1(KEYINPUT46), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(KEYINPUT46), .B2(new_n987), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n986), .B(new_n989), .C1(G311), .C2(new_n781), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n982), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n735), .B1(new_n993), .B2(new_n751), .ZN(new_n994));
  INV_X1    g0794(.A(new_n739), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n752), .B1(new_n224), .B2(new_n310), .C1(new_n995), .C2(new_n235), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n994), .B(new_n996), .C1(new_n800), .C2(new_n947), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n975), .A2(new_n997), .ZN(G387));
  AOI22_X1  g0798(.A1(new_n781), .A2(G322), .B1(G303), .B2(new_n772), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n821), .B2(new_n824), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G317), .B2(new_n767), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT48), .Z(new_n1002));
  OAI22_X1  g0802(.A1(new_n775), .A2(new_n755), .B1(new_n758), .B2(new_n817), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT111), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n763), .A2(G326), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n737), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G116), .B2(new_n794), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n762), .A2(new_n247), .ZN(new_n1011));
  INV_X1    g0811(.A(G159), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1012), .A2(new_n825), .B1(new_n824), .B2(new_n250), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n775), .A2(new_n310), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n239), .B2(new_n758), .C1(new_n213), .C2(new_n757), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1008), .B1(new_n202), .B2(new_n771), .C1(new_n408), .C2(new_n768), .ZN(new_n1016));
  OR3_X1    g0816(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1010), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n735), .B1(new_n1018), .B2(new_n751), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n250), .A2(G50), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT50), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n684), .B1(new_n202), .B2(new_n239), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g0822(.A(G45), .B(new_n1022), .C1(new_n1021), .C2(new_n1020), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n739), .B1(new_n232), .B2(new_n447), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n273), .B(new_n224), .C1(G116), .C2(new_n567), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n224), .A2(G107), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n752), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1019), .B(new_n1028), .C1(new_n674), .C2(new_n800), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT112), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n727), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(new_n963), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n683), .B1(new_n1031), .B2(new_n963), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1030), .B(new_n1034), .C1(new_n963), .C2(new_n968), .ZN(G393));
  AOI21_X1  g0835(.A(new_n683), .B1(new_n1032), .B2(new_n961), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n961), .B2(new_n1032), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n936), .A2(new_n750), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n752), .B1(new_n213), .B2(new_n224), .C1(new_n995), .C2(new_n244), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n762), .A2(new_n828), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n820), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n776), .A2(G77), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n202), .C2(new_n758), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1043), .A2(new_n737), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n408), .B2(new_n824), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT51), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n825), .A2(new_n247), .B1(new_n1012), .B2(new_n768), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n1046), .B2(new_n1047), .C1(new_n250), .C2(new_n771), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n781), .A2(G317), .B1(G311), .B2(new_n767), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT52), .Z(new_n1051));
  OAI22_X1  g0851(.A1(new_n775), .A2(new_n208), .B1(new_n757), .B2(new_n316), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n318), .B1(new_n762), .B2(new_n769), .C1(new_n817), .C2(new_n771), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(new_n783), .C2(G303), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1051), .B(new_n1054), .C1(new_n755), .C2(new_n758), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n735), .B1(new_n1056), .B2(new_n751), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1038), .A2(new_n1039), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n961), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n967), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1037), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(G390));
  NAND2_X1  g0862(.A1(new_n781), .A2(G283), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n767), .A2(G116), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n273), .B1(new_n763), .B2(G294), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1063), .A2(new_n1042), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n824), .A2(new_n316), .B1(new_n213), .B2(new_n771), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(KEYINPUT117), .B2(new_n1067), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(KEYINPUT117), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1068), .A2(new_n1069), .A3(new_n789), .A4(new_n831), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n781), .A2(G128), .B1(G132), .B2(new_n767), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT116), .Z(new_n1072));
  OR3_X1    g0872(.A1(new_n758), .A2(KEYINPUT53), .A3(new_n247), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT53), .B1(new_n758), .B2(new_n247), .ZN(new_n1074));
  XOR2_X1   g0874(.A(KEYINPUT54), .B(G143), .Z(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1073), .B(new_n1074), .C1(new_n771), .C2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G137), .B2(new_n783), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n273), .B1(new_n757), .B2(new_n408), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G125), .B2(new_n763), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT115), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1072), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n775), .A2(new_n1012), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1070), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n735), .B1(new_n1084), .B2(new_n751), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n308), .B2(new_n839), .C1(new_n919), .C2(new_n749), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n725), .A2(G330), .A3(new_n858), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n917), .B1(new_n903), .B2(new_n889), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n920), .B1(new_n924), .B2(new_n923), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n889), .A2(new_n917), .A3(new_n894), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n920), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n895), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n704), .A2(new_n672), .A3(new_n805), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n806), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1094), .B1(new_n923), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1088), .B1(new_n1092), .B2(new_n1097), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1095), .A2(new_n806), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n923), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1093), .B(new_n895), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1101), .B(new_n1087), .C1(new_n919), .C2(new_n1090), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1086), .B1(new_n1103), .B2(new_n968), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n433), .A2(new_n725), .A3(G330), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n927), .A2(new_n1106), .A3(new_n661), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n721), .A2(G330), .A3(new_n723), .A4(new_n810), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1100), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1087), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n924), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1099), .A2(new_n1087), .A3(new_n1109), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1107), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1098), .A2(new_n1102), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT113), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1098), .A2(new_n1102), .A3(new_n1113), .A4(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n683), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1113), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1103), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1121), .A2(KEYINPUT114), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(KEYINPUT114), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1105), .B1(new_n1122), .B2(new_n1123), .ZN(G378));
  AND4_X1   g0924(.A1(new_n899), .A2(new_n860), .A3(new_n864), .A4(new_n895), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n899), .B1(new_n898), .B2(new_n864), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n906), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n296), .A2(new_n302), .A3(new_n307), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n268), .A2(new_n669), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1130), .A2(KEYINPUT55), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(KEYINPUT55), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT56), .ZN(new_n1133));
  OR3_X1    g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1127), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n926), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n901), .A2(new_n1136), .A3(G330), .A4(new_n906), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1139), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1107), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(KEYINPUT121), .B1(new_n1146), .B2(new_n683), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1145), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1144), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1142), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n1152), .A3(KEYINPUT57), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT121), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n1154), .A3(new_n731), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1147), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1152), .A2(new_n967), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1076), .A2(new_n758), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n775), .A2(new_n247), .B1(new_n771), .B2(new_n977), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n781), .C2(G125), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n832), .B2(new_n824), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G128), .B2(new_n767), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G33), .B1(new_n763), .B2(G124), .ZN(new_n1165));
  AOI21_X1  g0965(.A(G41), .B1(new_n794), .B2(G159), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n279), .B1(new_n737), .B2(new_n269), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(KEYINPUT118), .A3(new_n408), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n776), .A2(G68), .B1(new_n794), .B2(G58), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n239), .B2(new_n758), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n279), .B1(new_n762), .B2(new_n755), .C1(new_n310), .C2(new_n771), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1171), .A2(new_n1008), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G97), .A2(new_n783), .B1(new_n781), .B2(G116), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n316), .C2(new_n768), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT119), .Z(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT118), .B1(new_n1168), .B2(new_n408), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1167), .A2(new_n1169), .A3(new_n1178), .A4(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n735), .B1(new_n1181), .B2(new_n751), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1182), .B1(G50), .B2(new_n839), .C1(new_n1136), .C2(new_n749), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1157), .A2(new_n1183), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1156), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(G375));
  NAND3_X1  g0986(.A1(new_n1111), .A2(new_n1107), .A3(new_n1112), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1119), .A2(new_n965), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n968), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n838), .A2(new_n202), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n923), .A2(new_n749), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G150), .A2(new_n772), .B1(new_n763), .B2(G128), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1192), .B1(new_n408), .B2(new_n775), .C1(new_n1012), .C2(new_n758), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n824), .A2(new_n1076), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(G132), .C2(new_n781), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1008), .B1(new_n201), .B2(new_n757), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT122), .Z(new_n1197));
  OAI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n977), .C2(new_n768), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n273), .B1(new_n772), .B2(G107), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n759), .B2(new_n762), .C1(new_n768), .C2(new_n755), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G97), .B2(new_n788), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n976), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(G116), .A2(new_n783), .B1(new_n781), .B2(G294), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1014), .A4(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n754), .B1(new_n1198), .B2(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1191), .A2(new_n735), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1189), .B1(new_n1190), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1188), .A2(new_n1207), .ZN(G381));
  AOI21_X1  g1008(.A(new_n1104), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(G375), .A2(new_n1210), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G381), .A2(G384), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(G407));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n670), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(G407), .A2(G213), .A3(new_n1215), .ZN(G409));
  NAND3_X1  g1016(.A1(new_n1156), .A2(G378), .A3(new_n1184), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1149), .A2(new_n965), .A3(new_n1152), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(new_n1152), .B(KEYINPUT123), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1183), .C1(new_n1219), .C2(new_n968), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(new_n1209), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n670), .A2(G213), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT60), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n683), .B1(new_n1187), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n1119), .C1(new_n1224), .C2(new_n1187), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1226), .A2(new_n1207), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1227), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1222), .A2(new_n1223), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(KEYINPUT62), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n670), .A2(G213), .A3(G2897), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1234), .B(new_n1238), .Z(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT61), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT62), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1222), .A2(new_n1242), .A3(new_n1223), .A4(new_n1234), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1236), .A2(new_n1240), .A3(new_n1241), .A4(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT126), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  XOR2_X1   g1046(.A(G393), .B(G396), .Z(new_n1247));
  AND3_X1   g1047(.A1(new_n975), .A2(new_n997), .A3(G390), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G390), .B1(new_n975), .B2(new_n997), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G387), .A2(new_n1061), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n975), .A2(new_n997), .A3(G390), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1247), .A2(KEYINPUT125), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1248), .A2(KEYINPUT125), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1250), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1257), .A2(new_n1236), .A3(KEYINPUT126), .A4(new_n1243), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1246), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1235), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT63), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1256), .A2(KEYINPUT61), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1240), .A2(KEYINPUT63), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1261), .B(new_n1262), .C1(new_n1263), .C2(new_n1260), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1259), .A2(new_n1264), .ZN(G405));
  NAND3_X1  g1065(.A1(new_n1250), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1266), .B(new_n1217), .C1(new_n1185), .C2(new_n1210), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1217), .B1(new_n1185), .B2(new_n1210), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1256), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(new_n1234), .ZN(G402));
endmodule


