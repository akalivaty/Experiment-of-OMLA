//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905;
  XNOR2_X1  g000(.A(G119), .B(G128), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT74), .ZN(new_n188));
  XOR2_X1   g002(.A(KEYINPUT24), .B(G110), .Z(new_n189));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(G119), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G128), .ZN(new_n194));
  OAI22_X1  g008(.A1(new_n192), .A2(new_n194), .B1(G119), .B2(new_n191), .ZN(new_n195));
  OAI22_X1  g009(.A1(new_n188), .A2(new_n189), .B1(G110), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT16), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n197), .A2(KEYINPUT75), .A3(G125), .ZN(new_n201));
  XNOR2_X1  g015(.A(G125), .B(G140), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n202), .B2(KEYINPUT75), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  OAI211_X1 g018(.A(G146), .B(new_n200), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n196), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n198), .A3(KEYINPUT75), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n197), .A2(KEYINPUT75), .A3(G125), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n204), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n206), .B1(new_n213), .B2(new_n199), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n205), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n188), .A2(new_n189), .B1(G110), .B2(new_n195), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT76), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n217), .B1(new_n215), .B2(new_n216), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n208), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT22), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(G137), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n208), .B(new_n224), .C1(new_n218), .C2(new_n219), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT78), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT77), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(KEYINPUT25), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT25), .B1(new_n233), .B2(KEYINPUT77), .ZN(new_n235));
  OAI22_X1  g049(.A1(new_n231), .A2(new_n234), .B1(new_n235), .B2(new_n229), .ZN(new_n236));
  INV_X1    g050(.A(G217), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(G234), .B2(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n228), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(G902), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n236), .A2(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n206), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT0), .A3(G128), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(G137), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT66), .B1(new_n256), .B2(G134), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n254), .A3(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n255), .A2(new_n257), .A3(new_n259), .A4(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT65), .B(G131), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n252), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(G143), .B2(new_n206), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n246), .B1(new_n269), .B2(new_n191), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n250), .A2(new_n268), .A3(G128), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n254), .A2(G137), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n256), .A2(G134), .ZN(new_n274));
  OAI21_X1  g088(.A(G131), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n272), .B(new_n275), .C1(new_n263), .C2(new_n261), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n252), .B(KEYINPUT67), .C1(new_n262), .C2(new_n264), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n267), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n193), .A2(G116), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n281), .B(KEYINPUT68), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT69), .B(G116), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(new_n193), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(KEYINPUT69), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(KEYINPUT69), .ZN(new_n288));
  OAI211_X1 g102(.A(KEYINPUT70), .B(G119), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT2), .B(G113), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n291), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n282), .A2(new_n285), .A3(new_n293), .A4(new_n289), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n265), .A2(new_n276), .A3(KEYINPUT30), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n280), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n298));
  INV_X1    g112(.A(G237), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n221), .A3(G210), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n298), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G101), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n265), .A2(new_n276), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n305), .A2(new_n295), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT31), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n278), .A2(new_n295), .ZN(new_n311));
  OR3_X1    g125(.A1(new_n305), .A2(new_n295), .A3(new_n309), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n303), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT31), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n297), .A2(new_n315), .A3(new_n304), .A4(new_n306), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT32), .ZN(new_n318));
  NOR2_X1   g132(.A1(G472), .A2(G902), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G472), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n313), .A2(new_n304), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n297), .A2(new_n303), .A3(new_n306), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n303), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n310), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n305), .B(new_n295), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT28), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n306), .A2(KEYINPUT73), .A3(new_n309), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n336), .A2(new_n324), .A3(new_n303), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G902), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n323), .B1(new_n330), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n242), .B1(new_n322), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n221), .A2(G952), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(G234), .B2(G237), .ZN(new_n343));
  XOR2_X1   g157(.A(KEYINPUT21), .B(G898), .Z(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(G234), .A2(G237), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G902), .A3(G953), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n343), .B1(new_n345), .B2(new_n348), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n252), .A2(new_n209), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n350), .A2(KEYINPUT88), .ZN(new_n351));
  INV_X1    g165(.A(new_n272), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n209), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(KEYINPUT88), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G224), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(G953), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT89), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT7), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n355), .A2(new_n360), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT5), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n193), .A3(G116), .ZN(new_n364));
  OAI211_X1 g178(.A(G113), .B(new_n364), .C1(new_n290), .C2(new_n363), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n294), .ZN(new_n366));
  INV_X1    g180(.A(G107), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT80), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G107), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT3), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT81), .B1(new_n367), .B2(G104), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n372), .A3(G107), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n371), .A2(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G101), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT3), .B1(new_n372), .B2(G107), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n367), .A2(G104), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n377), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n382), .B1(new_n371), .B2(G104), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G101), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n366), .B(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(G110), .B(G122), .Z(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT8), .ZN(new_n392));
  OAI22_X1  g206(.A1(new_n361), .A2(new_n362), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n393), .A2(KEYINPUT91), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n377), .A2(new_n384), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G101), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  AND4_X1   g213(.A1(new_n398), .A2(new_n395), .A3(new_n399), .A4(G101), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n378), .B1(new_n377), .B2(new_n384), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n398), .B1(new_n401), .B2(new_n399), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n295), .B(new_n397), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n389), .A2(new_n365), .A3(new_n294), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(new_n391), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n393), .B2(KEYINPUT91), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n394), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n403), .A2(new_n409), .A3(new_n404), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n403), .B2(new_n404), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n391), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(KEYINPUT87), .A2(KEYINPUT6), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n406), .A2(KEYINPUT6), .ZN(new_n415));
  INV_X1    g229(.A(new_n413), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n391), .B(new_n416), .C1(new_n410), .C2(new_n411), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n355), .B(new_n358), .Z(new_n419));
  AND3_X1   g233(.A1(new_n418), .A2(KEYINPUT90), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT90), .B1(new_n418), .B2(new_n419), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n408), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n423), .B(new_n408), .C1(new_n420), .C2(new_n421), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n349), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  INV_X1    g242(.A(G227), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(G953), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n428), .B(new_n430), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n252), .B(new_n397), .C1(new_n400), .C2(new_n402), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n262), .A2(new_n264), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n352), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(KEYINPUT1), .C1(new_n244), .C2(G146), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G128), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n246), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n271), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n385), .A3(new_n387), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n389), .A2(new_n436), .B1(new_n443), .B2(new_n435), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n433), .A2(new_n434), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n434), .B1(new_n433), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n432), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n388), .A2(new_n352), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n434), .B1(new_n449), .B2(new_n443), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n433), .A2(new_n444), .A3(new_n434), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n451), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n431), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n448), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G469), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n450), .B(KEYINPUT12), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n458), .A2(KEYINPUT84), .A3(new_n453), .A4(new_n431), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n456), .A2(new_n457), .A3(new_n227), .A4(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n458), .A2(new_n453), .A3(new_n432), .ZN(new_n461));
  INV_X1    g275(.A(new_n446), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n432), .B1(new_n462), .B2(new_n453), .ZN(new_n463));
  OAI21_X1  g277(.A(G469), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n457), .A2(new_n227), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT9), .B(G234), .Z(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G221), .B1(new_n469), .B2(G902), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n299), .A2(new_n221), .A3(G214), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(new_n244), .ZN(new_n473));
  NAND2_X1  g287(.A1(KEYINPUT18), .A2(G131), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n203), .A2(G146), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT92), .A3(new_n207), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n475), .B(new_n477), .C1(KEYINPUT92), .C2(new_n476), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(KEYINPUT17), .A3(new_n263), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n473), .B(new_n263), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(KEYINPUT17), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n478), .B1(new_n481), .B2(new_n215), .ZN(new_n482));
  XNOR2_X1  g296(.A(G113), .B(G122), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n372), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  MUX2_X1   g299(.A(new_n202), .B(new_n203), .S(KEYINPUT19), .Z(new_n486));
  OAI211_X1 g300(.A(new_n480), .B(new_n205), .C1(G146), .C2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n484), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(KEYINPUT93), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G475), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n485), .A2(new_n493), .A3(new_n227), .A4(new_n489), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n286), .A2(G122), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT95), .ZN(new_n497));
  INV_X1    g311(.A(G122), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n284), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n371), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n244), .A2(G128), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT96), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(G128), .B2(new_n244), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(G134), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(new_n284), .B2(new_n498), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT98), .Z(new_n508));
  NOR3_X1   g322(.A1(new_n284), .A2(KEYINPUT14), .A3(new_n498), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n508), .A2(new_n497), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n501), .B(new_n506), .C1(new_n510), .C2(new_n367), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n503), .A2(KEYINPUT13), .B1(G128), .B2(new_n244), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT97), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n503), .A2(KEYINPUT13), .ZN(new_n515));
  OAI221_X1 g329(.A(KEYINPUT97), .B1(G128), .B2(new_n244), .C1(new_n503), .C2(KEYINPUT13), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G134), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n500), .B(new_n371), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n518), .B(new_n519), .C1(G134), .C2(new_n505), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n469), .A2(new_n237), .A3(G953), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n511), .A2(new_n520), .A3(new_n522), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G478), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n526), .B(new_n227), .C1(KEYINPUT15), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n525), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n522), .B1(new_n511), .B2(new_n520), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n227), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT15), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(G478), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n484), .A2(KEYINPUT94), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n482), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n534), .B2(new_n482), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G475), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n495), .A2(new_n528), .A3(new_n533), .A4(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n471), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(G214), .B1(G237), .B2(G902), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT85), .ZN(new_n541));
  AND4_X1   g355(.A1(new_n341), .A2(new_n427), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n378), .ZN(G3));
  AND2_X1   g357(.A1(new_n427), .A2(new_n540), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT99), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n317), .A2(new_n227), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G472), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n236), .A2(new_n238), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n317), .A2(new_n319), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n240), .A2(new_n241), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n547), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n545), .B1(new_n551), .B2(new_n471), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n467), .A2(new_n470), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n546), .A2(G472), .B1(new_n317), .B2(new_n319), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n553), .A2(KEYINPUT99), .A3(new_n242), .A4(new_n554), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n495), .A2(new_n537), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(G478), .B1(new_n526), .B2(new_n227), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT101), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT33), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n561), .B1(new_n525), .B2(KEYINPUT100), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n526), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n526), .A2(new_n562), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(G478), .A3(new_n227), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n558), .B1(new_n560), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n544), .A2(new_n556), .A3(new_n567), .ZN(new_n568));
  XOR2_X1   g382(.A(KEYINPUT34), .B(G104), .Z(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(G6));
  NAND2_X1  g384(.A1(new_n533), .A2(new_n528), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n494), .A2(new_n491), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n494), .A2(new_n491), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n573), .A2(new_n537), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n544), .A2(new_n556), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT35), .B(G107), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G9));
  NOR2_X1   g396(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n220), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n241), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n548), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n554), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n427), .A2(new_n539), .A3(new_n541), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT37), .B(G110), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G12));
  INV_X1    g408(.A(G900), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n343), .B1(new_n348), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n572), .A2(new_n576), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n418), .A2(new_n419), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n418), .A2(KEYINPUT90), .A3(new_n419), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n423), .B1(new_n602), .B2(new_n408), .ZN(new_n603));
  INV_X1    g417(.A(new_n426), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n540), .B(new_n597), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT106), .ZN(new_n606));
  INV_X1    g420(.A(new_n321), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n330), .A2(new_n338), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n612), .A2(new_n553), .A3(new_n586), .ZN(new_n613));
  INV_X1    g427(.A(new_n540), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n425), .B2(new_n426), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT106), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n597), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n606), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  XOR2_X1   g433(.A(new_n596), .B(KEYINPUT39), .Z(new_n620));
  NAND2_X1  g434(.A1(new_n553), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT40), .Z(new_n622));
  NAND2_X1  g436(.A1(new_n297), .A2(new_n306), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n304), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n227), .B1(new_n333), .B2(new_n304), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n609), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n622), .A2(new_n540), .A3(new_n587), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n425), .A2(new_n426), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT38), .Z(new_n631));
  OR4_X1    g445(.A1(new_n572), .A2(new_n629), .A3(new_n558), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT107), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G143), .ZN(G45));
  INV_X1    g448(.A(new_n596), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n567), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n613), .A3(new_n615), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G146), .ZN(G48));
  NAND3_X1  g452(.A1(new_n456), .A2(new_n227), .A3(new_n459), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT108), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n456), .A2(KEYINPUT108), .A3(new_n227), .A4(new_n459), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n641), .A2(G469), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n460), .A2(KEYINPUT109), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n641), .A2(KEYINPUT109), .A3(G469), .A4(new_n642), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(new_n470), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(new_n340), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n648), .A2(new_n427), .A3(new_n540), .A4(new_n567), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT41), .B(G113), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G15));
  NAND4_X1  g465(.A1(new_n648), .A2(new_n427), .A3(new_n540), .A4(new_n577), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G116), .ZN(G18));
  AOI211_X1 g467(.A(new_n349), .B(new_n538), .C1(new_n609), .C2(new_n611), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n645), .A2(new_n470), .A3(new_n646), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n615), .A2(new_n654), .A3(new_n586), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G119), .ZN(G21));
  AND3_X1   g471(.A1(new_n655), .A2(new_n630), .A3(new_n540), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n558), .A2(new_n572), .ZN(new_n659));
  INV_X1    g473(.A(new_n242), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n336), .A2(new_n303), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n308), .A3(new_n316), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n319), .B(KEYINPUT110), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n547), .A2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n660), .A2(new_n665), .A3(new_n349), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n658), .A2(KEYINPUT111), .A3(new_n659), .A4(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n615), .A2(new_n659), .A3(new_n655), .A4(new_n666), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT111), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G122), .ZN(G24));
  INV_X1    g486(.A(new_n665), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n658), .A2(new_n586), .A3(new_n636), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G125), .ZN(G27));
  NAND4_X1  g489(.A1(new_n425), .A2(new_n470), .A3(new_n540), .A4(new_n426), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n464), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n464), .A2(new_n678), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n460), .A3(new_n466), .A4(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n677), .A2(new_n341), .A3(new_n636), .A4(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n567), .A2(new_n635), .ZN(new_n684));
  INV_X1    g498(.A(new_n681), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n676), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n340), .A2(KEYINPUT113), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n612), .A2(new_n688), .A3(new_n242), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n687), .A2(new_n689), .A3(KEYINPUT42), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n682), .A2(new_n683), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(G131), .Z(G33));
  NAND4_X1  g506(.A1(new_n677), .A2(new_n341), .A3(new_n597), .A4(new_n681), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G134), .ZN(G36));
  NOR2_X1   g508(.A1(new_n461), .A2(new_n463), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT114), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT114), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n696), .A2(new_n699), .A3(G469), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n466), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n460), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n702), .A2(new_n703), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n470), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n560), .A2(new_n566), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n558), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT43), .B1(new_n558), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n588), .A3(new_n586), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n708), .B(new_n620), .C1(new_n709), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n709), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n630), .A2(new_n614), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G137), .ZN(G39));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n707), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT47), .B(new_n470), .C1(new_n705), .C2(new_n706), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n684), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n612), .A2(new_n242), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n718), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G140), .ZN(G42));
  NAND2_X1  g542(.A1(new_n645), .A2(new_n646), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n729), .B(KEYINPUT116), .Z(new_n730));
  INV_X1    g544(.A(new_n470), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n723), .A2(new_n724), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n660), .A2(new_n665), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n714), .A2(new_n343), .A3(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n718), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n614), .A3(new_n631), .A4(new_n655), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT50), .ZN(new_n739));
  AND4_X1   g553(.A1(new_n343), .A2(new_n714), .A3(new_n655), .A4(new_n718), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n587), .A2(new_n665), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n738), .A2(KEYINPUT50), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n628), .A2(new_n660), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n718), .A2(new_n343), .A3(new_n655), .A4(new_n743), .ZN(new_n744));
  OR3_X1    g558(.A1(new_n744), .A2(new_n557), .A3(new_n710), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n737), .A2(new_n739), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n747), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n748), .A2(new_n750), .A3(new_n342), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n685), .A2(new_n731), .A3(new_n586), .A4(new_n596), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n752), .A2(new_n615), .A3(new_n659), .A4(new_n628), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n674), .A2(new_n618), .A3(new_n637), .A4(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n558), .A2(new_n571), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n556), .A2(new_n541), .A3(new_n427), .A4(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n759), .A2(KEYINPUT117), .A3(new_n590), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT117), .B1(new_n759), .B2(new_n590), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n649), .A2(new_n652), .A3(new_n656), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n349), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n541), .B(new_n765), .C1(new_n603), .C2(new_n604), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n552), .A2(new_n555), .ZN(new_n767));
  INV_X1    g581(.A(new_n567), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n542), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n671), .A2(new_n764), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n762), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n677), .A2(new_n636), .A3(new_n681), .A4(new_n741), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n571), .A2(new_n596), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n718), .A2(new_n575), .A3(new_n613), .A4(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n693), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n691), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n756), .A2(KEYINPUT53), .A3(new_n772), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n618), .A2(new_n637), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n755), .A3(new_n674), .A4(new_n753), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n754), .A2(KEYINPUT52), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n784));
  INV_X1    g598(.A(new_n590), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n766), .A2(new_n767), .A3(new_n757), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n759), .A2(KEYINPUT117), .A3(new_n590), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n763), .B1(new_n670), .B2(new_n667), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n777), .A2(new_n789), .A3(new_n790), .A4(new_n770), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n779), .B1(new_n783), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n778), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n783), .A2(new_n791), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(KEYINPUT118), .A3(KEYINPUT53), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT54), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n778), .B2(new_n792), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n744), .A2(new_n768), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n736), .A2(new_n658), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n751), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n687), .A2(new_n689), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n740), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT48), .Z(new_n806));
  OAI22_X1  g620(.A1(new_n803), .A2(new_n806), .B1(G952), .B2(G953), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n730), .B(KEYINPUT49), .ZN(new_n808));
  AND4_X1   g622(.A1(new_n470), .A2(new_n808), .A3(new_n541), .A4(new_n631), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(new_n558), .A3(new_n710), .A4(new_n743), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n807), .A2(new_n810), .ZN(G75));
  NOR2_X1   g625(.A1(new_n221), .A2(G952), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n418), .B(new_n419), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT55), .Z(new_n814));
  NAND4_X1  g628(.A1(new_n794), .A2(G210), .A3(G902), .A4(new_n796), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n794), .A2(G902), .A3(new_n796), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n794), .A2(KEYINPUT120), .A3(G902), .A4(new_n796), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n424), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n814), .A2(new_n816), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n812), .B(new_n817), .C1(new_n823), .C2(new_n824), .ZN(G51));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n794), .A2(new_n796), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n798), .ZN(new_n828));
  INV_X1    g642(.A(new_n797), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n794), .A2(KEYINPUT121), .A3(KEYINPUT54), .A4(new_n796), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n465), .B(KEYINPUT57), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n456), .A2(new_n459), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT122), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n822), .A2(new_n700), .A3(new_n698), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n812), .B1(new_n836), .B2(new_n837), .ZN(G54));
  AND2_X1   g652(.A1(KEYINPUT58), .A2(G475), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n820), .A2(new_n821), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n485), .A2(new_n489), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n812), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT123), .B1(new_n840), .B2(new_n841), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n846));
  INV_X1    g660(.A(new_n841), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n822), .A2(new_n846), .A3(new_n847), .A4(new_n839), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n845), .B2(new_n848), .ZN(G60));
  NAND2_X1  g663(.A1(G478), .A2(G902), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT59), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n831), .A2(new_n565), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n797), .B2(new_n799), .ZN(new_n853));
  INV_X1    g667(.A(new_n565), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n812), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n852), .A2(new_n855), .ZN(G63));
  NAND2_X1  g670(.A1(G217), .A2(G902), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT60), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n827), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n812), .B1(new_n859), .B2(new_n239), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n827), .A2(new_n858), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n584), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT61), .B1(new_n862), .B2(KEYINPUT124), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n860), .B(new_n862), .C1(KEYINPUT124), .C2(KEYINPUT61), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(G66));
  OAI21_X1  g681(.A(G953), .B1(new_n345), .B2(new_n356), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(new_n772), .B2(G953), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT125), .ZN(new_n870));
  INV_X1    g684(.A(new_n418), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(G898), .B2(new_n221), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n870), .B(new_n872), .ZN(G69));
  NAND3_X1  g687(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n280), .A2(new_n296), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n486), .ZN(new_n876));
  AOI211_X1 g690(.A(new_n340), .B(new_n621), .C1(new_n768), .C2(new_n757), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n718), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n716), .B2(new_n719), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT126), .Z(new_n880));
  AND2_X1   g694(.A1(new_n780), .A2(new_n674), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n632), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT62), .Z(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n727), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n874), .B(new_n876), .C1(new_n884), .C2(G953), .ZN(new_n885));
  INV_X1    g699(.A(new_n691), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n727), .A2(new_n886), .A3(new_n693), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n615), .A2(new_n659), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n708), .A2(new_n620), .A3(new_n804), .A4(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n887), .A2(new_n720), .A3(new_n881), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n221), .ZN(new_n891));
  INV_X1    g705(.A(new_n876), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n429), .A2(G900), .A3(G953), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n885), .A2(new_n894), .ZN(G72));
  NAND2_X1  g709(.A1(G472), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT63), .Z(new_n897));
  INV_X1    g711(.A(new_n772), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(new_n890), .B2(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n327), .B(KEYINPUT127), .Z(new_n900));
  AOI21_X1  g714(.A(new_n812), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n778), .A2(new_n792), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n902), .A2(new_n327), .A3(new_n624), .A4(new_n897), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n897), .B1(new_n884), .B2(new_n898), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n625), .B2(new_n905), .ZN(G57));
endmodule


