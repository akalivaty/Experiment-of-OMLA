//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT74), .B(G211gat), .ZN(new_n203));
  AOI21_X1  g002(.A(KEYINPUT22), .B1(new_n203), .B2(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  OAI22_X1  g009(.A1(new_n205), .A2(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT75), .B1(new_n204), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G211gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT74), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT74), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G211gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n216), .A3(G218gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT22), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT75), .ZN(new_n220));
  INV_X1    g019(.A(new_n205), .ZN(new_n221));
  INV_X1    g020(.A(G218gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n221), .A2(new_n206), .B1(new_n223), .B2(new_n208), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n219), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n212), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n219), .B1(new_n205), .B2(new_n207), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n223), .A3(new_n208), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G226gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n233));
  AND2_X1   g032(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n234));
  AND2_X1   g033(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n236));
  OAI22_X1  g035(.A1(new_n233), .A2(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT28), .ZN(new_n238));
  NOR2_X1   g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT26), .ZN(new_n240));
  NAND2_X1  g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n239), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT66), .B(G190gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT27), .B(G183gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n238), .A2(new_n242), .A3(new_n243), .A4(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  INV_X1    g048(.A(G183gat), .ZN(new_n250));
  INV_X1    g049(.A(G190gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT25), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT23), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT23), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n255), .A2(new_n257), .A3(new_n241), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n255), .A2(new_n241), .A3(new_n257), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n244), .A2(new_n250), .B1(KEYINPUT65), .B2(new_n249), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n253), .B1(new_n249), .B2(KEYINPUT65), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT25), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n248), .B(new_n259), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n232), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n250), .B1(new_n234), .B2(new_n233), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n258), .B1(new_n271), .B2(new_n262), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(KEYINPUT25), .B1(new_n258), .B2(new_n254), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n231), .B1(new_n273), .B2(new_n248), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n230), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n266), .A2(new_n232), .ZN(new_n276));
  AOI21_X1  g075(.A(KEYINPUT29), .B1(new_n273), .B2(new_n248), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n229), .B(new_n276), .C1(new_n277), .C2(new_n232), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n275), .A2(KEYINPUT76), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT76), .B1(new_n275), .B2(new_n278), .ZN(new_n280));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT77), .ZN(new_n282));
  XNOR2_X1  g081(.A(G64gat), .B(G92gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT78), .ZN(new_n285));
  OR3_X1    g084(.A1(new_n279), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n275), .A2(new_n278), .ZN(new_n288));
  INV_X1    g087(.A(new_n284), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n275), .A2(new_n278), .A3(KEYINPUT30), .A4(new_n284), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OR3_X1    g091(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  INV_X1    g093(.A(G148gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G141gat), .ZN(new_n296));
  INV_X1    g095(.A(G141gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G148gat), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n293), .A2(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n297), .A2(G148gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n295), .A2(G141gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n296), .A2(new_n298), .A3(KEYINPUT79), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  XOR2_X1   g105(.A(G155gat), .B(G162gat), .Z(new_n307));
  AOI21_X1  g106(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G113gat), .ZN(new_n309));
  OR3_X1    g108(.A1(new_n309), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n310));
  INV_X1    g109(.A(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G113gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(G120gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G127gat), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n315), .A2(new_n316), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n309), .A2(G120gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n311), .A2(G113gat), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT69), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n312), .A2(new_n314), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n316), .A3(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n318), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n320), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n317), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n319), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n329), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n327), .A2(KEYINPUT70), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT70), .B1(new_n327), .B2(new_n334), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n308), .B(new_n321), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n327), .A2(new_n334), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n327), .A2(KEYINPUT70), .A3(new_n334), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n308), .A4(new_n321), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n306), .A2(new_n307), .ZN(new_n348));
  INV_X1    g147(.A(new_n299), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI211_X1 g149(.A(KEYINPUT80), .B(new_n299), .C1(new_n306), .C2(new_n307), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(new_n321), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n308), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT82), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n346), .A2(new_n357), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n350), .A2(new_n351), .ZN(new_n363));
  INV_X1    g162(.A(new_n321), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n341), .B2(new_n342), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n337), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n366), .B2(new_n359), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(G57gat), .B(G85gat), .Z(new_n369));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n346), .A2(new_n357), .A3(new_n362), .A4(new_n360), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT6), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n368), .A2(new_n374), .ZN(new_n379));
  INV_X1    g178(.A(new_n373), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n379), .A2(KEYINPUT84), .A3(new_n380), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n378), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n386));
  AOI211_X1 g185(.A(new_n202), .B(new_n292), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G15gat), .B(G43gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  OR2_X1    g189(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(KEYINPUT72), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(KEYINPUT33), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n353), .A2(new_n266), .ZN(new_n394));
  INV_X1    g193(.A(new_n266), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n365), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT64), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT32), .B(new_n393), .C1(new_n397), .C2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n394), .B2(new_n396), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT33), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT32), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n390), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n399), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(KEYINPUT34), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n397), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n394), .A2(new_n396), .A3(new_n398), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n400), .A2(new_n404), .A3(new_n410), .A4(new_n408), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(KEYINPUT31), .B(G50gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n212), .A2(new_n419), .A3(new_n225), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n228), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n212), .B2(new_n225), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n267), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n355), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT86), .ZN(new_n425));
  INV_X1    g224(.A(new_n308), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n204), .A2(new_n211), .A3(KEYINPUT75), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n220), .B1(new_n219), .B2(new_n224), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT85), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n228), .A3(new_n420), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n354), .B1(new_n431), .B2(new_n267), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT86), .B1(new_n432), .B2(new_n308), .ZN(new_n433));
  NAND2_X1  g232(.A1(G228gat), .A2(G233gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n356), .A2(new_n267), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n230), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n427), .A2(new_n433), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT3), .B1(new_n229), .B2(new_n267), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(new_n363), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(G228gat), .A3(G233gat), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n437), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n438), .B1(new_n437), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n418), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n434), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n308), .B1(new_n423), .B2(new_n355), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n436), .B1(new_n446), .B2(new_n425), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n441), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G22gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n437), .A2(new_n438), .A3(new_n441), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n417), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n414), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n379), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n368), .A2(KEYINPUT87), .A3(new_n374), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n373), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n386), .B1(new_n456), .B2(new_n377), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n444), .A2(new_n451), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT73), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n412), .A2(new_n459), .A3(new_n413), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n411), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n292), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n457), .A2(new_n458), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n387), .A2(new_n452), .B1(new_n464), .B2(new_n202), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n368), .A2(KEYINPUT87), .A3(new_n374), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT87), .B1(new_n368), .B2(new_n374), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n380), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n378), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n275), .A2(new_n278), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n275), .A2(new_n278), .A3(new_n474), .A4(new_n471), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n279), .A2(new_n280), .A3(new_n471), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT38), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n289), .B1(new_n288), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n471), .B1(new_n275), .B2(new_n278), .ZN(new_n481));
  AOI211_X1 g280(.A(KEYINPUT38), .B(new_n481), .C1(new_n473), .C2(new_n475), .ZN(new_n482));
  INV_X1    g281(.A(new_n285), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n470), .A2(new_n386), .A3(new_n478), .A4(new_n484), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n366), .A2(new_n359), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n360), .B1(new_n346), .B2(new_n357), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n488), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n373), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  OR3_X1    g292(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n493), .B1(new_n490), .B2(new_n492), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n495), .A3(new_n292), .A4(new_n469), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n485), .A2(new_n458), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g296(.A1(new_n444), .A2(new_n451), .ZN(new_n498));
  INV_X1    g297(.A(new_n386), .ZN(new_n499));
  AOI211_X1 g298(.A(new_n382), .B(new_n373), .C1(new_n368), .C2(new_n374), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(new_n377), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n499), .B1(new_n501), .B2(new_n383), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n498), .B1(new_n502), .B2(new_n292), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n412), .A2(KEYINPUT36), .A3(new_n413), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n462), .B2(KEYINPUT36), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n497), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n465), .A2(new_n466), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n466), .B1(new_n465), .B2(new_n506), .ZN(new_n508));
  XNOR2_X1  g307(.A(G127gat), .B(G155gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(G231gat), .A2(G233gat), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g315(.A1(G71gat), .A2(G78gat), .ZN(new_n517));
  OR2_X1    g316(.A1(G71gat), .A2(G78gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n517), .B(new_n518), .C1(new_n515), .C2(new_n519), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT92), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT21), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529));
  XNOR2_X1  g328(.A(G15gat), .B(G22gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(G1gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G1gat), .B2(new_n530), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G8gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n528), .A2(new_n529), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n529), .B1(new_n528), .B2(new_n535), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n514), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n523), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n541));
  XOR2_X1   g340(.A(G183gat), .B(G211gat), .Z(new_n542));
  XOR2_X1   g341(.A(new_n541), .B(new_n542), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n535), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT93), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(new_n536), .A3(new_n513), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n539), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n544), .B1(new_n539), .B2(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n512), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n539), .A2(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n543), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n511), .A3(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT95), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n559), .A2(G85gat), .A3(G92gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n560), .A3(KEYINPUT7), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G99gat), .B(G106gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n570), .A2(KEYINPUT96), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(KEYINPUT96), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n565), .B(new_n566), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n564), .B(new_n563), .C1(new_n571), .C2(new_n572), .ZN(new_n574));
  INV_X1    g373(.A(new_n566), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n576), .A3(KEYINPUT97), .ZN(new_n577));
  OR3_X1    g376(.A1(new_n574), .A2(KEYINPUT97), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OR3_X1    g378(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n580), .A2(new_n581), .B1(G29gat), .B2(G36gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT15), .ZN(new_n583));
  XOR2_X1   g382(.A(G43gat), .B(G50gat), .Z(new_n584));
  OR3_X1    g383(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n583), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n583), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT17), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT17), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n579), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n579), .B2(new_n589), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n594), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n594), .B2(new_n596), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT94), .ZN(new_n602));
  XOR2_X1   g401(.A(G134gat), .B(G162gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OR3_X1    g404(.A1(new_n599), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n605), .B1(new_n599), .B2(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n556), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G230gat), .ZN(new_n610));
  INV_X1    g409(.A(G233gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n577), .A2(new_n578), .A3(new_n523), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n540), .A2(new_n573), .A3(new_n576), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n579), .A2(KEYINPUT10), .A3(new_n527), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n612), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n619), .A2(new_n621), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n609), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n507), .A2(new_n508), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n534), .A2(new_n589), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n593), .B2(new_n534), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT18), .ZN(new_n635));
  NAND2_X1  g434(.A1(G229gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n635), .B1(new_n634), .B2(new_n637), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n534), .B(new_n589), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n636), .B(KEYINPUT13), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n644));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G169gat), .B(G197gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n638), .A2(new_n642), .A3(new_n639), .A4(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n632), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n502), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g456(.A1(new_n654), .A2(new_n463), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT98), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n654), .B2(new_n463), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  OAI211_X1 g461(.A(new_n659), .B(new_n661), .C1(KEYINPUT42), .C2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n663), .B1(new_n664), .B2(G8gat), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n658), .A2(KEYINPUT42), .A3(new_n662), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(G1325gat));
  AOI21_X1  g466(.A(G15gat), .B1(new_n655), .B2(new_n462), .ZN(new_n668));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n505), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT99), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n668), .B1(new_n655), .B2(new_n671), .ZN(G1326gat));
  NOR2_X1   g471(.A1(new_n654), .A2(new_n458), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676));
  INV_X1    g475(.A(new_n608), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n292), .B1(new_n385), .B2(new_n386), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n680), .B1(new_n681), .B2(new_n458), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n498), .B(KEYINPUT101), .C1(new_n502), .C2(new_n292), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n682), .A2(new_n497), .A3(new_n683), .A4(new_n505), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n677), .B(new_n679), .C1(new_n684), .C2(new_n465), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n497), .A2(new_n503), .A3(new_n505), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n464), .A2(new_n202), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n681), .A2(KEYINPUT35), .A3(new_n452), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT89), .B1(new_n686), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n465), .A2(new_n506), .A3(new_n466), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n608), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n685), .B1(new_n692), .B2(KEYINPUT44), .ZN(new_n693));
  INV_X1    g492(.A(new_n653), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n555), .B(KEYINPUT100), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n630), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n502), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n676), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(KEYINPUT103), .A3(new_n502), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(G29gat), .A3(new_n701), .ZN(new_n702));
  NOR4_X1   g501(.A1(new_n692), .A2(new_n694), .A3(new_n555), .A4(new_n629), .ZN(new_n703));
  INV_X1    g502(.A(G29gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n502), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(G1328gat));
  INV_X1    g506(.A(G36gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n703), .A2(new_n708), .A3(new_n292), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n698), .B2(new_n463), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(G43gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n703), .A2(new_n713), .A3(new_n462), .ZN(new_n714));
  NOR4_X1   g513(.A1(new_n693), .A2(new_n694), .A3(new_n505), .A4(new_n696), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n715), .B2(new_n713), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI221_X1 g519(.A(new_n714), .B1(new_n717), .B2(KEYINPUT47), .C1(new_n715), .C2(new_n713), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1330gat));
  NAND3_X1  g521(.A1(new_n697), .A2(G50gat), .A3(new_n498), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n703), .A2(new_n498), .ZN(new_n724));
  INV_X1    g523(.A(G50gat), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT48), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n723), .A2(new_n729), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n684), .A2(new_n465), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n609), .A2(new_n629), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n694), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n732), .A2(KEYINPUT105), .A3(new_n694), .A4(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n502), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g541(.A1(new_n739), .A2(new_n463), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n743), .B2(new_n744), .ZN(G1333gat));
  INV_X1    g546(.A(new_n462), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT106), .B1(new_n739), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(G71gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n737), .A2(new_n751), .A3(new_n462), .A4(new_n738), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  OR3_X1    g552(.A1(new_n739), .A2(new_n750), .A3(new_n505), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n498), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G78gat), .ZN(G1335gat));
  INV_X1    g558(.A(new_n685), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n507), .A2(new_n508), .A3(new_n677), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n555), .A2(new_n653), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n629), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n699), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n732), .A2(new_n608), .A3(new_n764), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n732), .A2(KEYINPUT51), .A3(new_n608), .A4(new_n764), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(KEYINPUT108), .A3(new_n772), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n775), .A2(new_n568), .A3(new_n629), .A4(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n768), .B1(new_n699), .B2(new_n777), .ZN(G1336gat));
  NAND3_X1  g577(.A1(new_n629), .A2(new_n292), .A3(new_n569), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(KEYINPUT110), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(KEYINPUT110), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n463), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n569), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  OAI221_X1 g587(.A(new_n782), .B1(new_n786), .B2(new_n785), .C1(new_n783), .C2(new_n569), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n767), .B2(new_n505), .ZN(new_n791));
  INV_X1    g590(.A(G99gat), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n775), .A2(new_n792), .A3(new_n629), .A4(new_n776), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n748), .B2(new_n793), .ZN(G1338gat));
  NOR3_X1   g593(.A1(new_n458), .A2(new_n630), .A3(G106gat), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n771), .B2(new_n772), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT113), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n693), .A2(new_n458), .A3(new_n765), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n804), .B(new_n805), .C1(new_n771), .C2(new_n772), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n763), .A2(new_n498), .A3(new_n766), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(G106gat), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n808), .A2(new_n809), .A3(new_n799), .ZN(new_n810));
  INV_X1    g609(.A(new_n805), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n773), .A2(new_n803), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n801), .B2(new_n800), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT112), .B1(new_n813), .B2(KEYINPUT53), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n802), .B1(new_n810), .B2(new_n814), .ZN(G1339gat));
  NAND2_X1  g614(.A1(new_n502), .A2(new_n463), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n616), .A2(new_n612), .A3(new_n617), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n619), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n618), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(new_n820), .B2(new_n625), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n822));
  AOI211_X1 g621(.A(new_n822), .B(new_n627), .C1(new_n618), .C2(new_n819), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n818), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(KEYINPUT55), .B(new_n818), .C1(new_n821), .C2(new_n823), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n826), .A2(new_n653), .A3(new_n628), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n634), .A2(new_n829), .A3(new_n637), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n640), .A2(new_n641), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n829), .B1(new_n634), .B2(new_n637), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n652), .B1(new_n833), .B2(new_n648), .ZN(new_n834));
  OR2_X1    g633(.A1(new_n630), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n608), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n606), .B2(new_n607), .ZN(new_n837));
  AND4_X1   g636(.A1(new_n628), .A2(new_n837), .A3(new_n826), .A4(new_n827), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n695), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n609), .A2(new_n694), .A3(new_n630), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n816), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n452), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n842), .A2(new_n309), .A3(new_n653), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n748), .A2(new_n498), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n694), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(G1340gat));
  NAND2_X1  g646(.A1(new_n629), .A2(new_n311), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT117), .Z(new_n849));
  NAND2_X1  g648(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n841), .A2(new_n629), .A3(new_n844), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n851), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT116), .B1(new_n851), .B2(G120gat), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT118), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n842), .A2(new_n317), .A3(new_n555), .ZN(new_n856));
  OAI21_X1  g655(.A(G127gat), .B1(new_n845), .B2(new_n695), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT119), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n319), .A3(new_n608), .ZN(new_n860));
  XOR2_X1   g659(.A(new_n860), .B(KEYINPUT56), .Z(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n845), .B2(new_n677), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1343gat));
  OAI21_X1  g662(.A(new_n556), .B1(new_n836), .B2(new_n838), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n840), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(KEYINPUT57), .A3(new_n498), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n458), .B1(new_n839), .B2(new_n840), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n866), .B(KEYINPUT120), .C1(KEYINPUT57), .C2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n816), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n505), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  AOI211_X1 g670(.A(new_n871), .B(new_n458), .C1(new_n864), .C2(new_n840), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G141gat), .B1(new_n875), .B2(new_n694), .ZN(new_n876));
  INV_X1    g675(.A(new_n870), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n867), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(new_n297), .A3(new_n653), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n295), .A3(new_n629), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n865), .B2(new_n498), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n871), .B(new_n458), .C1(new_n839), .C2(new_n840), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n629), .B(new_n877), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(G148gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT121), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT59), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n875), .A2(new_n630), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(KEYINPUT59), .A3(new_n295), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n883), .B1(new_n892), .B2(new_n894), .ZN(G1345gat));
  AOI21_X1  g694(.A(G155gat), .B1(new_n879), .B2(new_n555), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n875), .A2(new_n695), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(G155gat), .ZN(G1346gat));
  NOR3_X1   g697(.A1(new_n878), .A2(G162gat), .A3(new_n677), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n868), .A2(new_n874), .A3(new_n608), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(G162gat), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT122), .ZN(G1347gat));
  AOI21_X1  g701(.A(new_n502), .B1(new_n839), .B2(new_n840), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI211_X1 g704(.A(KEYINPUT123), .B(new_n502), .C1(new_n839), .C2(new_n840), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n452), .A2(new_n292), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT124), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(G169gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n653), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n903), .A2(new_n292), .A3(new_n844), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n694), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n909), .B2(new_n629), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n912), .A2(new_n630), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(G176gat), .B2(new_n916), .ZN(G1349gat));
  NAND2_X1  g716(.A1(new_n839), .A2(new_n840), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n699), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n904), .ZN(new_n921));
  INV_X1    g720(.A(new_n908), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n920), .A2(new_n245), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT125), .B1(new_n923), .B2(new_n556), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n925), .A3(new_n245), .A4(new_n555), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G183gat), .B1(new_n912), .B2(new_n695), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT60), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT60), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(G1350gat));
  OAI21_X1  g732(.A(G190gat), .B1(new_n912), .B2(new_n677), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT61), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n909), .A2(new_n244), .A3(new_n608), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n905), .A2(new_n906), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n458), .A2(new_n463), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n505), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(KEYINPUT126), .B(G197gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n653), .A3(new_n942), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n884), .A2(new_n885), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n944), .A2(new_n699), .A3(new_n292), .A4(new_n505), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n694), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n946), .B2(new_n942), .ZN(G1352gat));
  OAI21_X1  g746(.A(KEYINPUT127), .B1(new_n945), .B2(new_n630), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n292), .B(new_n505), .C1(new_n884), .C2(new_n885), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  NAND4_X1  g750(.A1(new_n950), .A2(new_n951), .A3(new_n699), .A4(new_n629), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(G204gat), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n940), .A2(G204gat), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT62), .B1(new_n954), .B2(new_n630), .ZN(new_n955));
  OR4_X1    g754(.A1(KEYINPUT62), .A2(new_n940), .A3(G204gat), .A4(new_n630), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G1353gat));
  OR3_X1    g756(.A1(new_n940), .A2(new_n203), .A3(new_n556), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n950), .A2(new_n699), .A3(new_n555), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n959), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n959), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(G218gat), .B1(new_n945), .B2(new_n677), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n941), .A2(new_n222), .A3(new_n608), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1355gat));
endmodule


