//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G211gat), .ZN(new_n203));
  INV_X1    g002(.A(G218gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G211gat), .A2(G218gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(KEYINPUT70), .A3(new_n206), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT71), .ZN(new_n212));
  INV_X1    g011(.A(G197gat), .ZN(new_n213));
  INV_X1    g012(.A(G204gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G197gat), .A2(G204gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n206), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n211), .A2(new_n212), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n209), .B(new_n210), .C1(new_n218), .C2(KEYINPUT71), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT79), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT2), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(new_n227), .B2(new_n226), .ZN(new_n229));
  INV_X1    g028(.A(G155gat), .ZN(new_n230));
  INV_X1    g029(.A(G162gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n230), .A2(new_n231), .A3(KEYINPUT78), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n233), .B1(G155gat), .B2(G162gat), .ZN(new_n234));
  AOI22_X1  g033(.A1(new_n232), .A2(new_n234), .B1(G155gat), .B2(G162gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n226), .B(KEYINPUT80), .ZN(new_n237));
  NAND2_X1  g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT81), .B1(new_n238), .B2(KEYINPUT2), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n230), .A3(new_n231), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n236), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT87), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n202), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n225), .A2(KEYINPUT87), .A3(new_n244), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n229), .A2(new_n235), .B1(new_n237), .B2(new_n242), .ZN(new_n249));
  XOR2_X1   g048(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n250));
  AOI21_X1  g049(.A(KEYINPUT29), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n220), .A2(new_n222), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT88), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n243), .A3(new_n250), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(new_n221), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT88), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n247), .A2(new_n248), .A3(new_n253), .A4(new_n257), .ZN(new_n258));
  AOI211_X1 g057(.A(KEYINPUT86), .B(new_n218), .C1(new_n209), .C2(new_n210), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n219), .B1(new_n211), .B2(new_n260), .ZN(new_n261));
  OAI22_X1  g060(.A1(new_n259), .A2(new_n261), .B1(new_n260), .B2(new_n211), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n221), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n249), .B1(new_n263), .B2(new_n250), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n202), .B1(new_n264), .B2(new_n255), .ZN(new_n265));
  INV_X1    g064(.A(G22gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n258), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n258), .B2(new_n265), .ZN(new_n269));
  OAI21_X1  g068(.A(G78gat), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n258), .A2(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G22gat), .ZN(new_n272));
  INV_X1    g071(.A(G78gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n267), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT31), .B(G50gat), .ZN(new_n276));
  INV_X1    g075(.A(G106gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n276), .B(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n270), .A2(new_n274), .A3(new_n278), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n284));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(KEYINPUT23), .B2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n285), .A2(KEYINPUT23), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT24), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n292), .A2(new_n294), .B1(new_n290), .B2(new_n291), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n284), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n292), .A2(new_n294), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT66), .B(G190gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n297), .B1(new_n299), .B2(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(KEYINPUT23), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n287), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n300), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n296), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT28), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n298), .A2(new_n309), .A3(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT26), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n302), .A2(new_n315), .A3(new_n303), .ZN(new_n316));
  INV_X1    g115(.A(new_n286), .ZN(new_n317));
  INV_X1    g116(.A(new_n285), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n318), .B2(KEYINPUT26), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n316), .A2(new_n319), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(KEYINPUT67), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT67), .B1(new_n314), .B2(new_n320), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n308), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G113gat), .B(G120gat), .Z(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n330), .A2(new_n331), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n334), .B(new_n308), .C1(new_n322), .C2(new_n323), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n283), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT68), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT34), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n333), .A2(new_n335), .A3(new_n337), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G15gat), .B(G43gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n344), .B(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n337), .B1(new_n333), .B2(new_n335), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n346), .B1(new_n347), .B2(KEYINPUT33), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI221_X4 g150(.A(new_n349), .B1(KEYINPUT33), .B2(new_n346), .C1(new_n336), .C2(new_n338), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n343), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT33), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n357), .A3(new_n346), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n348), .A2(new_n350), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n339), .A2(new_n342), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n353), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT36), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n358), .A2(KEYINPUT69), .A3(new_n360), .A4(new_n359), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n353), .A2(new_n361), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n282), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n296), .A2(new_n307), .B1(new_n314), .B2(new_n320), .ZN(new_n370));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(KEYINPUT72), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n314), .A2(new_n320), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n376), .A2(new_n321), .B1(new_n296), .B2(new_n307), .ZN(new_n377));
  INV_X1    g176(.A(new_n372), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(new_n221), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n373), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT73), .B1(new_n380), .B2(new_n252), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n324), .A2(new_n221), .A3(new_n378), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n383));
  INV_X1    g182(.A(new_n252), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n373), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n378), .B1(new_n370), .B2(KEYINPUT29), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n252), .C1(new_n377), .C2(new_n378), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n324), .A2(new_n372), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(KEYINPUT74), .A3(new_n252), .A4(new_n387), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(new_n397), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n386), .A2(new_n393), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT30), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n393), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n398), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n386), .A2(new_n393), .A3(KEYINPUT30), .A4(new_n399), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n406), .A2(new_n407), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n405), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n249), .A2(KEYINPUT84), .A3(new_n334), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT84), .B1(new_n249), .B2(new_n334), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT4), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n330), .A2(KEYINPUT82), .A3(new_n331), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT82), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n332), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n415), .A2(new_n416), .A3(new_n418), .A4(new_n254), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n334), .A2(new_n236), .A3(new_n243), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n414), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n244), .A2(new_n416), .A3(new_n418), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n411), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n426), .B(KEYINPUT39), .C1(new_n425), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G1gat), .B(G29gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT0), .ZN(new_n433));
  XNOR2_X1  g232(.A(G57gat), .B(G85gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n433), .B(new_n434), .Z(new_n435));
  XOR2_X1   g234(.A(KEYINPUT89), .B(KEYINPUT39), .Z(new_n436));
  NAND3_X1  g235(.A1(new_n423), .A2(new_n425), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n431), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n431), .A2(KEYINPUT40), .A3(new_n435), .A4(new_n437), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT5), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n430), .B2(new_n425), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n421), .A3(new_n411), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n334), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n444), .A2(new_n419), .A3(new_n424), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n254), .A2(new_n416), .A3(new_n418), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n425), .B1(new_n448), .B2(new_n415), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n449), .A2(new_n414), .A3(new_n442), .A4(new_n422), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n435), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n440), .A2(new_n441), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n403), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n399), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT38), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(new_n403), .B2(KEYINPUT37), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n391), .A2(new_n384), .A3(new_n387), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n460), .B(KEYINPUT37), .C1(new_n384), .C2(new_n380), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n398), .B(new_n461), .C1(new_n403), .C2(KEYINPUT37), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n457), .A2(new_n459), .B1(new_n462), .B2(new_n458), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n435), .A3(new_n450), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT6), .B1(new_n466), .B2(new_n453), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n447), .A2(KEYINPUT85), .A3(new_n450), .A4(new_n435), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n468), .A2(new_n469), .B1(new_n451), .B2(new_n452), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n400), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n410), .A2(new_n454), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n369), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n270), .A2(new_n274), .A3(new_n278), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n278), .B1(new_n270), .B2(new_n274), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n363), .A2(new_n365), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n409), .A2(new_n408), .ZN(new_n480));
  INV_X1    g279(.A(new_n405), .ZN(new_n481));
  INV_X1    g280(.A(new_n467), .ZN(new_n482));
  INV_X1    g281(.A(new_n470), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n474), .B1(new_n479), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n366), .A2(new_n368), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n353), .A2(new_n361), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n475), .A2(new_n476), .A3(new_n487), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n486), .A2(new_n282), .B1(new_n488), .B2(KEYINPUT35), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n473), .B(new_n485), .C1(new_n489), .C2(new_n484), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n491));
  INV_X1    g290(.A(G50gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(G43gat), .ZN(new_n493));
  INV_X1    g292(.A(G43gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G50gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OR3_X1    g297(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(KEYINPUT90), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n506), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n499), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n508), .A2(new_n503), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n491), .B(new_n504), .C1(new_n509), .C2(new_n502), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n500), .ZN(new_n512));
  NOR3_X1   g311(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n513));
  OAI22_X1  g312(.A1(new_n511), .A2(KEYINPUT15), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n502), .A2(new_n503), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n502), .B1(new_n508), .B2(new_n503), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT91), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(G1gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT16), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(G1gat), .B2(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G8gat), .ZN(new_n524));
  INV_X1    g323(.A(G8gat), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n522), .B(new_n525), .C1(G1gat), .C2(new_n519), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n518), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n510), .A2(new_n518), .A3(KEYINPUT93), .A4(new_n527), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT92), .B(KEYINPUT17), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n510), .A2(new_n518), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n527), .ZN(new_n537));
  OAI211_X1 g336(.A(KEYINPUT17), .B(new_n504), .C1(new_n509), .C2(new_n502), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n532), .A2(new_n533), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT18), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n540), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n510), .A2(new_n518), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n532), .B1(new_n546), .B2(new_n527), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n533), .B(KEYINPUT13), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n543), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT12), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n543), .A2(new_n555), .A3(new_n545), .A4(new_n549), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(G64gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n562), .B(new_n564), .C1(G57gat), .C2(new_n563), .ZN(new_n565));
  INV_X1    g364(.A(G71gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n273), .A3(KEYINPUT9), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n567), .B1(new_n566), .B2(new_n273), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n561), .A2(G64gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n563), .A2(G57gat), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT9), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G71gat), .B(G78gat), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT96), .ZN(new_n578));
  XOR2_X1   g377(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G183gat), .B(G211gat), .Z(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT98), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n580), .B(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n568), .A2(new_n565), .B1(new_n572), .B2(new_n573), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n527), .B1(KEYINPUT21), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT97), .ZN(new_n586));
  XNOR2_X1  g385(.A(G127gat), .B(G155gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n586), .B(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT8), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT100), .ZN(new_n599));
  OR2_X1    g398(.A1(G85gat), .A2(G92gat), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G99gat), .B(G106gat), .ZN(new_n602));
  AND2_X1   g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n603), .A2(new_n604), .A3(new_n605), .A4(KEYINPUT7), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT7), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n598), .B2(KEYINPUT101), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n601), .A2(new_n602), .A3(new_n606), .A4(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n602), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n605), .A2(G85gat), .A3(G92gat), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n604), .A2(KEYINPUT7), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n599), .A3(new_n600), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n595), .B1(new_n546), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n536), .A2(new_n538), .A3(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n620), .B(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT99), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n623), .A2(new_n627), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n632));
  NOR2_X1   g431(.A1(G85gat), .A2(G92gat), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(KEYINPUT100), .B2(new_n598), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n634), .A2(new_n606), .A3(new_n597), .A4(new_n608), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT102), .B1(new_n635), .B2(new_n610), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n616), .A2(new_n584), .A3(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n609), .B(new_n615), .C1(new_n575), .C2(KEYINPUT102), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  NOR3_X1   g439(.A1(new_n616), .A2(new_n640), .A3(new_n575), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n631), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n637), .A2(new_n638), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n642), .B(new_n645), .C1(new_n631), .C2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n631), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n650), .B(new_n631), .C1(new_n639), .C2(new_n641), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n648), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n647), .B1(new_n652), .B2(new_n645), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT105), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655));
  OAI211_X1 g454(.A(new_n655), .B(new_n647), .C1(new_n652), .C2(new_n645), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n594), .A2(new_n630), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n490), .A2(new_n559), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n482), .A2(new_n483), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(new_n520), .ZN(G1324gat));
  NOR2_X1   g462(.A1(new_n659), .A2(new_n410), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(KEYINPUT42), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(G8gat), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n665), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n667), .B2(new_n668), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n666), .B(new_n669), .C1(new_n671), .C2(KEYINPUT42), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n659), .B2(new_n486), .ZN(new_n673));
  INV_X1    g472(.A(new_n478), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n659), .B2(new_n675), .ZN(G1326gat));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n477), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT43), .B(G22gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(new_n630), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(new_n657), .A3(new_n593), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n490), .A2(new_n559), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(G29gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n660), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT107), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n473), .A2(new_n485), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n486), .A2(new_n282), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n484), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n630), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n688), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n490), .A2(KEYINPUT108), .A3(KEYINPUT44), .A4(new_n630), .ZN(new_n696));
  INV_X1    g495(.A(new_n559), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(new_n593), .A3(new_n657), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G29gat), .B1(new_n699), .B2(new_n661), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n686), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n687), .A2(new_n700), .A3(new_n701), .ZN(G1328gat));
  INV_X1    g501(.A(G36gat), .ZN(new_n703));
  INV_X1    g502(.A(new_n410), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n682), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT109), .B(KEYINPUT46), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(G36gat), .B1(new_n699), .B2(new_n410), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1329gat));
  NOR2_X1   g508(.A1(new_n674), .A2(G43gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n682), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G43gat), .B1(new_n699), .B2(new_n486), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1330gat));
  INV_X1    g516(.A(KEYINPUT111), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n682), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n282), .A2(new_n492), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n682), .B2(new_n718), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n719), .A2(new_n721), .B1(KEYINPUT112), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G50gat), .B1(new_n699), .B2(new_n477), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n722), .A2(KEYINPUT112), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1331gat));
  INV_X1    g526(.A(new_n490), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n697), .A2(new_n593), .A3(new_n680), .A4(new_n657), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n660), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g531(.A1(new_n728), .A2(new_n410), .A3(new_n729), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  AND2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n734), .ZN(G1333gat));
  INV_X1    g536(.A(new_n486), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n566), .B1(new_n730), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n674), .A2(G71gat), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n730), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g541(.A1(new_n730), .A2(new_n282), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G78gat), .ZN(G1335gat));
  INV_X1    g543(.A(new_n657), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n593), .A3(new_n559), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n695), .A2(new_n696), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(G85gat), .B1(new_n747), .B2(new_n661), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n749), .B(new_n630), .C1(new_n689), .C2(new_n692), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n593), .A2(new_n559), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n749), .B1(new_n490), .B2(new_n630), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT51), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n693), .A2(KEYINPUT113), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(new_n756), .A3(new_n751), .A4(new_n750), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n661), .A2(G85gat), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n754), .A2(new_n757), .A3(new_n657), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n748), .A2(new_n759), .ZN(G1336gat));
  OAI21_X1  g559(.A(G92gat), .B1(new_n747), .B2(new_n410), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n410), .A2(new_n745), .A3(G92gat), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n752), .B2(new_n753), .ZN(new_n765));
  INV_X1    g564(.A(new_n764), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n755), .A2(new_n751), .A3(new_n750), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n763), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n761), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI211_X1 g569(.A(KEYINPUT115), .B(new_n763), .C1(new_n765), .C2(new_n767), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT52), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n754), .A2(new_n757), .A3(new_n762), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n761), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n747), .B2(new_n486), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n674), .A2(new_n745), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(G99gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n754), .A2(new_n757), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n777), .A2(new_n781), .ZN(G1338gat));
  NAND4_X1  g581(.A1(new_n695), .A2(new_n282), .A3(new_n696), .A4(new_n746), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(G106gat), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n477), .A2(G106gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n657), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n765), .B2(new_n767), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT53), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n754), .A2(new_n757), .A3(new_n657), .A4(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT53), .B1(new_n783), .B2(G106gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n789), .A2(new_n790), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n658), .A2(new_n697), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n547), .A2(new_n548), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n533), .B1(new_n532), .B2(new_n539), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n554), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n654), .A2(new_n558), .A3(new_n656), .A4(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n649), .A2(new_n802), .A3(new_n651), .ZN(new_n803));
  INV_X1    g602(.A(new_n645), .ZN(new_n804));
  OR3_X1    g603(.A1(new_n639), .A2(new_n631), .A3(new_n641), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n805), .A2(KEYINPUT54), .A3(new_n642), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n803), .A2(new_n806), .A3(KEYINPUT55), .A4(new_n804), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n647), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n801), .B1(new_n697), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n680), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n558), .A2(new_n800), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n680), .A2(new_n814), .A3(new_n811), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n797), .B1(new_n594), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n282), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n704), .A2(new_n661), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n478), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(G113gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n697), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n818), .A2(new_n661), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n488), .A3(new_n410), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n559), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n823), .B1(new_n822), .B2(new_n827), .ZN(G1340gat));
  OR3_X1    g627(.A1(new_n825), .A2(G120gat), .A3(new_n745), .ZN(new_n829));
  OAI21_X1  g628(.A(G120gat), .B1(new_n821), .B2(new_n745), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n829), .B1(new_n832), .B2(new_n833), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n821), .B2(new_n594), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n594), .A2(G127gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT118), .Z(G1342gat));
  OR3_X1    g637(.A1(new_n825), .A2(G134gat), .A3(new_n680), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  OAI21_X1  g639(.A(G134gat), .B1(new_n821), .B2(new_n680), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(G1343gat));
  INV_X1    g642(.A(new_n820), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n738), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n477), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n807), .A2(new_n808), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n810), .A2(new_n647), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n809), .A2(KEYINPUT119), .A3(new_n647), .A4(new_n810), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n559), .A3(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n856), .A3(new_n801), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n680), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n856), .B1(new_n855), .B2(new_n801), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n849), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n801), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT120), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(KEYINPUT121), .A3(new_n680), .A4(new_n857), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(new_n816), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n594), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n848), .B1(new_n865), .B2(new_n796), .ZN(new_n866));
  INV_X1    g665(.A(new_n818), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT57), .B1(new_n867), .B2(new_n282), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n559), .B(new_n845), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G141gat), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873));
  AOI211_X1 g672(.A(new_n690), .B(new_n704), .C1(new_n824), .C2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT122), .B1(new_n818), .B2(new_n661), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n697), .A2(G141gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n872), .A2(new_n878), .A3(KEYINPUT58), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT58), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n870), .B(new_n877), .C1(new_n871), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n881), .ZN(G1344gat));
  NOR3_X1   g681(.A1(new_n844), .A2(new_n738), .A3(new_n745), .ZN(new_n883));
  AND4_X1   g682(.A1(new_n558), .A2(new_n654), .A3(new_n656), .A4(new_n800), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n811), .A2(new_n850), .B1(new_n557), .B2(new_n558), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n854), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n630), .B1(new_n886), .B2(new_n856), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n815), .B1(new_n887), .B2(new_n862), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n796), .B1(new_n888), .B2(new_n593), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n889), .B2(new_n282), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n818), .A2(new_n848), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT125), .B(new_n883), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G148gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n816), .B1(new_n858), .B2(new_n859), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n797), .B1(new_n894), .B2(new_n594), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n846), .B1(new_n895), .B2(new_n477), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n896), .B1(new_n818), .B2(new_n848), .ZN(new_n897));
  AOI21_X1  g696(.A(KEYINPUT125), .B1(new_n897), .B2(new_n883), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT59), .B1(new_n893), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n657), .B(new_n845), .C1(new_n866), .C2(new_n868), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901));
  INV_X1    g700(.A(G148gat), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(KEYINPUT59), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n874), .A2(new_n875), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n902), .A3(new_n657), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n230), .A3(new_n593), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n866), .A2(new_n868), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n738), .A3(new_n844), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n912), .A2(new_n593), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n230), .ZN(G1346gat));
  AOI21_X1  g713(.A(G162gat), .B1(new_n907), .B2(new_n630), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n680), .A2(new_n231), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n912), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n818), .A2(new_n660), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n282), .A2(new_n410), .A3(new_n487), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n559), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n410), .A2(new_n660), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n819), .A2(new_n478), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(G169gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(new_n697), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n922), .A2(new_n926), .ZN(G1348gat));
  AOI21_X1  g726(.A(G176gat), .B1(new_n921), .B2(new_n657), .ZN(new_n928));
  AND4_X1   g727(.A1(G176gat), .A2(new_n819), .A3(new_n778), .A4(new_n923), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n924), .B2(new_n594), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n593), .A2(new_n309), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n931), .B(new_n933), .C1(new_n920), .C2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n936));
  XOR2_X1   g735(.A(new_n935), .B(new_n936), .Z(G1350gat));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n298), .A3(new_n630), .ZN(new_n938));
  OAI21_X1  g737(.A(G190gat), .B1(new_n924), .B2(new_n680), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  NOR2_X1   g741(.A1(new_n690), .A2(new_n410), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n918), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n559), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n897), .A2(new_n486), .A3(new_n923), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n697), .A2(new_n213), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  NOR3_X1   g748(.A1(new_n944), .A2(G204gat), .A3(new_n745), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n947), .A2(new_n657), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n214), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n945), .A2(new_n203), .A3(new_n593), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n897), .A2(new_n486), .A3(new_n593), .A4(new_n923), .ZN(new_n956));
  AND4_X1   g755(.A1(new_n955), .A2(new_n956), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(G211gat), .B1(new_n955), .B2(KEYINPUT63), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n956), .A2(new_n959), .B1(new_n955), .B2(KEYINPUT63), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n954), .B1(new_n957), .B2(new_n960), .ZN(G1354gat));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n204), .A3(new_n630), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n947), .A2(new_n630), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n963), .B2(new_n204), .ZN(G1355gat));
endmodule


