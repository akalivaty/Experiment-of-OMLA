

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725;

  INV_X1 U368 ( .A(n542), .ZN(n519) );
  XNOR2_X1 U369 ( .A(n372), .B(n504), .ZN(n542) );
  AND2_X1 U370 ( .A1(n578), .A2(n577), .ZN(n364) );
  INV_X1 U371 ( .A(G953), .ZN(n713) );
  NAND2_X1 U372 ( .A1(n541), .A2(n519), .ZN(n532) );
  XNOR2_X2 U373 ( .A(n587), .B(n586), .ZN(n391) );
  NOR2_X2 U374 ( .A1(n723), .A2(n725), .ZN(n539) );
  NOR2_X2 U375 ( .A1(n589), .A2(n550), .ZN(n630) );
  NOR2_X1 U376 ( .A1(n639), .A2(n638), .ZN(n640) );
  AND2_X2 U377 ( .A1(n609), .A2(n608), .ZN(n693) );
  INV_X1 U378 ( .A(n532), .ZN(n624) );
  XNOR2_X1 U379 ( .A(G472), .B(n470), .ZN(n592) );
  AND2_X2 U380 ( .A1(n594), .A2(n364), .ZN(n579) );
  XNOR2_X1 U381 ( .A(n449), .B(G107), .ZN(n473) );
  XNOR2_X1 U382 ( .A(n460), .B(n398), .ZN(n475) );
  INV_X1 U383 ( .A(KEYINPUT78), .ZN(n418) );
  XNOR2_X1 U384 ( .A(n468), .B(n448), .ZN(n709) );
  XNOR2_X1 U385 ( .A(n475), .B(n395), .ZN(n703) );
  XNOR2_X1 U386 ( .A(n396), .B(n473), .ZN(n395) );
  XNOR2_X1 U387 ( .A(n474), .B(n397), .ZN(n396) );
  INV_X1 U388 ( .A(KEYINPUT73), .ZN(n397) );
  XOR2_X1 U389 ( .A(G137), .B(G140), .Z(n448) );
  XNOR2_X1 U390 ( .A(n485), .B(n419), .ZN(n501) );
  INV_X1 U391 ( .A(KEYINPUT10), .ZN(n419) );
  XNOR2_X1 U392 ( .A(n446), .B(n445), .ZN(n636) );
  NOR2_X1 U393 ( .A1(G902), .A2(n694), .ZN(n446) );
  OR2_X1 U394 ( .A1(n626), .A2(n624), .ZN(n528) );
  XNOR2_X1 U395 ( .A(G116), .B(G101), .ZN(n457) );
  XNOR2_X1 U396 ( .A(G119), .B(G113), .ZN(n461) );
  XOR2_X1 U397 ( .A(KEYINPUT23), .B(G128), .Z(n435) );
  XNOR2_X1 U398 ( .A(G119), .B(G110), .ZN(n434) );
  XNOR2_X1 U399 ( .A(G140), .B(G122), .ZN(n492) );
  XNOR2_X1 U400 ( .A(G110), .B(G104), .ZN(n449) );
  XOR2_X1 U401 ( .A(G146), .B(G101), .Z(n451) );
  NOR2_X1 U402 ( .A1(n521), .A2(n418), .ZN(n413) );
  OR2_X1 U403 ( .A1(n688), .A2(G902), .ZN(n372) );
  XNOR2_X1 U404 ( .A(n454), .B(G469), .ZN(n455) );
  NOR2_X1 U405 ( .A1(G902), .A2(n681), .ZN(n456) );
  XNOR2_X1 U406 ( .A(n515), .B(n387), .ZN(n468) );
  XNOR2_X1 U407 ( .A(n388), .B(G131), .ZN(n387) );
  INV_X1 U408 ( .A(KEYINPUT4), .ZN(n388) );
  XNOR2_X1 U409 ( .A(n484), .B(n367), .ZN(n486) );
  XNOR2_X1 U410 ( .A(n485), .B(n483), .ZN(n367) );
  AND2_X1 U411 ( .A1(n543), .A2(n652), .ZN(n491) );
  NAND2_X1 U412 ( .A1(n573), .A2(n345), .ZN(n375) );
  AND2_X1 U413 ( .A1(n377), .A2(KEYINPUT35), .ZN(n376) );
  INV_X1 U414 ( .A(n639), .ZN(n589) );
  XNOR2_X1 U415 ( .A(n441), .B(n440), .ZN(n694) );
  XNOR2_X1 U416 ( .A(n420), .B(n501), .ZN(n441) );
  AND2_X1 U417 ( .A1(n528), .A2(KEYINPUT74), .ZN(n526) );
  NOR2_X1 U418 ( .A1(G953), .A2(G237), .ZN(n494) );
  XNOR2_X1 U419 ( .A(n403), .B(KEYINPUT48), .ZN(n554) );
  XOR2_X1 U420 ( .A(KEYINPUT16), .B(G122), .Z(n474) );
  OR2_X1 U421 ( .A1(n600), .A2(n356), .ZN(n363) );
  XOR2_X1 U422 ( .A(G128), .B(G143), .Z(n482) );
  XNOR2_X1 U423 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n476) );
  INV_X1 U424 ( .A(KEYINPUT18), .ZN(n478) );
  OR2_X1 U425 ( .A1(G902), .A2(G237), .ZN(n487) );
  XNOR2_X1 U426 ( .A(n366), .B(KEYINPUT107), .ZN(n655) );
  AND2_X1 U427 ( .A1(n652), .A2(n651), .ZN(n366) );
  INV_X1 U428 ( .A(KEYINPUT35), .ZN(n381) );
  NAND2_X1 U429 ( .A1(n639), .A2(n638), .ZN(n593) );
  NOR2_X1 U430 ( .A1(n576), .A2(n636), .ZN(n638) );
  XNOR2_X1 U431 ( .A(n461), .B(n399), .ZN(n398) );
  INV_X1 U432 ( .A(KEYINPUT3), .ZN(n399) );
  XOR2_X1 U433 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n463) );
  XNOR2_X1 U434 ( .A(G137), .B(G146), .ZN(n464) );
  XOR2_X1 U435 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n465) );
  NAND2_X1 U436 ( .A1(n359), .A2(n357), .ZN(n712) );
  NOR2_X1 U437 ( .A1(n633), .A2(n358), .ZN(n357) );
  INV_X1 U438 ( .A(n554), .ZN(n359) );
  INV_X1 U439 ( .A(n634), .ZN(n358) );
  INV_X1 U440 ( .A(n501), .ZN(n710) );
  XNOR2_X1 U441 ( .A(n436), .B(n433), .ZN(n420) );
  XNOR2_X1 U442 ( .A(n482), .B(n447), .ZN(n515) );
  INV_X1 U443 ( .A(G134), .ZN(n447) );
  XNOR2_X1 U444 ( .A(G116), .B(G107), .ZN(n505) );
  XOR2_X1 U445 ( .A(KEYINPUT101), .B(G122), .Z(n506) );
  XNOR2_X1 U446 ( .A(KEYINPUT7), .B(KEYINPUT102), .ZN(n507) );
  XOR2_X1 U447 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n508) );
  XNOR2_X1 U448 ( .A(n500), .B(n373), .ZN(n688) );
  XNOR2_X1 U449 ( .A(n501), .B(n346), .ZN(n373) );
  XNOR2_X1 U450 ( .A(G113), .B(G104), .ZN(n498) );
  XNOR2_X1 U451 ( .A(n473), .B(n452), .ZN(n453) );
  NAND2_X1 U452 ( .A1(n411), .A2(n410), .ZN(n543) );
  NAND2_X1 U453 ( .A1(n693), .A2(G475), .ZN(n370) );
  XNOR2_X1 U454 ( .A(n676), .B(n675), .ZN(n677) );
  NOR2_X1 U455 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U456 ( .A1(n383), .A2(n382), .ZN(n720) );
  AND2_X1 U457 ( .A1(n380), .A2(n379), .ZN(n383) );
  NAND2_X1 U458 ( .A1(n376), .A2(n375), .ZN(n382) );
  NAND2_X1 U459 ( .A1(n588), .A2(n582), .ZN(n583) );
  OR2_X1 U460 ( .A1(n639), .A2(n401), .ZN(n400) );
  NAND2_X1 U461 ( .A1(n402), .A2(n636), .ZN(n401) );
  INV_X1 U462 ( .A(n645), .ZN(n402) );
  AND2_X1 U463 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U464 ( .A1(n393), .A2(n368), .ZN(n392) );
  XNOR2_X1 U465 ( .A(n394), .B(n354), .ZN(n393) );
  NAND2_X1 U466 ( .A1(n407), .A2(n368), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n407) );
  INV_X1 U468 ( .A(n694), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n362), .B(n361), .ZN(G60) );
  INV_X1 U470 ( .A(KEYINPUT60), .ZN(n361) );
  NAND2_X1 U471 ( .A1(n369), .A2(n368), .ZN(n362) );
  XNOR2_X1 U472 ( .A(n370), .B(n355), .ZN(n369) );
  XNOR2_X1 U473 ( .A(n384), .B(KEYINPUT118), .ZN(n672) );
  AND2_X1 U474 ( .A1(n575), .A2(n572), .ZN(n345) );
  XOR2_X1 U475 ( .A(n493), .B(n492), .Z(n346) );
  XNOR2_X1 U476 ( .A(KEYINPUT117), .B(n671), .ZN(n347) );
  NOR2_X1 U477 ( .A1(n611), .A2(n363), .ZN(n348) );
  AND2_X1 U478 ( .A1(n575), .A2(KEYINPUT34), .ZN(n349) );
  AND2_X1 U479 ( .A1(n531), .A2(n530), .ZN(n350) );
  NOR2_X1 U480 ( .A1(n581), .A2(n400), .ZN(n351) );
  AND2_X1 U481 ( .A1(n345), .A2(n381), .ZN(n352) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT72), .Z(n353) );
  XOR2_X1 U483 ( .A(n610), .B(KEYINPUT62), .Z(n354) );
  XNOR2_X1 U484 ( .A(n709), .B(n453), .ZN(n681) );
  XOR2_X1 U485 ( .A(n688), .B(n687), .Z(n355) );
  AND2_X1 U486 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n356) );
  NOR2_X1 U487 ( .A1(G952), .A2(n713), .ZN(n695) );
  INV_X1 U488 ( .A(n695), .ZN(n368) );
  NAND2_X1 U489 ( .A1(n585), .A2(n421), .ZN(n587) );
  AND2_X2 U490 ( .A1(n584), .A2(n721), .ZN(n421) );
  NOR2_X2 U491 ( .A1(n581), .A2(n580), .ZN(n588) );
  NAND2_X1 U492 ( .A1(n624), .A2(n546), .ZN(n555) );
  XNOR2_X2 U493 ( .A(n360), .B(KEYINPUT86), .ZN(n548) );
  NAND2_X1 U494 ( .A1(n540), .A2(n651), .ZN(n360) );
  XNOR2_X1 U495 ( .A(n365), .B(n680), .ZN(G51) );
  NOR2_X2 U496 ( .A1(n679), .A2(n695), .ZN(n365) );
  INV_X1 U497 ( .A(n528), .ZN(n656) );
  XNOR2_X1 U498 ( .A(n517), .B(n371), .ZN(n626) );
  INV_X1 U499 ( .A(KEYINPUT103), .ZN(n371) );
  NAND2_X1 U500 ( .A1(n374), .A2(n638), .ZN(n597) );
  NAND2_X1 U501 ( .A1(n525), .A2(n374), .ZN(n536) );
  XNOR2_X2 U502 ( .A(n374), .B(KEYINPUT1), .ZN(n639) );
  XNOR2_X2 U503 ( .A(n456), .B(n455), .ZN(n374) );
  NAND2_X1 U504 ( .A1(n574), .A2(n349), .ZN(n377) );
  NAND2_X1 U505 ( .A1(n574), .A2(n378), .ZN(n380) );
  AND2_X1 U506 ( .A1(n349), .A2(n381), .ZN(n378) );
  NAND2_X1 U507 ( .A1(n573), .A2(n352), .ZN(n379) );
  NAND2_X1 U508 ( .A1(n386), .A2(n385), .ZN(n384) );
  XNOR2_X1 U509 ( .A(n667), .B(KEYINPUT2), .ZN(n385) );
  AND2_X1 U510 ( .A1(n668), .A2(n347), .ZN(n386) );
  XNOR2_X2 U511 ( .A(n389), .B(KEYINPUT0), .ZN(n594) );
  NOR2_X2 U512 ( .A1(n565), .A2(n564), .ZN(n389) );
  XNOR2_X2 U513 ( .A(n548), .B(n520), .ZN(n565) );
  NOR2_X4 U514 ( .A1(n696), .A2(n712), .ZN(n667) );
  XNOR2_X2 U515 ( .A(n390), .B(n601), .ZN(n696) );
  NAND2_X1 U516 ( .A1(n348), .A2(n391), .ZN(n390) );
  XNOR2_X1 U517 ( .A(n392), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U518 ( .A1(n693), .A2(G472), .ZN(n394) );
  XNOR2_X2 U519 ( .A(n579), .B(n353), .ZN(n581) );
  NAND2_X1 U520 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U521 ( .A(n539), .B(n538), .ZN(n404) );
  AND2_X1 U522 ( .A1(n553), .A2(n350), .ZN(n405) );
  XNOR2_X1 U523 ( .A(n406), .B(KEYINPUT121), .ZN(G66) );
  NAND2_X1 U524 ( .A1(n693), .A2(G217), .ZN(n409) );
  NAND2_X1 U525 ( .A1(n415), .A2(n472), .ZN(n410) );
  NAND2_X1 U526 ( .A1(n412), .A2(n472), .ZN(n411) );
  AND2_X1 U527 ( .A1(n414), .A2(n413), .ZN(n412) );
  INV_X1 U528 ( .A(n597), .ZN(n414) );
  NAND2_X1 U529 ( .A1(n417), .A2(n416), .ZN(n415) );
  NAND2_X1 U530 ( .A1(n521), .A2(n418), .ZN(n416) );
  NAND2_X1 U531 ( .A1(n597), .A2(n418), .ZN(n417) );
  XNOR2_X1 U532 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U533 ( .A1(n602), .A2(n674), .ZN(n489) );
  XNOR2_X1 U534 ( .A(n467), .B(n466), .ZN(n422) );
  XNOR2_X1 U535 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n538) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n481), .B(n480), .ZN(n484) );
  INV_X1 U538 ( .A(KEYINPUT91), .ZN(n432) );
  XNOR2_X1 U539 ( .A(n569), .B(KEYINPUT70), .ZN(n570) );
  XNOR2_X1 U540 ( .A(n432), .B(KEYINPUT24), .ZN(n433) );
  XNOR2_X1 U541 ( .A(n475), .B(n422), .ZN(n469) );
  XNOR2_X1 U542 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U543 ( .A1(n607), .A2(n606), .ZN(n609) );
  XNOR2_X1 U544 ( .A(G902), .B(KEYINPUT15), .ZN(n603) );
  INV_X1 U545 ( .A(n603), .ZN(n602) );
  NAND2_X1 U546 ( .A1(G237), .A2(G234), .ZN(n423) );
  XNOR2_X1 U547 ( .A(n423), .B(KEYINPUT14), .ZN(n424) );
  NAND2_X1 U548 ( .A1(G952), .A2(n424), .ZN(n665) );
  NOR2_X1 U549 ( .A1(G953), .A2(n665), .ZN(n563) );
  NAND2_X1 U550 ( .A1(G902), .A2(n424), .ZN(n425) );
  XNOR2_X1 U551 ( .A(KEYINPUT89), .B(n425), .ZN(n426) );
  NAND2_X1 U552 ( .A1(n426), .A2(G953), .ZN(n560) );
  NOR2_X1 U553 ( .A1(G900), .A2(n560), .ZN(n427) );
  XOR2_X1 U554 ( .A(KEYINPUT105), .B(n427), .Z(n428) );
  NOR2_X1 U555 ( .A1(n563), .A2(n428), .ZN(n521) );
  XOR2_X1 U556 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n430) );
  NAND2_X1 U557 ( .A1(G234), .A2(n603), .ZN(n429) );
  XNOR2_X1 U558 ( .A(n430), .B(n429), .ZN(n442) );
  NAND2_X1 U559 ( .A1(n442), .A2(G221), .ZN(n431) );
  XNOR2_X1 U560 ( .A(KEYINPUT21), .B(n431), .ZN(n635) );
  XOR2_X1 U561 ( .A(KEYINPUT95), .B(n635), .Z(n576) );
  XOR2_X1 U562 ( .A(G125), .B(G146), .Z(n485) );
  XNOR2_X1 U563 ( .A(n435), .B(n434), .ZN(n436) );
  NAND2_X1 U564 ( .A1(G234), .A2(n713), .ZN(n437) );
  XOR2_X1 U565 ( .A(KEYINPUT8), .B(n437), .Z(n511) );
  NAND2_X1 U566 ( .A1(n511), .A2(G221), .ZN(n439) );
  XNOR2_X1 U567 ( .A(n448), .B(KEYINPUT92), .ZN(n438) );
  XOR2_X1 U568 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n444) );
  NAND2_X1 U569 ( .A1(n442), .A2(G217), .ZN(n443) );
  XNOR2_X1 U570 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U571 ( .A1(G227), .A2(n713), .ZN(n450) );
  XNOR2_X1 U572 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U573 ( .A(KEYINPUT67), .B(KEYINPUT68), .ZN(n454) );
  INV_X1 U574 ( .A(n457), .ZN(n459) );
  XNOR2_X1 U575 ( .A(KEYINPUT87), .B(KEYINPUT69), .ZN(n458) );
  XNOR2_X1 U576 ( .A(n459), .B(n458), .ZN(n460) );
  NAND2_X1 U577 ( .A1(n494), .A2(G210), .ZN(n462) );
  XNOR2_X1 U578 ( .A(n463), .B(n462), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U580 ( .A(n469), .B(n468), .ZN(n610) );
  NOR2_X1 U581 ( .A1(G902), .A2(n610), .ZN(n470) );
  INV_X1 U582 ( .A(n592), .ZN(n645) );
  NAND2_X1 U583 ( .A1(G214), .A2(n487), .ZN(n651) );
  NAND2_X1 U584 ( .A1(n645), .A2(n651), .ZN(n471) );
  XOR2_X1 U585 ( .A(KEYINPUT30), .B(n471), .Z(n472) );
  XNOR2_X1 U586 ( .A(KEYINPUT38), .B(KEYINPUT75), .ZN(n490) );
  XOR2_X1 U587 ( .A(KEYINPUT80), .B(KEYINPUT88), .Z(n477) );
  XNOR2_X1 U588 ( .A(n477), .B(n476), .ZN(n481) );
  NAND2_X1 U589 ( .A1(G224), .A2(n713), .ZN(n479) );
  INV_X1 U590 ( .A(n482), .ZN(n483) );
  XNOR2_X1 U591 ( .A(n703), .B(n486), .ZN(n674) );
  NAND2_X1 U592 ( .A1(G210), .A2(n487), .ZN(n488) );
  XNOR2_X2 U593 ( .A(n489), .B(n488), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n490), .B(n540), .ZN(n652) );
  XNOR2_X1 U595 ( .A(n491), .B(KEYINPUT39), .ZN(n533) );
  XOR2_X1 U596 ( .A(KEYINPUT97), .B(G143), .Z(n493) );
  XOR2_X1 U597 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n496) );
  NAND2_X1 U598 ( .A1(n494), .A2(G214), .ZN(n495) );
  XNOR2_X1 U599 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U600 ( .A(n497), .B(G131), .Z(n499) );
  XNOR2_X1 U601 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U602 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n503) );
  XNOR2_X1 U603 ( .A(KEYINPUT98), .B(G475), .ZN(n502) );
  XNOR2_X1 U604 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U605 ( .A(n506), .B(n505), .ZN(n510) );
  XNOR2_X1 U606 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U607 ( .A(n510), .B(n509), .Z(n513) );
  NAND2_X1 U608 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U609 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U610 ( .A(n515), .B(n514), .ZN(n689) );
  NOR2_X1 U611 ( .A1(n689), .A2(G902), .ZN(n516) );
  XNOR2_X1 U612 ( .A(n516), .B(G478), .ZN(n541) );
  NOR2_X1 U613 ( .A1(n519), .A2(n541), .ZN(n517) );
  INV_X1 U614 ( .A(n626), .ZN(n518) );
  NOR2_X1 U615 ( .A1(n533), .A2(n518), .ZN(n633) );
  XNOR2_X1 U616 ( .A(KEYINPUT79), .B(KEYINPUT19), .ZN(n520) );
  NOR2_X1 U617 ( .A1(n635), .A2(n521), .ZN(n522) );
  NAND2_X1 U618 ( .A1(n522), .A2(n636), .ZN(n545) );
  NOR2_X1 U619 ( .A1(n592), .A2(n545), .ZN(n524) );
  XNOR2_X1 U620 ( .A(KEYINPUT106), .B(KEYINPUT28), .ZN(n523) );
  XNOR2_X1 U621 ( .A(n524), .B(n523), .ZN(n525) );
  NOR2_X1 U622 ( .A1(n565), .A2(n536), .ZN(n622) );
  NAND2_X1 U623 ( .A1(n526), .A2(n622), .ZN(n527) );
  XOR2_X1 U624 ( .A(n527), .B(KEYINPUT47), .Z(n531) );
  NOR2_X1 U625 ( .A1(KEYINPUT74), .A2(n528), .ZN(n529) );
  NAND2_X1 U626 ( .A1(n529), .A2(n622), .ZN(n530) );
  NOR2_X1 U627 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U628 ( .A(n534), .B(KEYINPUT40), .ZN(n723) );
  NAND2_X1 U629 ( .A1(n542), .A2(n541), .ZN(n654) );
  NOR2_X1 U630 ( .A1(n654), .A2(n655), .ZN(n535) );
  XNOR2_X1 U631 ( .A(n535), .B(KEYINPUT41), .ZN(n670) );
  NOR2_X1 U632 ( .A1(n536), .A2(n670), .ZN(n537) );
  XNOR2_X1 U633 ( .A(n537), .B(KEYINPUT42), .ZN(n725) );
  INV_X1 U634 ( .A(n540), .ZN(n558) );
  NOR2_X1 U635 ( .A1(n542), .A2(n541), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n543), .A2(n575), .ZN(n544) );
  NOR2_X1 U637 ( .A1(n558), .A2(n544), .ZN(n621) );
  XOR2_X1 U638 ( .A(KEYINPUT81), .B(n621), .Z(n552) );
  XOR2_X1 U639 ( .A(n592), .B(KEYINPUT6), .Z(n567) );
  NOR2_X1 U640 ( .A1(n567), .A2(n545), .ZN(n546) );
  XNOR2_X1 U641 ( .A(KEYINPUT108), .B(n555), .ZN(n547) );
  XOR2_X1 U642 ( .A(KEYINPUT36), .B(n549), .Z(n550) );
  XNOR2_X1 U643 ( .A(KEYINPUT84), .B(n630), .ZN(n551) );
  NOR2_X1 U644 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U645 ( .A1(n639), .A2(n555), .ZN(n556) );
  NAND2_X1 U646 ( .A1(n556), .A2(n651), .ZN(n557) );
  XNOR2_X1 U647 ( .A(n557), .B(KEYINPUT43), .ZN(n559) );
  NAND2_X1 U648 ( .A1(n559), .A2(n558), .ZN(n634) );
  NOR2_X1 U649 ( .A1(G898), .A2(n560), .ZN(n561) );
  XNOR2_X1 U650 ( .A(n561), .B(KEYINPUT90), .ZN(n562) );
  NOR2_X1 U651 ( .A1(n563), .A2(n562), .ZN(n564) );
  INV_X1 U652 ( .A(n594), .ZN(n596) );
  INV_X1 U653 ( .A(KEYINPUT104), .ZN(n566) );
  XNOR2_X1 U654 ( .A(n593), .B(n566), .ZN(n568) );
  INV_X1 U655 ( .A(n567), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n568), .A2(n580), .ZN(n571) );
  INV_X1 U657 ( .A(KEYINPUT33), .ZN(n569) );
  XNOR2_X2 U658 ( .A(n571), .B(n570), .ZN(n669) );
  NOR2_X2 U659 ( .A1(n596), .A2(n669), .ZN(n574) );
  INV_X1 U660 ( .A(n574), .ZN(n573) );
  INV_X1 U661 ( .A(KEYINPUT34), .ZN(n572) );
  INV_X1 U662 ( .A(n720), .ZN(n585) );
  INV_X1 U663 ( .A(n576), .ZN(n577) );
  INV_X1 U664 ( .A(n654), .ZN(n578) );
  INV_X1 U665 ( .A(n351), .ZN(n584) );
  AND2_X1 U666 ( .A1(n639), .A2(n636), .ZN(n582) );
  XNOR2_X2 U667 ( .A(n583), .B(KEYINPUT32), .ZN(n721) );
  NOR2_X1 U668 ( .A1(KEYINPUT71), .A2(KEYINPUT44), .ZN(n586) );
  XNOR2_X1 U669 ( .A(n590), .B(KEYINPUT85), .ZN(n591) );
  NOR2_X1 U670 ( .A1(n636), .A2(n591), .ZN(n611) );
  NOR2_X1 U671 ( .A1(n593), .A2(n592), .ZN(n647) );
  NAND2_X1 U672 ( .A1(n647), .A2(n594), .ZN(n595) );
  XNOR2_X1 U673 ( .A(KEYINPUT31), .B(n595), .ZN(n627) );
  OR2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U675 ( .A1(n645), .A2(n598), .ZN(n614) );
  NOR2_X1 U676 ( .A1(n627), .A2(n614), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n656), .A2(n599), .ZN(n600) );
  XNOR2_X1 U678 ( .A(KEYINPUT45), .B(KEYINPUT65), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n667), .ZN(n607) );
  XOR2_X1 U680 ( .A(n603), .B(KEYINPUT82), .Z(n604) );
  NAND2_X1 U681 ( .A1(n604), .A2(KEYINPUT2), .ZN(n605) );
  XNOR2_X1 U682 ( .A(KEYINPUT66), .B(n605), .ZN(n606) );
  NAND2_X1 U683 ( .A1(KEYINPUT2), .A2(n667), .ZN(n608) );
  XOR2_X1 U684 ( .A(G101), .B(n611), .Z(G3) );
  XOR2_X1 U685 ( .A(G104), .B(KEYINPUT109), .Z(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n624), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n613), .B(n612), .ZN(G6) );
  XNOR2_X1 U688 ( .A(G107), .B(KEYINPUT110), .ZN(n618) );
  XOR2_X1 U689 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n616) );
  NAND2_X1 U690 ( .A1(n614), .A2(n626), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(G9) );
  XOR2_X1 U693 ( .A(G110), .B(n351), .Z(G12) );
  XOR2_X1 U694 ( .A(G128), .B(KEYINPUT29), .Z(n620) );
  NAND2_X1 U695 ( .A1(n622), .A2(n626), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n620), .B(n619), .ZN(G30) );
  XOR2_X1 U697 ( .A(G143), .B(n621), .Z(G45) );
  NAND2_X1 U698 ( .A1(n622), .A2(n624), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n623), .B(G146), .ZN(G48) );
  NAND2_X1 U700 ( .A1(n627), .A2(n624), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n625), .B(G113), .ZN(G15) );
  XOR2_X1 U702 ( .A(G116), .B(KEYINPUT111), .Z(n629) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U704 ( .A(n629), .B(n628), .ZN(G18) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT112), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT37), .ZN(n632) );
  XNOR2_X1 U707 ( .A(G125), .B(n632), .ZN(G27) );
  XOR2_X1 U708 ( .A(G134), .B(n633), .Z(G36) );
  XNOR2_X1 U709 ( .A(G140), .B(n634), .ZN(G42) );
  AND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U711 ( .A(KEYINPUT49), .B(n637), .ZN(n643) );
  XNOR2_X1 U712 ( .A(KEYINPUT50), .B(KEYINPUT113), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U717 ( .A(n648), .B(KEYINPUT51), .Z(n649) );
  XNOR2_X1 U718 ( .A(KEYINPUT114), .B(n649), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n670), .A2(n650), .ZN(n661) );
  NOR2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n658) );
  NOR2_X1 U722 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U724 ( .A1(n669), .A2(n659), .ZN(n660) );
  NOR2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U726 ( .A(n662), .B(KEYINPUT115), .Z(n663) );
  XNOR2_X1 U727 ( .A(KEYINPUT52), .B(n663), .ZN(n664) );
  NOR2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U729 ( .A(KEYINPUT116), .B(n666), .Z(n668) );
  NOR2_X1 U730 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U731 ( .A1(G953), .A2(n672), .ZN(n673) );
  XNOR2_X1 U732 ( .A(KEYINPUT53), .B(n673), .ZN(G75) );
  NAND2_X1 U733 ( .A1(n693), .A2(G210), .ZN(n678) );
  BUF_X1 U734 ( .A(n674), .Z(n676) );
  XOR2_X1 U735 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n675) );
  XOR2_X1 U736 ( .A(KEYINPUT83), .B(KEYINPUT56), .Z(n680) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n683) );
  XNOR2_X1 U738 ( .A(n681), .B(KEYINPUT119), .ZN(n682) );
  XNOR2_X1 U739 ( .A(n683), .B(n682), .ZN(n685) );
  NAND2_X1 U740 ( .A1(n693), .A2(G469), .ZN(n684) );
  XOR2_X1 U741 ( .A(n685), .B(n684), .Z(n686) );
  NOR2_X1 U742 ( .A1(n695), .A2(n686), .ZN(G54) );
  INV_X1 U743 ( .A(KEYINPUT59), .ZN(n687) );
  XNOR2_X1 U744 ( .A(n689), .B(KEYINPUT120), .ZN(n691) );
  NAND2_X1 U745 ( .A1(G478), .A2(n693), .ZN(n690) );
  XNOR2_X1 U746 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U747 ( .A1(n695), .A2(n692), .ZN(G63) );
  NOR2_X1 U748 ( .A1(G953), .A2(n696), .ZN(n702) );
  XOR2_X1 U749 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n698) );
  NAND2_X1 U750 ( .A1(G224), .A2(G953), .ZN(n697) );
  XNOR2_X1 U751 ( .A(n698), .B(n697), .ZN(n700) );
  INV_X1 U752 ( .A(G898), .ZN(n699) );
  NOR2_X1 U753 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(n708) );
  NOR2_X1 U755 ( .A1(G898), .A2(n713), .ZN(n705) );
  XOR2_X1 U756 ( .A(n703), .B(KEYINPUT124), .Z(n704) );
  NOR2_X1 U757 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U758 ( .A(KEYINPUT123), .B(n706), .Z(n707) );
  XOR2_X1 U759 ( .A(n708), .B(n707), .Z(G69) );
  XOR2_X1 U760 ( .A(n710), .B(n709), .Z(n711) );
  XNOR2_X1 U761 ( .A(n711), .B(KEYINPUT125), .ZN(n715) );
  XNOR2_X1 U762 ( .A(n712), .B(n715), .ZN(n714) );
  NAND2_X1 U763 ( .A1(n714), .A2(n713), .ZN(n719) );
  XNOR2_X1 U764 ( .A(G227), .B(n715), .ZN(n716) );
  NAND2_X1 U765 ( .A1(n716), .A2(G900), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n717), .A2(G953), .ZN(n718) );
  NAND2_X1 U767 ( .A1(n719), .A2(n718), .ZN(G72) );
  XOR2_X1 U768 ( .A(n720), .B(G122), .Z(G24) );
  XNOR2_X1 U769 ( .A(G119), .B(n721), .ZN(n722) );
  XNOR2_X1 U770 ( .A(n722), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U771 ( .A(G131), .B(KEYINPUT127), .ZN(n724) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(G33) );
  XOR2_X1 U773 ( .A(G137), .B(n725), .Z(G39) );
endmodule

