//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n567, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n479), .A2(new_n475), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(new_n475), .B2(G112), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n482), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n464), .A2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G102), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n479), .B2(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n492), .B1(new_n495), .B2(new_n475), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n475), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n479), .A2(KEYINPUT4), .A3(G138), .A4(new_n475), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n490), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n492), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n493), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n506), .A2(KEYINPUT66), .A3(new_n499), .A4(new_n500), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n502), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  OAI211_X1 g091(.A(new_n513), .B(new_n514), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(new_n512), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n516), .A2(new_n515), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT67), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(new_n520), .A3(G88), .ZN(new_n521));
  INV_X1    g096(.A(G75), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT68), .B1(new_n522), .B2(new_n509), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G75), .A3(G543), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n525), .C1(new_n518), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n519), .A2(new_n509), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(G651), .B1(new_n528), .B2(G50), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT69), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n521), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G166));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n528), .A2(G51), .B1(new_n513), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n517), .A2(new_n520), .A3(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(KEYINPUT70), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT70), .B1(new_n537), .B2(new_n539), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n528), .A2(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n517), .A2(new_n520), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  INV_X1    g124(.A(G77), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n518), .A2(new_n549), .B1(new_n550), .B2(new_n509), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI221_X1 g128(.A(KEYINPUT71), .B1(new_n550), .B2(new_n509), .C1(new_n518), .C2(new_n549), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(G651), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n548), .A2(new_n556), .ZN(G171));
  AND2_X1   g132(.A1(new_n517), .A2(new_n520), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G81), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n518), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n528), .B2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  AND3_X1   g141(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G36), .ZN(G176));
  XOR2_X1   g143(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n569));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n518), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  OAI211_X1 g151(.A(G53), .B(G543), .C1(new_n516), .C2(new_n515), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n577), .B(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G91), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n576), .B(new_n580), .C1(new_n546), .C2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G171), .ZN(G301));
  INV_X1    g158(.A(G166), .ZN(G303));
  OAI21_X1  g159(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n528), .A2(G49), .ZN(new_n586));
  INV_X1    g161(.A(G87), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n546), .C2(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n518), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n528), .B2(G48), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n546), .B2(new_n593), .ZN(G305));
  NAND3_X1  g169(.A1(new_n517), .A2(new_n520), .A3(G85), .ZN(new_n595));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n518), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n528), .B2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n595), .A2(new_n599), .A3(KEYINPUT74), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT75), .Z(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n558), .A2(new_n607), .A3(G92), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT76), .ZN(new_n610));
  XNOR2_X1  g185(.A(KEYINPUT77), .B(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n518), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(new_n528), .B2(G54), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT10), .B1(new_n546), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n608), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n606), .B1(G868), .B2(new_n617), .ZN(G284));
  OAI21_X1  g193(.A(new_n606), .B1(G868), .B2(new_n617), .ZN(G321));
  MUX2_X1   g194(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g195(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g196(.A(KEYINPUT78), .B(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n617), .B1(G860), .B2(new_n622), .ZN(G148));
  NAND2_X1  g198(.A1(new_n617), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n479), .A2(new_n491), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT79), .B(G2100), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G123), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n484), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n633), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2435), .ZN(new_n642));
  XOR2_X1   g217(.A(G2427), .B(G2438), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(KEYINPUT14), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n651), .B(new_n652), .Z(new_n653));
  AND2_X1   g228(.A1(new_n653), .A2(G14), .ZN(G401));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT83), .Z(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n656), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n659), .B2(new_n658), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT84), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n658), .A2(new_n659), .A3(new_n656), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  INV_X1    g240(.A(new_n656), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n658), .A3(new_n660), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2096), .Z(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(G2100), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT85), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  OAI221_X1 g259(.A(new_n679), .B1(new_n677), .B2(new_n675), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT87), .B(G1981), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT86), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n687), .B(new_n692), .ZN(G229));
  NAND3_X1  g268(.A1(new_n479), .A2(G128), .A3(G2105), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n479), .A2(G140), .A3(new_n475), .ZN(new_n695));
  OR2_X1    g270(.A1(G104), .A2(G2105), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n696), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT95), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT95), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(G26), .ZN(new_n706));
  OAI21_X1  g281(.A(KEYINPUT28), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(KEYINPUT28), .B2(new_n706), .ZN(new_n708));
  INV_X1    g283(.A(G2067), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G29), .A2(G33), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n491), .A2(G103), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n484), .A2(G139), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n714), .B(new_n715), .C1(new_n475), .C2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT97), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n711), .B1(new_n719), .B2(G29), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(G2072), .Z(new_n721));
  INV_X1    g296(.A(KEYINPUT93), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G4), .B2(G16), .ZN(new_n723));
  OR3_X1    g298(.A1(new_n722), .A2(G4), .A3(G16), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n723), .B(new_n724), .C1(new_n616), .C2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1348), .ZN(new_n727));
  NAND2_X1  g302(.A1(G299), .A2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT88), .B(G16), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT23), .ZN(new_n730));
  INV_X1    g305(.A(G20), .ZN(new_n731));
  OR3_X1    g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n729), .B2(new_n731), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1956), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n710), .A2(new_n721), .A3(new_n727), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n729), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n565), .B2(new_n729), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT94), .B(G1341), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n725), .A2(G5), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G171), .B2(new_n725), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n742), .B1(G1961), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n744), .A2(G1961), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n739), .A2(new_n741), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT24), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(G34), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(G34), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n477), .B2(G29), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT30), .B(G28), .Z(new_n763));
  MUX2_X1   g338(.A(new_n763), .B(new_n637), .S(G29), .Z(new_n764));
  NAND4_X1  g339(.A1(new_n753), .A2(new_n761), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n737), .A2(new_n752), .A3(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT90), .B(KEYINPUT34), .Z(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n725), .A2(G23), .ZN(new_n770));
  INV_X1    g345(.A(G288), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n725), .ZN(new_n772));
  AND2_X1   g347(.A1(new_n772), .A2(KEYINPUT91), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(KEYINPUT91), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT33), .B(G1976), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n776), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n773), .B2(new_n774), .ZN(new_n779));
  INV_X1    g354(.A(G1971), .ZN(new_n780));
  NAND2_X1  g355(.A1(G166), .A2(new_n729), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n729), .A2(G22), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n781), .A2(new_n780), .A3(new_n782), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n777), .B(new_n779), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n725), .A2(G6), .ZN(new_n786));
  INV_X1    g361(.A(G305), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(new_n725), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT32), .B(G1981), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n769), .B1(new_n785), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n784), .A2(new_n783), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n776), .B2(new_n775), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n794), .A2(new_n768), .A3(new_n779), .A4(new_n790), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(G290), .A2(new_n729), .ZN(new_n797));
  INV_X1    g372(.A(G24), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT89), .B1(new_n729), .B2(new_n798), .ZN(new_n799));
  OR3_X1    g374(.A1(new_n729), .A2(KEYINPUT89), .A3(new_n798), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1986), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n481), .A2(G119), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n484), .A2(G131), .ZN(new_n804));
  NOR2_X1   g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  OAI21_X1  g380(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  MUX2_X1   g382(.A(G25), .B(new_n807), .S(G29), .Z(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n808), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(KEYINPUT92), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n802), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n796), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT92), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(KEYINPUT36), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n767), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n819));
  INV_X1    g394(.A(G129), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n480), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n479), .A2(KEYINPUT98), .A3(G129), .A4(G2105), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n491), .A2(G105), .ZN(new_n824));
  INV_X1    g399(.A(G141), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n483), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT99), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n830), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT26), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n823), .A2(new_n827), .A3(new_n833), .ZN(new_n834));
  MUX2_X1   g409(.A(G32), .B(new_n834), .S(G29), .Z(new_n835));
  XOR2_X1   g410(.A(KEYINPUT27), .B(G1996), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(G16), .A2(G21), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G168), .B2(G16), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT100), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1966), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n814), .ZN(new_n844));
  AOI211_X1 g419(.A(new_n817), .B(new_n844), .C1(new_n792), .C2(new_n795), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n818), .A2(new_n838), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n704), .A2(G35), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G162), .B2(new_n704), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT29), .B(G2090), .Z(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n847), .A2(new_n851), .ZN(G311));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n847), .B2(new_n851), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n844), .B1(new_n792), .B2(new_n795), .ZN(new_n855));
  INV_X1    g430(.A(new_n817), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n766), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n857), .A2(new_n845), .A3(new_n842), .ZN(new_n858));
  INV_X1    g433(.A(new_n851), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n858), .A2(KEYINPUT101), .A3(new_n859), .A4(new_n838), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n854), .A2(new_n860), .ZN(G150));
  NAND2_X1  g436(.A1(G80), .A2(G543), .ZN(new_n862));
  INV_X1    g437(.A(G67), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n518), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(G651), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n528), .A2(G55), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n558), .B2(G93), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n565), .A2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n564), .A2(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n617), .A2(G559), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n871), .B1(new_n878), .B2(G860), .ZN(G145));
  NAND3_X1  g454(.A1(new_n834), .A2(new_n700), .A3(new_n701), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n826), .B1(new_n821), .B2(new_n822), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n702), .A2(new_n881), .A3(new_n833), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n496), .A2(new_n501), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n883), .B1(new_n880), .B2(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n719), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n882), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n506), .A2(new_n499), .A3(new_n500), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n880), .A2(new_n882), .A3(new_n883), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n717), .A3(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n629), .B(KEYINPUT103), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n886), .B2(new_n891), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n807), .B(KEYINPUT104), .ZN(new_n896));
  INV_X1    g471(.A(G142), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n483), .A2(KEYINPUT102), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT102), .B1(new_n483), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n481), .A2(G130), .ZN(new_n900));
  OR2_X1    g475(.A1(G106), .A2(G2105), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n901), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n896), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n894), .A2(new_n895), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n886), .A2(new_n891), .ZN(new_n907));
  INV_X1    g482(.A(new_n892), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n904), .B1(new_n909), .B2(new_n893), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT105), .B1(new_n906), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n907), .A2(KEYINPUT105), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n637), .B(new_n477), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n488), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n914), .B1(new_n906), .B2(new_n910), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n874), .B(new_n624), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n616), .A2(G299), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n616), .A2(G299), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(KEYINPUT41), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(new_n930), .A3(new_n924), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(new_n921), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n920), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT106), .B1(new_n922), .B2(new_n926), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(G290), .A2(new_n787), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n602), .A2(G305), .A3(new_n603), .ZN(new_n939));
  AOI21_X1  g514(.A(G166), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n938), .A2(G166), .A3(new_n939), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n941), .A2(new_n771), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n771), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT42), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n937), .A2(new_n946), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n868), .A2(G868), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(G295));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n949), .A2(new_n953), .A3(new_n951), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n949), .B2(new_n951), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(G331));
  NAND2_X1  g531(.A1(new_n558), .A2(G90), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(KEYINPUT109), .A3(new_n545), .A4(new_n555), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n548), .B2(new_n556), .ZN(new_n960));
  NAND3_X1  g535(.A1(G286), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n537), .A2(new_n539), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT70), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n540), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(KEYINPUT109), .A3(new_n536), .A4(G171), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n872), .A2(new_n873), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n874), .A2(new_n966), .A3(new_n961), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n874), .A2(new_n961), .A3(KEYINPUT110), .A4(new_n966), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n972), .A2(new_n932), .A3(new_n933), .A4(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n926), .A3(new_n971), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n945), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G37), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n945), .B1(new_n974), .B2(new_n975), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n925), .B1(new_n972), .B2(new_n973), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n971), .A2(new_n969), .B1(new_n928), .B2(new_n931), .ZN(new_n982));
  OAI22_X1  g557(.A1(new_n981), .A2(new_n982), .B1(new_n943), .B2(new_n944), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n976), .A3(new_n984), .A4(new_n977), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n984), .B1(new_n978), .B2(new_n979), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n976), .A3(new_n977), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n984), .B2(new_n988), .ZN(new_n989));
  MUX2_X1   g564(.A(new_n986), .B(new_n989), .S(KEYINPUT44), .Z(G397));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n502), .A2(new_n507), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n471), .A2(new_n476), .A3(G40), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n496), .B2(new_n501), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n996));
  AOI21_X1  g571(.A(G1956), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT119), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n999));
  NAND2_X1  g574(.A1(G299), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT120), .Z(new_n1001));
  NOR2_X1   g576(.A1(G299), .A2(new_n999), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT121), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n502), .A2(new_n507), .A3(new_n992), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(KEYINPUT114), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n994), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n998), .A2(new_n1004), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1009), .B1(new_n995), .B2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1348), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n995), .A2(new_n994), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1022), .A2(new_n1023), .B1(new_n709), .B2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1018), .A2(new_n616), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT114), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1016), .ZN(new_n1029));
  NOR4_X1   g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1012), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n993), .A2(new_n996), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT119), .B1(new_n1031), .B2(new_n735), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n1033), .B(G1956), .C1(new_n993), .C2(new_n996), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT122), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT122), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n998), .A2(new_n1037), .A3(new_n1017), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1004), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1026), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT61), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1004), .B1(new_n998), .B2(new_n1017), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1018), .B2(new_n1042), .ZN(new_n1043));
  NOR4_X1   g618(.A1(new_n1027), .A2(new_n1028), .A3(G1996), .A4(new_n1012), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT58), .B(G1341), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1024), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n565), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT59), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(new_n565), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1025), .B1(KEYINPUT60), .B2(new_n617), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n617), .A2(KEYINPUT60), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1043), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1039), .A2(new_n1041), .A3(new_n1018), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1040), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1027), .A2(new_n1028), .A3(new_n1012), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT53), .B1(new_n1060), .B2(new_n750), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1019), .B1(KEYINPUT50), .B2(new_n1005), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(G1961), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT45), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n995), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1009), .B(new_n1066), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(G171), .B(KEYINPUT54), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G286), .A2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1062), .A2(new_n760), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G8), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT51), .B(new_n1073), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1020), .A2(new_n1021), .A3(new_n760), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1078), .B(G8), .C1(new_n1081), .C2(G286), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1073), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT124), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1085), .B(new_n1073), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1077), .B(new_n1082), .C1(new_n1084), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1072), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1006), .B1(new_n888), .B2(new_n992), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1068), .B1(new_n1009), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n1011), .C1(new_n1090), .C2(new_n1009), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1064), .B(new_n1070), .C1(new_n1089), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(G303), .B2(G8), .ZN(new_n1095));
  NOR3_X1   g670(.A1(G166), .A2(KEYINPUT55), .A3(new_n1076), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT115), .B(G1971), .Z(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1022), .A2(G2090), .ZN(new_n1100));
  OAI211_X1 g675(.A(G8), .B(new_n1097), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1100), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1060), .B2(new_n1098), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1105), .A2(KEYINPUT116), .A3(G8), .A4(new_n1097), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1024), .A2(new_n1076), .ZN(new_n1108));
  INV_X1    g683(.A(G1976), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(G288), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n771), .A2(G1976), .ZN(new_n1111));
  OR3_X1    g686(.A1(new_n1110), .A2(KEYINPUT52), .A3(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(G305), .B(G1981), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n1114));
  OR2_X1    g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n1108), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1110), .A2(KEYINPUT52), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1112), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1031), .A2(G2090), .ZN(new_n1120));
  OAI21_X1  g695(.A(G8), .B1(new_n1099), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1097), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1093), .A2(new_n1107), .A3(new_n1119), .A4(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1088), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT123), .B(new_n1040), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1059), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1103), .A2(new_n1106), .A3(new_n1119), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1117), .A2(new_n1109), .A3(new_n771), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G305), .A2(G1981), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1130), .B(KEYINPUT117), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1108), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1128), .A2(KEYINPUT118), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT118), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1085), .B1(new_n1075), .B2(new_n1073), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1081), .A2(new_n1083), .A3(KEYINPUT124), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1082), .A4(new_n1077), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1107), .A2(new_n1119), .A3(new_n1139), .A4(new_n1123), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1087), .A2(KEYINPUT62), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(G171), .A3(new_n1069), .ZN(new_n1142));
  OAI22_X1  g717(.A1(new_n1133), .A2(new_n1134), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT63), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1105), .A2(G8), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n1122), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1107), .A2(new_n1146), .A3(new_n1119), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1075), .A2(new_n1076), .A3(G286), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1107), .A2(new_n1119), .A3(new_n1123), .A4(new_n1148), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1147), .A2(new_n1148), .B1(new_n1149), .B2(new_n1144), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1143), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1127), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n702), .B(new_n709), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1089), .A2(new_n1009), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n1155), .B(KEYINPUT113), .Z(new_n1156));
  INV_X1    g731(.A(new_n1154), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n834), .B(G1996), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n807), .B(new_n810), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1154), .A2(G290), .A3(G1986), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1157), .A2(G1986), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1162), .B1(new_n1163), .B2(G290), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT112), .Z(new_n1165));
  NOR2_X1   g740(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1152), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1154), .A2(G1996), .ZN(new_n1169));
  NAND2_X1  g744(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1169), .B(new_n1170), .Z(new_n1171));
  NAND3_X1  g746(.A1(new_n1153), .A2(new_n881), .A3(new_n833), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1168), .B(new_n1171), .C1(new_n1157), .C2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n807), .A2(new_n809), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1159), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n703), .A2(new_n709), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1154), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1162), .B(KEYINPUT48), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1161), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1174), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1167), .A2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g757(.A(new_n461), .B1(new_n916), .B2(new_n917), .ZN(new_n1184));
  NOR2_X1   g758(.A1(G401), .A2(G229), .ZN(new_n1185));
  NAND4_X1  g759(.A1(new_n986), .A2(new_n1184), .A3(new_n670), .A4(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g760(.A(new_n1186), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1188));
  XNOR2_X1  g762(.A(new_n1186), .B(new_n1188), .ZN(G225));
endmodule


