//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1233, new_n1234, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G107), .ZN(new_n220));
  INV_X1    g0020(.A(G264), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n211), .B1(new_n215), .B2(new_n216), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n218), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT67), .B(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G97), .B(G107), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  AND2_X1   g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(new_n212), .ZN(new_n250));
  INV_X1    g0050(.A(G274), .ZN(new_n251));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n257), .A2(G223), .B1(G77), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n255), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  AND3_X1   g0069(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(KEYINPUT70), .B1(new_n268), .B2(new_n269), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n254), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n253), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n268), .A2(new_n269), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n252), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT69), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n275), .A2(new_n280), .A3(new_n276), .A4(new_n277), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n273), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G200), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  INV_X1    g0086(.A(G190), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n284), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n286), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n212), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n204), .A2(new_n213), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n213), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n295), .A2(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n293), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G13), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n302), .A2(new_n213), .A3(G1), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n293), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n303), .A2(new_n293), .A3(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n252), .A2(G20), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n307), .A2(new_n308), .A3(G50), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n303), .A2(new_n202), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n301), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT9), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n289), .A2(new_n290), .A3(new_n291), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n291), .A2(new_n313), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT10), .B1(new_n315), .B2(new_n288), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n284), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n273), .A2(new_n321), .A3(new_n283), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G68), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n303), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n298), .A2(G50), .B1(G20), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n205), .B2(new_n296), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n303), .A2(new_n293), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G68), .A3(new_n309), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n327), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(KEYINPUT11), .B1(new_n329), .B2(new_n293), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n255), .A2(G226), .A3(new_n265), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n259), .A2(new_n261), .A3(G232), .A4(G1698), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n254), .B1(new_n339), .B2(new_n272), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n279), .A2(G238), .A3(new_n281), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(G179), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n343), .B2(new_n345), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n345), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n344), .B1(new_n340), .B2(new_n341), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n350), .B(new_n347), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n335), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n352), .A2(new_n353), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n335), .B1(new_n357), .B2(G190), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(G200), .C1(new_n352), .C2(new_n353), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n343), .A2(new_n345), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n359), .B1(new_n362), .B2(G200), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n295), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n295), .A2(new_n303), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT7), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n255), .A2(new_n370), .A3(G20), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT7), .B1(new_n262), .B2(new_n213), .ZN(new_n372));
  OAI21_X1  g0172(.A(G68), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n298), .A2(G159), .ZN(new_n374));
  AND3_X1   g0174(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT77), .B1(G58), .B2(G68), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n375), .A2(new_n376), .A3(new_n201), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n374), .B1(new_n377), .B2(new_n213), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n373), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n370), .B1(new_n255), .B2(G20), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n260), .A2(G33), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n384));
  OAI211_X1 g0184(.A(KEYINPUT7), .B(new_n213), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n325), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT16), .B1(new_n386), .B2(new_n378), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n369), .B1(new_n388), .B2(new_n293), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n219), .B1(new_n268), .B2(new_n269), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(new_n275), .A3(new_n277), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT79), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT79), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n390), .A2(new_n275), .A3(new_n393), .A4(new_n277), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n259), .A2(new_n261), .A3(G226), .A4(G1698), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n259), .A2(new_n261), .A3(G223), .A4(new_n265), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(KEYINPUT78), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT78), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n400), .A2(G33), .A3(G87), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n396), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n254), .B1(new_n403), .B2(new_n272), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n319), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(G179), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT18), .B1(new_n389), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n380), .B1(new_n373), .B2(new_n379), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n386), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n293), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n369), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n405), .A2(G179), .ZN(new_n415));
  AOI21_X1  g0215(.A(G169), .B1(new_n395), .B2(new_n404), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n408), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n395), .A2(new_n404), .A3(new_n287), .ZN(new_n420));
  AOI21_X1  g0220(.A(G200), .B1(new_n395), .B2(new_n404), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(G200), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n405), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n395), .A2(new_n404), .A3(new_n287), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT80), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n389), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT81), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n422), .B1(new_n420), .B2(new_n421), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n425), .A2(KEYINPUT80), .A3(new_n426), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n389), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n419), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI22_X1  g0238(.A1(new_n295), .A2(new_n299), .B1(new_n213), .B2(new_n205), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT15), .B(G87), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(new_n296), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n293), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n331), .A2(G77), .A3(new_n309), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n442), .B(new_n443), .C1(G77), .C2(new_n304), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT73), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n282), .A2(G244), .ZN(new_n446));
  INV_X1    g0246(.A(new_n254), .ZN(new_n447));
  INV_X1    g0247(.A(G238), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n256), .A2(new_n448), .B1(new_n220), .B2(new_n255), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n255), .A2(G232), .A3(new_n265), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n450), .A2(KEYINPUT72), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(KEYINPUT72), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n272), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n446), .B(new_n447), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n445), .B1(new_n319), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n455), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n321), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n424), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n445), .B1(new_n455), .B2(new_n287), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR4_X1   g0262(.A1(new_n324), .A2(new_n365), .A3(new_n438), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n259), .A2(new_n261), .A3(G250), .A4(G1698), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n259), .A2(new_n261), .A3(G244), .A4(new_n265), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n272), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n250), .A2(new_n251), .ZN(new_n472));
  INV_X1    g0272(.A(G45), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n473), .A2(G1), .ZN(new_n474));
  INV_X1    g0274(.A(G41), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n474), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(KEYINPUT5), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n252), .B(G45), .C1(new_n475), .C2(KEYINPUT5), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT83), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n472), .A2(new_n476), .A3(new_n477), .A4(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n480), .A3(new_n477), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G257), .A3(new_n276), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n471), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G179), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n299), .A2(new_n205), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT6), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n489), .A3(G107), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n487), .B1(new_n492), .B2(new_n213), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n220), .B1(new_n382), .B2(new_n385), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n293), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n489), .A2(new_n220), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n488), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n490), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n486), .B1(new_n502), .B2(G20), .ZN(new_n503));
  OAI21_X1  g0303(.A(G107), .B1(new_n371), .B2(new_n372), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT82), .A3(new_n293), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n497), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n304), .A2(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n252), .A2(G33), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n331), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n511), .B2(G97), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n485), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT84), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n483), .A2(new_n481), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(new_n471), .ZN(new_n517));
  AND4_X1   g0317(.A1(new_n514), .A2(new_n471), .A3(new_n481), .A4(new_n483), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n319), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n516), .A2(new_n514), .A3(new_n471), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(G190), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n484), .A2(G200), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(new_n507), .A4(new_n512), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n520), .A2(new_n525), .A3(KEYINPUT85), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT86), .B(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n499), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n213), .B1(new_n338), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n255), .A2(new_n213), .A3(G68), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n296), .B2(new_n489), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n293), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n440), .A2(new_n303), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n511), .A2(G87), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n474), .A2(new_n251), .ZN(new_n539));
  INV_X1    g0339(.A(G250), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n473), .B2(G1), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n539), .A2(new_n276), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n255), .A2(G244), .A3(G1698), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n255), .A2(G238), .A3(new_n265), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n542), .B1(new_n546), .B2(new_n272), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n538), .B1(G190), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n424), .B2(new_n547), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n535), .A2(new_n536), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n510), .A2(new_n440), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(new_n321), .B2(new_n547), .ZN(new_n552));
  INV_X1    g0352(.A(new_n547), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n319), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n526), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT21), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n510), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n331), .A2(KEYINPUT87), .A3(G116), .A4(new_n509), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n465), .B(new_n213), .C1(G33), .C2(new_n489), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n560), .A2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n293), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT20), .ZN(new_n567));
  OR2_X1    g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n567), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n302), .A2(G1), .ZN(new_n570));
  INV_X1    g0370(.A(new_n565), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n568), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n255), .A2(G257), .A3(new_n265), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n262), .A2(G303), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n575), .B(new_n576), .C1(new_n256), .C2(new_n221), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n272), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n482), .A2(G270), .A3(new_n276), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n481), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n558), .B1(new_n574), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(G200), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n574), .B(new_n583), .C1(new_n287), .C2(new_n580), .ZN(new_n584));
  INV_X1    g0384(.A(new_n580), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n585), .A2(new_n573), .A3(G179), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n573), .A2(KEYINPUT21), .A3(G169), .A4(new_n580), .ZN(new_n587));
  AND4_X1   g0387(.A1(new_n582), .A2(new_n584), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n482), .A2(G264), .A3(new_n276), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n259), .A2(new_n261), .A3(G257), .A4(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n259), .A2(new_n261), .A3(G250), .A4(new_n265), .ZN(new_n591));
  INV_X1    g0391(.A(G294), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n590), .B(new_n591), .C1(new_n258), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n272), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT89), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n596), .A3(G179), .A4(new_n481), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n589), .A2(new_n594), .A3(new_n481), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT89), .B1(new_n598), .B2(G169), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n321), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n255), .A2(new_n213), .A3(G87), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT22), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT22), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n255), .A2(new_n604), .A3(new_n213), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT24), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT23), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(new_n220), .A3(G20), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT23), .B1(new_n213), .B2(G107), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  OAI221_X1 g0411(.A(new_n609), .B1(G20), .B2(new_n545), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n610), .A2(new_n611), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n606), .A2(new_n607), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n607), .B1(new_n606), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n293), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(KEYINPUT25), .B1(new_n303), .B2(new_n220), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n220), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n511), .A2(G107), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n601), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n598), .A2(new_n424), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n598), .A2(G190), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n617), .B(new_n621), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT82), .B1(new_n505), .B2(new_n293), .ZN(new_n628));
  AOI211_X1 g0428(.A(new_n496), .B(new_n305), .C1(new_n503), .C2(new_n504), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n524), .B(new_n512), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n523), .B1(new_n513), .B2(new_n519), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n588), .B(new_n627), .C1(new_n632), .C2(KEYINPUT85), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n464), .A2(new_n557), .A3(new_n633), .ZN(G372));
  INV_X1    g0434(.A(new_n542), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n546), .A2(KEYINPUT90), .A3(new_n272), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT90), .B1(new_n546), .B2(new_n272), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n319), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n552), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n587), .A2(new_n586), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n582), .ZN(new_n642));
  INV_X1    g0442(.A(new_n623), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(G200), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n552), .A2(new_n639), .B1(new_n548), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n520), .A2(new_n646), .A3(new_n525), .A4(new_n626), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n520), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n650), .A3(new_n646), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n549), .A2(new_n555), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT26), .B1(new_n652), .B2(new_n520), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n463), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n323), .ZN(new_n657));
  INV_X1    g0457(.A(new_n419), .ZN(new_n658));
  INV_X1    g0458(.A(new_n356), .ZN(new_n659));
  INV_X1    g0459(.A(new_n459), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n364), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n434), .A2(new_n389), .A3(new_n435), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n434), .A2(new_n389), .B1(KEYINPUT81), .B2(new_n429), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n658), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n657), .B1(new_n665), .B2(new_n317), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n656), .A2(new_n666), .ZN(G369));
  NAND2_X1  g0467(.A1(new_n570), .A2(new_n213), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT27), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(G213), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n622), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n627), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT91), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n627), .A2(KEYINPUT91), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n673), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n623), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G330), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n588), .B1(new_n574), .B2(new_n680), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n642), .A2(new_n573), .A3(new_n673), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n643), .A2(new_n680), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n673), .B1(new_n641), .B2(new_n582), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n677), .A2(new_n678), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(G399));
  NAND3_X1  g0492(.A1(new_n209), .A2(KEYINPUT92), .A3(new_n475), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT92), .B1(new_n209), .B2(new_n475), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n528), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n216), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n655), .A2(new_n680), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n556), .A2(new_n649), .A3(new_n650), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n548), .A2(new_n645), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n640), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(KEYINPUT26), .B1(new_n707), .B2(new_n520), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n680), .B1(new_n648), .B2(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n547), .A2(new_n589), .A3(new_n594), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n578), .A2(new_n579), .A3(G179), .A4(new_n481), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n522), .A3(new_n521), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n715), .A2(new_n522), .A3(KEYINPUT30), .A4(new_n521), .ZN(new_n719));
  AOI21_X1  g0519(.A(G179), .B1(new_n516), .B2(new_n471), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n580), .A3(new_n598), .A4(new_n638), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT31), .B1(new_n722), .B2(new_n673), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n652), .B1(new_n632), .B2(KEYINPUT85), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n623), .A2(new_n626), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n520), .A2(new_n525), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT85), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n727), .A2(new_n731), .A3(new_n588), .A4(new_n680), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n712), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n702), .B1(new_n735), .B2(new_n252), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT94), .ZN(G364));
  AOI21_X1  g0537(.A(new_n212), .B1(G20), .B2(new_n319), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n287), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n213), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n489), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n213), .A2(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(G190), .A3(G200), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n527), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n213), .A2(new_n321), .ZN(new_n746));
  NOR2_X1   g0546(.A1(G190), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n262), .B1(new_n749), .B2(G77), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n746), .A2(G190), .A3(new_n424), .ZN(new_n751));
  OAI211_X1 g0551(.A(new_n745), .B(new_n750), .C1(new_n218), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n742), .A2(new_n747), .ZN(new_n753));
  INV_X1    g0553(.A(G159), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT32), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n746), .A2(G200), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n287), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n742), .A2(new_n287), .A3(G200), .ZN(new_n760));
  OAI221_X1 g0560(.A(new_n756), .B1(new_n202), .B2(new_n759), .C1(new_n220), .C2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n746), .A2(new_n287), .A3(G200), .ZN(new_n762));
  AND2_X1   g0562(.A1(new_n762), .A2(KEYINPUT97), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n757), .A2(KEYINPUT97), .A3(G190), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n752), .B(new_n761), .C1(G68), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n740), .ZN(new_n767));
  INV_X1    g0567(.A(new_n743), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n767), .A2(G294), .B1(new_n768), .B2(G303), .ZN(new_n769));
  INV_X1    g0569(.A(new_n760), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n758), .A2(G326), .B1(new_n770), .B2(G283), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n753), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n255), .B1(new_n773), .B2(G329), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(new_n775), .B2(new_n748), .C1(new_n776), .C2(new_n751), .ZN(new_n777));
  XNOR2_X1  g0577(.A(KEYINPUT33), .B(G317), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n772), .B(new_n777), .C1(new_n765), .C2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n738), .B1(new_n766), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT96), .Z(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n738), .ZN(new_n784));
  INV_X1    g0584(.A(new_n209), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n255), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n216), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n244), .B2(G45), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n255), .A2(new_n209), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT95), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G355), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(G116), .B2(new_n209), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n784), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n302), .A2(G20), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n252), .B1(new_n794), .B2(G45), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n696), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n780), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT98), .Z(new_n799));
  NAND3_X1  g0599(.A1(new_n685), .A2(new_n686), .A3(new_n783), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n687), .A2(new_n797), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n685), .A2(new_n684), .A3(new_n686), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  AND3_X1   g0606(.A1(new_n456), .A2(new_n458), .A3(new_n680), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n460), .A2(new_n461), .B1(new_n445), .B2(new_n680), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n807), .B1(new_n459), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n782), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n751), .ZN(new_n813));
  XOR2_X1   g0613(.A(KEYINPUT100), .B(G143), .Z(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n813), .A2(new_n815), .B1(new_n749), .B2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(G137), .ZN(new_n817));
  INV_X1    g0617(.A(new_n765), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n817), .B2(new_n759), .C1(new_n818), .C2(new_n297), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n255), .B1(new_n753), .B2(new_n823), .C1(new_n325), .C2(new_n760), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n740), .A2(new_n218), .B1(new_n743), .B2(new_n202), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n821), .A2(new_n822), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G87), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n827), .A2(new_n760), .B1(new_n743), .B2(new_n220), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n741), .B(new_n828), .C1(G303), .C2(new_n758), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n751), .A2(new_n592), .B1(new_n753), .B2(new_n775), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n255), .B(new_n830), .C1(G116), .C2(new_n749), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n829), .B(new_n831), .C1(new_n832), .C2(new_n818), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT99), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n738), .B1(new_n826), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n738), .A2(new_n781), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n205), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n812), .A2(new_n797), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n703), .A2(new_n810), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n680), .B(new_n809), .C1(new_n648), .C2(new_n654), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(new_n734), .ZN(new_n842));
  INV_X1    g0642(.A(new_n797), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n841), .A2(new_n734), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n838), .B1(new_n846), .B2(new_n847), .ZN(G384));
  NOR2_X1   g0648(.A1(new_n794), .A2(new_n252), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n413), .B1(new_n432), .B2(new_n433), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n389), .B1(new_n407), .B2(new_n671), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n671), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n413), .B1(new_n417), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n850), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n428), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n389), .A2(new_n671), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(KEYINPUT38), .C1(new_n437), .C2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT104), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n664), .B2(new_n419), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT104), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT38), .A4(new_n858), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n431), .A2(new_n436), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n860), .B1(new_n867), .B2(new_n658), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n853), .A2(new_n857), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n862), .A2(new_n865), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n335), .A2(new_n673), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n356), .A2(new_n364), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n356), .A2(new_n364), .A3(KEYINPUT102), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n351), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n364), .A2(new_n354), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n335), .A3(new_n673), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n810), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT106), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n633), .A2(new_n557), .A3(new_n673), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n722), .A2(new_n673), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT31), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n723), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n882), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n726), .A2(new_n732), .A3(KEYINPUT106), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n871), .A2(new_n881), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT107), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n891), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT105), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT37), .B1(new_n852), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n428), .A2(new_n855), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n428), .A2(new_n855), .A3(new_n897), .A4(KEYINPUT37), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n866), .B1(new_n868), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n891), .B1(new_n903), .B2(new_n861), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(new_n881), .A3(new_n888), .A4(new_n889), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n463), .A2(new_n888), .A3(new_n889), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n908), .A2(new_n909), .A3(new_n684), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n861), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n862), .A2(new_n865), .A3(new_n870), .A4(KEYINPUT39), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n356), .A2(new_n673), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n807), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n840), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n877), .A2(new_n880), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n922), .A2(new_n871), .B1(new_n419), .B2(new_n671), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n463), .B1(new_n704), .B2(new_n711), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n925), .A2(new_n666), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n924), .B(new_n926), .Z(new_n927));
  AOI21_X1  g0727(.A(new_n849), .B1(new_n911), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n927), .B2(new_n911), .ZN(new_n929));
  AOI211_X1 g0729(.A(new_n560), .B(new_n215), .C1(new_n502), .C2(KEYINPUT35), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(KEYINPUT35), .B2(new_n502), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n376), .A2(new_n375), .A3(new_n216), .A4(new_n205), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n325), .A2(G50), .ZN(new_n934));
  OAI211_X1 g0734(.A(G1), .B(new_n302), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n932), .A3(new_n935), .ZN(G367));
  NAND2_X1  g0736(.A1(new_n507), .A2(new_n512), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n673), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n632), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n520), .B2(new_n680), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n691), .A2(new_n689), .A3(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n940), .B1(new_n691), .B2(new_n689), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(KEYINPUT44), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n944), .A2(KEYINPUT44), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n943), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n688), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n943), .B(new_n688), .C1(new_n945), .C2(new_n946), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n691), .B1(new_n683), .B2(new_n690), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(new_n687), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n734), .A3(new_n712), .ZN(new_n954));
  OAI21_X1  g0754(.A(KEYINPUT109), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n954), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT109), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n956), .A2(new_n949), .A3(new_n957), .A4(new_n950), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n735), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n696), .B(KEYINPUT41), .Z(new_n960));
  OAI21_X1  g0760(.A(new_n795), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n940), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n691), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n520), .B1(new_n939), .B2(new_n623), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n963), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n538), .A2(new_n673), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n646), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n640), .A2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n964), .A2(new_n966), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n948), .A2(new_n940), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n961), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n784), .B1(new_n209), .B2(new_n440), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n239), .A2(new_n786), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n797), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G50), .A2(new_n749), .B1(new_n773), .B2(G137), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n980), .B(new_n255), .C1(new_n297), .C2(new_n751), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n760), .A2(new_n205), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n758), .B2(new_n815), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n218), .B2(new_n743), .C1(new_n325), .C2(new_n740), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n981), .B(new_n984), .C1(G159), .C2(new_n765), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G283), .A2(new_n749), .B1(new_n773), .B2(G317), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n255), .B1(new_n813), .B2(G303), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n768), .A2(KEYINPUT46), .A3(G116), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT46), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n743), .B2(new_n560), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G107), .A2(new_n767), .B1(new_n758), .B2(G311), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n489), .B2(new_n760), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n991), .B(new_n993), .C1(G294), .C2(new_n765), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n979), .B1(new_n996), .B2(new_n738), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n968), .A2(new_n969), .A3(new_n783), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n976), .A2(new_n999), .ZN(G387));
  INV_X1    g0800(.A(new_n698), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n790), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(G107), .B2(new_n209), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n236), .A2(G45), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1004), .B(KEYINPUT110), .Z(new_n1005));
  INV_X1    g0805(.A(new_n786), .ZN(new_n1006));
  AOI211_X1 g0806(.A(G45), .B(new_n1001), .C1(G68), .C2(G77), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n295), .A2(G50), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1003), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n784), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n797), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT111), .Z(new_n1014));
  INV_X1    g0814(.A(new_n783), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(KEYINPUT112), .B(G150), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n813), .A2(G50), .B1(new_n773), .B2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n255), .C1(new_n325), .C2(new_n748), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n740), .A2(new_n440), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n743), .A2(new_n205), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n489), .B2(new_n760), .C1(new_n754), .C2(new_n759), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1018), .B(new_n1022), .C1(new_n366), .C2(new_n765), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT113), .Z(new_n1024));
  AOI22_X1  g0824(.A1(new_n813), .A2(G317), .B1(new_n749), .B2(G303), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n776), .B2(new_n759), .C1(new_n818), .C2(new_n775), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT115), .Z(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(KEYINPUT48), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1027), .A2(KEYINPUT48), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n740), .A2(new_n832), .B1(new_n743), .B2(new_n592), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT114), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT49), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n255), .B1(new_n773), .B2(G326), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n560), .B2(new_n760), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT116), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1032), .B2(KEYINPUT49), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1024), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n738), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1014), .B1(new_n683), .B2(new_n1015), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT117), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n953), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n735), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1043), .A2(new_n696), .A3(new_n954), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1041), .B(new_n1044), .C1(new_n795), .C2(new_n1042), .ZN(G393));
  INV_X1    g0845(.A(KEYINPUT118), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n795), .B1(new_n951), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n951), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n784), .B1(new_n489), .B2(new_n209), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n247), .A2(new_n1006), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n797), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n255), .B1(new_n814), .B2(new_n753), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n366), .B2(new_n749), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n740), .A2(new_n205), .B1(new_n760), .B2(new_n827), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G68), .B2(new_n768), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(new_n818), .C2(new_n202), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G150), .A2(new_n758), .B1(new_n813), .B2(G159), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT51), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n765), .A2(G303), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n262), .B1(new_n753), .B2(new_n776), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G294), .B2(new_n749), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n220), .A2(new_n760), .B1(new_n743), .B2(new_n832), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G116), .B2(new_n767), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G317), .A2(new_n758), .B1(new_n813), .B2(G311), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1056), .A2(new_n1058), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1051), .B1(new_n1067), .B2(new_n738), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n940), .B2(new_n1015), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1048), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n955), .A2(new_n958), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT119), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n697), .B1(new_n951), .B2(new_n954), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1073), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1071), .B1(new_n1076), .B2(new_n1077), .ZN(G390));
  NAND2_X1  g0878(.A1(new_n808), .A2(new_n459), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n919), .B1(new_n710), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n921), .A2(new_n733), .A3(G330), .A4(new_n809), .ZN(new_n1083));
  AND4_X1   g0883(.A1(G330), .A2(new_n888), .A3(new_n809), .A4(new_n889), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1083), .C1(new_n1084), .C2(new_n921), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n921), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n734), .B2(new_n810), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n888), .A2(new_n881), .A3(G330), .A4(new_n889), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n920), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1085), .A2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n463), .A2(G330), .A3(new_n888), .A4(new_n889), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n925), .A2(new_n666), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n917), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n912), .C1(new_n1082), .C2(new_n1086), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1083), .C1(new_n916), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1088), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n920), .A2(new_n921), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1100), .A2(new_n1095), .B1(new_n914), .B2(new_n915), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n912), .A2(new_n1095), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n921), .B2(new_n1081), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1099), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1094), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1091), .A2(new_n1093), .A3(new_n1098), .A4(new_n1104), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n696), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1098), .A2(new_n796), .A3(new_n1104), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n836), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n797), .B1(new_n366), .B2(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n751), .A2(new_n560), .B1(new_n753), .B2(new_n592), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n255), .B(new_n1112), .C1(G97), .C2(new_n749), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n765), .A2(G107), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n767), .A2(G77), .B1(new_n770), .B2(G68), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n758), .A2(G283), .B1(new_n768), .B2(G87), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n768), .A2(new_n1016), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT53), .Z(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n818), .B2(new_n817), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G159), .A2(new_n767), .B1(new_n758), .B2(G128), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n262), .B1(new_n749), .B2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n813), .A2(G132), .B1(new_n773), .B2(G125), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n770), .A2(G50), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1121), .A2(new_n1124), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1117), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1111), .B1(new_n1128), .B2(new_n738), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n916), .B2(new_n782), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1108), .A2(new_n1109), .A3(new_n1130), .ZN(G378));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n1107), .B2(new_n1093), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n905), .A2(G330), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n891), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT107), .B1(new_n890), .B2(new_n891), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n657), .B1(new_n314), .B2(new_n316), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n312), .A2(new_n854), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT55), .Z(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1140), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1147), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(new_n1139), .A3(new_n1145), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1138), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n924), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1151), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n1135), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1133), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n696), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT123), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1107), .A2(new_n1093), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1154), .B1(new_n896), .B2(new_n1135), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1134), .B(new_n1151), .C1(new_n894), .C2(new_n895), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n924), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(KEYINPUT123), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1161), .A2(new_n1162), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1159), .B1(new_n1168), .B2(new_n1132), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1161), .A2(new_n796), .A3(new_n1167), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1151), .A2(new_n811), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n797), .B1(G50), .B2(new_n1110), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n770), .A2(G58), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n759), .B2(new_n560), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1020), .B(new_n1174), .C1(G68), .C2(new_n767), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n262), .A2(new_n475), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n748), .A2(new_n440), .B1(new_n753), .B2(new_n832), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G107), .C2(new_n813), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(new_n489), .C2(new_n818), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT58), .ZN(new_n1180));
  AOI21_X1  g0980(.A(G50), .B1(new_n258), .B2(new_n475), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1179), .A2(new_n1180), .B1(new_n1176), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(G128), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n751), .A2(new_n1183), .B1(new_n748), .B2(new_n817), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(G150), .B2(new_n767), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n758), .A2(G125), .B1(new_n768), .B2(new_n1123), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n818), .C2(new_n823), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT59), .Z(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1189), .A2(KEYINPUT120), .ZN(new_n1190));
  AOI211_X1 g0990(.A(G33), .B(G41), .C1(new_n773), .C2(G124), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n754), .B2(new_n760), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT121), .Z(new_n1193));
  INV_X1    g0993(.A(KEYINPUT120), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1193), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1182), .B1(new_n1180), .B2(new_n1179), .C1(new_n1190), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1172), .B1(new_n1196), .B2(new_n738), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1171), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1170), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1169), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(G375));
  INV_X1    g1001(.A(new_n1091), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1093), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n960), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1094), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n255), .B1(new_n773), .B2(G303), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n220), .B2(new_n748), .C1(new_n832), .C2(new_n751), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n759), .A2(new_n592), .B1(new_n743), .B2(new_n489), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1208), .A2(new_n1209), .A3(new_n982), .A4(new_n1019), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n765), .A2(G116), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n759), .A2(KEYINPUT124), .A3(new_n823), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT124), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n758), .B2(G132), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n255), .B1(new_n748), .B2(new_n297), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n751), .A2(new_n817), .B1(new_n753), .B2(new_n1183), .ZN(new_n1216));
  NOR4_X1   g1016(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1173), .B1(new_n754), .B2(new_n743), .C1(new_n202), .C2(new_n740), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n765), .B2(new_n1123), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1210), .A2(new_n1211), .B1(new_n1217), .B2(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n797), .B1(G68), .B2(new_n1110), .C1(new_n1220), .C2(new_n1039), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1086), .B2(new_n781), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1202), .B2(new_n795), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1206), .A2(new_n1225), .ZN(G381));
  AOI22_X1  g1026(.A1(new_n961), .A2(new_n975), .B1(new_n998), .B2(new_n997), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1077), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1070), .B1(new_n1228), .B2(new_n1075), .ZN(new_n1229));
  OR2_X1    g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1230), .A2(G378), .A3(G381), .A4(G384), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1200), .A2(new_n1227), .A3(new_n1229), .A4(new_n1231), .ZN(G407));
  NAND2_X1  g1032(.A1(new_n672), .A2(G213), .ZN(new_n1233));
  OR2_X1    g1033(.A1(G378), .A2(new_n1233), .ZN(new_n1234));
  OAI211_X1 g1034(.A(G407), .B(G213), .C1(G375), .C2(new_n1234), .ZN(G409));
  NAND2_X1  g1035(.A1(G387), .A2(new_n1229), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1227), .A2(G390), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(G393), .B(new_n805), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1236), .A2(new_n1239), .A3(new_n1237), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT63), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1202), .A2(KEYINPUT60), .A3(new_n1203), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1245), .A2(new_n696), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1204), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1224), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(G384), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(G384), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G378), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1169), .A2(new_n1254), .A3(new_n1199), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n795), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1171), .B2(new_n1197), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1161), .A2(new_n1167), .A3(new_n1205), .A4(new_n1162), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G378), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1233), .B(new_n1253), .C1(new_n1255), .C2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1243), .B1(new_n1244), .B2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n672), .A2(G213), .A3(G2897), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT125), .Z(new_n1263));
  XNOR2_X1  g1063(.A(new_n1252), .B(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1233), .B1(new_n1255), .B2(new_n1259), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1261), .B(new_n1266), .C1(new_n1244), .C2(new_n1260), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1168), .A2(new_n1132), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1159), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1199), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1270), .A2(G378), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1259), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1272), .A2(new_n1273), .B1(G213), .B2(new_n672), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT62), .B1(new_n1274), .B2(new_n1253), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT62), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1260), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(KEYINPUT126), .B(new_n1266), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1243), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1274), .A2(KEYINPUT62), .A3(new_n1253), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1260), .A2(new_n1276), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT126), .B1(new_n1282), .B2(new_n1266), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1267), .B1(new_n1279), .B2(new_n1283), .ZN(G405));
  INV_X1    g1084(.A(new_n1242), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1239), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1252), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1253), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT127), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1200), .A2(G378), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(new_n1255), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1252), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1241), .A2(new_n1253), .A3(new_n1242), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n1289), .A2(new_n1291), .A3(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1291), .B1(new_n1289), .B2(new_n1295), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(new_n1297), .ZN(G402));
endmodule


