//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G122), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT3), .A2(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT3), .A2(G107), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(G104), .B2(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(KEYINPUT3), .A2(G107), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT79), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G104), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n196), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n198), .B1(G104), .B2(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n199), .A2(KEYINPUT80), .A3(new_n203), .ZN(new_n208));
  XNOR2_X1  g022(.A(G116), .B(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT5), .ZN(new_n210));
  INV_X1    g024(.A(G116), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT5), .A3(G119), .ZN(new_n212));
  INV_X1    g026(.A(G113), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n210), .A2(new_n214), .B1(new_n216), .B2(new_n209), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n217), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n192), .A2(new_n194), .A3(new_n196), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT3), .A2(G107), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n192), .B2(new_n193), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT4), .A3(new_n199), .ZN(new_n223));
  INV_X1    g037(.A(new_n209), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT69), .A3(new_n215), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT69), .B1(new_n216), .B2(new_n209), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n215), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n229), .B(G101), .C1(new_n219), .C2(new_n221), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n223), .A2(new_n225), .A3(new_n228), .A4(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n218), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n206), .A2(new_n208), .A3(new_n217), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT81), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n188), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT6), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n188), .A3(new_n231), .A4(new_n218), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT82), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n232), .A2(new_n240), .A3(new_n188), .A4(new_n234), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n237), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n236), .B1(new_n242), .B2(new_n235), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT65), .B(G143), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(G146), .ZN(new_n248));
  INV_X1    g062(.A(G143), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G146), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT1), .ZN(new_n251));
  OAI21_X1  g065(.A(G128), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n250), .B1(new_n247), .B2(G146), .ZN(new_n254));
  INV_X1    g068(.A(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT1), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G125), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n249), .A2(KEYINPUT65), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT65), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n245), .B1(new_n265), .B2(new_n244), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NOR3_X1   g083(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n261), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n267), .ZN(new_n273));
  OR3_X1    g087(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(new_n268), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n248), .A2(new_n275), .A3(KEYINPUT66), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n272), .A2(new_n276), .B1(new_n273), .B2(new_n254), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n260), .B1(new_n259), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G953), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G224), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n278), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n243), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G210), .B1(G237), .B2(G902), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n199), .A2(new_n203), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n233), .B1(new_n285), .B2(new_n217), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n188), .B(KEYINPUT8), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT84), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n289), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n290), .B2(new_n281), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n288), .B1(new_n278), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n278), .B1(new_n289), .B2(new_n281), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n278), .B(KEYINPUT83), .C1(new_n289), .C2(new_n281), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n239), .A2(new_n241), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n283), .A2(new_n284), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n284), .B1(new_n283), .B2(new_n300), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n187), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OR2_X1    g117(.A1(new_n303), .A2(KEYINPUT85), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n305));
  XNOR2_X1  g119(.A(G113), .B(G122), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(new_n193), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n259), .A2(G140), .ZN(new_n310));
  INV_X1    g124(.A(G140), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G125), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT19), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n259), .A2(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT74), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT88), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n313), .A2(KEYINPUT88), .A3(new_n314), .A4(new_n317), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT19), .B1(new_n310), .B2(new_n312), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n320), .A2(new_n244), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT16), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n310), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(G146), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n329));
  INV_X1    g143(.A(G237), .ZN(new_n330));
  AND4_X1   g144(.A1(G143), .A2(new_n330), .A3(new_n279), .A4(G214), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n279), .A3(G214), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n247), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G131), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n262), .A3(new_n264), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n279), .A3(G143), .A4(G214), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT86), .A3(G131), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n333), .A2(new_n334), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n335), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT87), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT86), .B1(new_n338), .B2(G131), .ZN(new_n343));
  AOI211_X1 g157(.A(new_n329), .B(new_n334), .C1(new_n336), .C2(new_n337), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT87), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n340), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n328), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(KEYINPUT18), .A2(G131), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n338), .B(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n313), .A2(new_n244), .A3(new_n317), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n244), .B1(new_n315), .B2(new_n316), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n308), .B1(new_n348), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT17), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n335), .A2(new_n358), .A3(new_n339), .A4(new_n340), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n324), .A2(G146), .A3(new_n326), .ZN(new_n360));
  AOI21_X1  g174(.A(G146), .B1(new_n324), .B2(new_n326), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT17), .B1(new_n343), .B2(new_n344), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n355), .A3(new_n307), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n357), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n305), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  AOI211_X1 g183(.A(KEYINPUT20), .B(new_n369), .C1(new_n357), .C2(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n364), .A2(new_n355), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n308), .ZN(new_n372));
  AOI21_X1  g186(.A(G902), .B1(new_n372), .B2(new_n365), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(KEYINPUT89), .ZN(new_n374));
  INV_X1    g188(.A(G902), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n364), .A2(new_n307), .A3(new_n355), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n307), .B1(new_n364), .B2(new_n355), .ZN(new_n377));
  OAI211_X1 g191(.A(KEYINPUT89), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G475), .ZN(new_n379));
  OAI22_X1  g193(.A1(new_n368), .A2(new_n370), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(KEYINPUT9), .B(G234), .ZN(new_n381));
  INV_X1    g195(.A(G217), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n381), .A2(new_n382), .A3(G953), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n384));
  INV_X1    g198(.A(G122), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G116), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n211), .A2(G122), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT90), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n386), .B2(new_n387), .ZN(new_n390));
  OAI21_X1  g204(.A(G107), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(new_n387), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT90), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(new_n200), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n249), .A2(G128), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n397), .B1(new_n247), .B2(G128), .ZN(new_n398));
  INV_X1    g212(.A(G134), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n262), .A2(new_n264), .A3(G128), .ZN(new_n401));
  INV_X1    g215(.A(new_n397), .ZN(new_n402));
  AND3_X1   g216(.A1(new_n401), .A2(KEYINPUT13), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT13), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n262), .A2(new_n264), .A3(new_n404), .A4(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G134), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n400), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n384), .B1(new_n396), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n406), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(KEYINPUT13), .A3(new_n402), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n409), .A2(new_n410), .B1(new_n399), .B2(new_n398), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n391), .A2(new_n395), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(KEYINPUT91), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n200), .B1(new_n386), .B2(KEYINPUT14), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n415), .A2(new_n392), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n392), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n398), .A2(new_n399), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n400), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n383), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n383), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n423), .B(new_n420), .C1(new_n408), .C2(new_n413), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n375), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT15), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(G478), .ZN(new_n427));
  INV_X1    g241(.A(G478), .ZN(new_n428));
  OAI221_X1 g242(.A(new_n375), .B1(KEYINPUT15), .B2(new_n428), .C1(new_n422), .C2(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT21), .B(G898), .Z(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT92), .ZN(new_n432));
  AOI211_X1 g246(.A(new_n375), .B(new_n279), .C1(G234), .C2(G237), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n279), .A2(G952), .ZN(new_n436));
  INV_X1    g250(.A(G234), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n330), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT93), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n380), .A2(new_n430), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n303), .A2(KEYINPUT85), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT67), .ZN(new_n445));
  INV_X1    g259(.A(G137), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(KEYINPUT67), .A2(G137), .ZN(new_n448));
  AND2_X1   g262(.A1(KEYINPUT11), .A2(G134), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(KEYINPUT11), .A2(G134), .ZN(new_n451));
  NOR2_X1   g265(.A1(KEYINPUT11), .A2(G134), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n451), .B1(new_n452), .B2(G137), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n334), .A2(KEYINPUT68), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n455), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n450), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n254), .A2(new_n273), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n266), .A2(new_n271), .A3(new_n261), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT66), .B1(new_n248), .B2(new_n275), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n253), .A2(new_n257), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n450), .A2(new_n453), .A3(new_n334), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n447), .A2(new_n399), .A3(new_n448), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n334), .B1(G134), .B2(G137), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n464), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n228), .A2(new_n225), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT28), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n465), .A2(new_n468), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n475), .B1(new_n253), .B2(new_n257), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT70), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n450), .A2(new_n457), .A3(new_n453), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n457), .B1(new_n450), .B2(new_n453), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n456), .A2(KEYINPUT70), .A3(new_n458), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n476), .B1(new_n482), .B2(new_n277), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n474), .B1(new_n483), .B2(new_n471), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n272), .A2(new_n276), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n485), .A2(new_n460), .A3(new_n481), .A4(new_n480), .ZN(new_n486));
  AND4_X1   g300(.A1(new_n474), .A2(new_n486), .A3(new_n471), .A4(new_n469), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n473), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n489));
  NAND3_X1  g303(.A1(new_n330), .A2(new_n279), .A3(G210), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT26), .B(G101), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n491), .B(new_n492), .Z(new_n493));
  NAND2_X1  g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n470), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n486), .A2(KEYINPUT30), .A3(new_n469), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n472), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n483), .A2(new_n471), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT31), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT31), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n498), .A2(new_n504), .A3(new_n499), .A4(new_n501), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n494), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(G472), .A2(G902), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n506), .A2(KEYINPUT32), .A3(new_n507), .ZN(new_n511));
  INV_X1    g325(.A(new_n493), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n488), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n498), .A2(new_n499), .A3(new_n493), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT29), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n484), .A2(new_n487), .B1(new_n471), .B2(new_n483), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(KEYINPUT29), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n375), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G472), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n510), .A2(new_n511), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G469), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n277), .A2(new_n230), .A3(new_n223), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n254), .B1(G128), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n254), .A2(new_n256), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n285), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n480), .A2(new_n481), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n206), .A2(new_n464), .A3(KEYINPUT10), .A4(new_n208), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n522), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n464), .B1(new_n206), .B2(new_n208), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n523), .A2(G128), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n265), .A2(new_n244), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n250), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n204), .B1(new_n536), .B2(new_n257), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n532), .B(new_n482), .C1(new_n533), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n208), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT80), .B1(new_n199), .B2(new_n203), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n258), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n526), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n532), .B1(new_n543), .B2(new_n459), .ZN(new_n544));
  XOR2_X1   g358(.A(G110), .B(G140), .Z(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT78), .ZN(new_n546));
  INV_X1    g360(.A(G227), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(G953), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n546), .B(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n539), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n549), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n522), .A2(new_n528), .A3(new_n530), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n482), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n551), .B1(new_n553), .B2(new_n531), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n521), .B(new_n375), .C1(new_n550), .C2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n521), .A2(new_n375), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n549), .B1(new_n539), .B2(new_n544), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n553), .A2(new_n531), .A3(new_n551), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n555), .B(new_n557), .C1(new_n521), .C2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G221), .B1(new_n381), .B2(G902), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT77), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT75), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(G119), .A3(new_n255), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n255), .A2(G119), .ZN(new_n572));
  INV_X1    g386(.A(G119), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G128), .ZN(new_n574));
  AND2_X1   g388(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n572), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n571), .A2(G110), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n568), .B(new_n577), .C1(new_n360), .C2(new_n361), .ZN(new_n578));
  AOI21_X1  g392(.A(G110), .B1(new_n571), .B2(new_n576), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n566), .A2(new_n567), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n351), .B(new_n327), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT22), .B(G137), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n279), .A2(G221), .A3(G234), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n578), .A2(new_n581), .A3(new_n585), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n587), .A2(new_n375), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n565), .B1(new_n589), .B2(KEYINPUT25), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT76), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n591), .A3(KEYINPUT25), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n587), .A2(KEYINPUT25), .A3(new_n375), .A4(new_n588), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n375), .A3(new_n588), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT25), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n590), .A2(new_n592), .A3(new_n594), .A4(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n382), .B1(G234), .B2(new_n375), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n587), .A2(new_n588), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n599), .A2(G902), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n520), .A2(new_n564), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n304), .A2(new_n443), .A3(new_n444), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(KEYINPUT94), .A2(G472), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n506), .A2(new_n375), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n506), .A2(new_n375), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(KEYINPUT94), .A3(G472), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n564), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n604), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n187), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n283), .A2(new_n300), .ZN(new_n616));
  INV_X1    g430(.A(new_n284), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n283), .A2(new_n300), .A3(new_n284), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n615), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT33), .B1(new_n422), .B2(new_n424), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n396), .A2(new_n407), .A3(new_n384), .ZN(new_n622));
  AOI21_X1  g436(.A(KEYINPUT91), .B1(new_n411), .B2(new_n412), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n421), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n423), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n414), .A2(new_n421), .A3(new_n383), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n621), .A2(new_n628), .A3(G478), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n428), .B(new_n375), .C1(new_n422), .C2(new_n424), .ZN(new_n630));
  NAND2_X1  g444(.A1(G478), .A2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n323), .A2(new_n327), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n346), .B1(new_n345), .B2(new_n340), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n346), .A2(new_n335), .A3(new_n339), .A4(new_n340), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n633), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n355), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n376), .B1(new_n637), .B2(new_n308), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT20), .B1(new_n638), .B2(new_n369), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n366), .A2(new_n305), .A3(new_n367), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT89), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(G475), .A3(new_n378), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n632), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n614), .A2(new_n441), .A3(new_n620), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT34), .B(G104), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(G475), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n373), .B2(KEYINPUT89), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n639), .A2(new_n640), .B1(new_n651), .B2(new_n644), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n620), .A2(new_n652), .A3(new_n430), .A4(new_n441), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n613), .A3(new_n612), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G107), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT95), .B(KEYINPUT35), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n586), .A2(KEYINPUT36), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n582), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n602), .ZN(new_n661));
  AOI21_X1  g475(.A(KEYINPUT96), .B1(new_n600), .B2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT96), .ZN(new_n663));
  INV_X1    g477(.A(new_n661), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n663), .B(new_n664), .C1(new_n598), .C2(new_n599), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n658), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n599), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n595), .A2(KEYINPUT75), .A3(new_n596), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT75), .B1(new_n595), .B2(new_n596), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n593), .B(new_n591), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n663), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n600), .A2(KEYINPUT96), .A3(new_n661), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(KEYINPUT97), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n612), .B1(new_n666), .B2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n444), .A3(new_n443), .A4(new_n304), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G12));
  INV_X1    g493(.A(KEYINPUT98), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n430), .B(new_n645), .C1(new_n368), .C2(new_n370), .ZN(new_n681));
  INV_X1    g495(.A(G900), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n433), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n438), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n680), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n652), .A2(KEYINPUT98), .A3(new_n430), .A4(new_n684), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n561), .A2(new_n563), .ZN(new_n689));
  AND3_X1   g503(.A1(new_n506), .A2(KEYINPUT32), .A3(new_n507), .ZN(new_n690));
  AOI21_X1  g504(.A(KEYINPUT32), .B1(new_n506), .B2(new_n507), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n689), .B1(new_n692), .B2(new_n519), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n666), .A2(new_n675), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n688), .A2(new_n693), .A3(new_n620), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NAND2_X1  g510(.A1(new_n499), .A2(new_n493), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n483), .A2(new_n471), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n375), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n510), .A2(new_n511), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT100), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n510), .A2(new_n704), .A3(new_n511), .A4(new_n701), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n684), .B(KEYINPUT39), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n564), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT40), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n673), .A2(new_n674), .ZN(new_n710));
  INV_X1    g524(.A(new_n430), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n710), .A2(new_n652), .A3(new_n711), .A4(new_n615), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n301), .A2(new_n302), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n706), .A2(new_n709), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n247), .ZN(G45));
  NAND2_X1  g531(.A1(new_n646), .A2(new_n684), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n693), .A2(new_n620), .A3(new_n694), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  OAI21_X1  g535(.A(new_n375), .B1(new_n550), .B2(new_n554), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G469), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n723), .A2(new_n555), .A3(new_n562), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n520), .A2(new_n604), .A3(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n646), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n725), .A2(new_n303), .A3(new_n442), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT41), .B(G113), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT101), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n727), .B(new_n729), .ZN(G15));
  OR3_X1    g544(.A1(new_n653), .A2(KEYINPUT102), .A3(new_n725), .ZN(new_n731));
  OAI21_X1  g545(.A(KEYINPUT102), .B1(new_n653), .B2(new_n725), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  OAI211_X1 g548(.A(new_n724), .B(new_n187), .C1(new_n301), .C2(new_n302), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n443), .A3(new_n520), .A4(new_n694), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  NAND2_X1  g552(.A1(new_n610), .A2(G472), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n516), .A2(new_n493), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n503), .A3(new_n505), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n507), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n604), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n724), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n442), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT103), .B1(new_n652), .B2(new_n711), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT103), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n380), .A2(new_n747), .A3(new_n430), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n303), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G122), .ZN(G24));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n646), .B2(new_n684), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n755));
  AND4_X1   g569(.A1(new_n753), .A2(new_n380), .A3(new_n755), .A4(new_n684), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n710), .A2(new_n742), .A3(new_n739), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n736), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  INV_X1    g575(.A(new_n562), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n555), .A2(new_n557), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT105), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n559), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(G469), .A3(new_n558), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n762), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n713), .A2(new_n187), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n613), .B1(new_n692), .B2(new_n519), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n757), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT42), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n769), .A2(KEYINPUT42), .A3(new_n770), .A4(new_n757), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NAND3_X1  g590(.A1(new_n769), .A2(new_n688), .A3(new_n770), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n652), .A2(new_n755), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT43), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n611), .A2(new_n609), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n710), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT44), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n301), .A2(new_n302), .A3(new_n615), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n783), .B2(KEYINPUT44), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n766), .A2(KEYINPUT45), .A3(new_n558), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n521), .B1(new_n560), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n556), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n555), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT46), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT106), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n762), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n707), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n788), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n446), .ZN(G39));
  NOR3_X1   g616(.A1(new_n520), .A2(new_n718), .A3(new_n604), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n785), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n799), .A2(KEYINPUT47), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n798), .B2(new_n762), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n804), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(new_n311), .ZN(G42));
  NOR4_X1   g623(.A1(new_n780), .A2(new_n786), .A3(new_n438), .A4(new_n744), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n770), .ZN(new_n811));
  XOR2_X1   g625(.A(new_n811), .B(KEYINPUT48), .Z(new_n812));
  OR3_X1    g626(.A1(new_n780), .A2(new_n438), .A3(new_n743), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n706), .A2(new_n438), .A3(new_n613), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n724), .A3(new_n785), .ZN(new_n815));
  OAI221_X1 g629(.A(new_n436), .B1(new_n813), .B2(new_n735), .C1(new_n815), .C2(new_n726), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  OR4_X1    g632(.A1(new_n187), .A2(new_n813), .A3(new_n715), .A4(new_n744), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n818), .B1(new_n821), .B2(KEYINPUT114), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n815), .A2(new_n380), .A3(new_n755), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n810), .A2(new_n759), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT113), .B1(new_n818), .B2(KEYINPUT114), .ZN(new_n825));
  AOI211_X1 g639(.A(new_n823), .B(new_n824), .C1(new_n819), .C2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n826), .A3(KEYINPUT115), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n723), .A2(new_n555), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n805), .B(new_n807), .C1(new_n563), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n813), .A2(new_n786), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n827), .A2(KEYINPUT51), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT115), .B1(new_n822), .B2(new_n826), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n822), .A2(new_n826), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n830), .B2(new_n831), .ZN(new_n836));
  OAI221_X1 g650(.A(new_n817), .B1(new_n833), .B2(new_n834), .C1(KEYINPUT51), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n737), .A2(new_n751), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n727), .ZN(new_n839));
  AND4_X1   g653(.A1(KEYINPUT53), .A2(new_n733), .A3(new_n775), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n430), .B(KEYINPUT107), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(new_n380), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n442), .B1(new_n842), .B2(new_n726), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n304), .A3(new_n614), .A4(new_n444), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n677), .A2(new_n606), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n652), .A2(new_n684), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n841), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT108), .B1(new_n786), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n694), .A2(new_n520), .A3(new_n564), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT108), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n785), .A2(new_n851), .A3(new_n841), .A4(new_n847), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n754), .A2(new_n758), .A3(new_n756), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n769), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n853), .A2(new_n777), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n845), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n677), .A2(new_n606), .A3(new_n844), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n853), .A2(new_n777), .A3(new_n855), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT112), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n840), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n672), .A2(new_n664), .A3(new_n685), .ZN(new_n864));
  INV_X1    g678(.A(new_n767), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n864), .B(new_n562), .C1(new_n865), .C2(new_n763), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n704), .B1(new_n692), .B2(new_n701), .ZN(new_n868));
  INV_X1    g682(.A(new_n705), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n620), .A2(new_n746), .A3(new_n748), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n760), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n695), .A2(new_n720), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT110), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n866), .B1(new_n703), .B2(new_n705), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n750), .A2(new_n876), .B1(new_n854), .B2(new_n736), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n850), .B(new_n620), .C1(new_n688), .C2(new_n719), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT110), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n863), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT52), .B1(new_n872), .B2(new_n873), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n862), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n874), .B1(new_n872), .B2(new_n873), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n877), .A2(KEYINPUT110), .A3(new_n878), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT52), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT111), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n845), .A2(new_n856), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n775), .A2(new_n733), .A3(new_n839), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT111), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n885), .A2(new_n886), .A3(KEYINPUT52), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n880), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n889), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n883), .B1(new_n884), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT109), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n900), .B1(new_n890), .B2(new_n891), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n733), .A2(new_n839), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n859), .A2(new_n860), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT109), .A4(new_n775), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n884), .B1(new_n905), .B2(new_n882), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n884), .B2(new_n896), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n899), .B1(new_n908), .B2(new_n898), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n837), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(G952), .A2(G953), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n828), .B(KEYINPUT49), .Z(new_n912));
  NAND3_X1  g726(.A1(new_n604), .A2(new_n187), .A3(new_n563), .ZN(new_n913));
  OR4_X1    g727(.A1(new_n706), .A2(new_n912), .A3(new_n779), .A4(new_n913), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n910), .A2(new_n911), .B1(new_n715), .B2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n897), .A2(new_n375), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(G210), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT56), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n243), .B(new_n282), .ZN(new_n919));
  XOR2_X1   g733(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n917), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(new_n917), .B2(new_n918), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n279), .A2(G952), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(G51));
  XNOR2_X1  g739(.A(new_n556), .B(KEYINPUT57), .ZN(new_n926));
  INV_X1    g740(.A(new_n899), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n897), .A2(new_n898), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n550), .A2(new_n554), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT117), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n916), .A2(new_n789), .A3(new_n791), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n924), .B1(new_n932), .B2(new_n933), .ZN(G54));
  NAND3_X1  g748(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(new_n638), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n638), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n924), .ZN(G60));
  AND2_X1   g752(.A1(new_n621), .A2(new_n628), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n631), .B(KEYINPUT59), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n940), .B(new_n941), .C1(new_n927), .C2(new_n928), .ZN(new_n942));
  INV_X1    g756(.A(new_n924), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n940), .B1(new_n909), .B2(new_n941), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(G63));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n896), .A2(new_n884), .ZN(new_n952));
  INV_X1    g766(.A(new_n883), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n601), .B(KEYINPUT119), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n948), .B(new_n943), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n660), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n955), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n897), .B2(new_n951), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n948), .B1(new_n960), .B2(new_n943), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n947), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n960), .A2(KEYINPUT121), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(KEYINPUT121), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n924), .A2(new_n947), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n957), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n962), .A2(new_n966), .ZN(G66));
  AOI21_X1  g781(.A(new_n279), .B1(new_n432), .B2(G224), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n902), .A2(new_n845), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(new_n279), .ZN(new_n970));
  INV_X1    g784(.A(new_n243), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(G898), .B2(new_n279), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n970), .B(new_n973), .ZN(G69));
  OAI21_X1  g788(.A(G953), .B1(new_n547), .B2(new_n682), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n775), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n878), .A2(new_n760), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n808), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n777), .B1(new_n788), .B2(new_n800), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n707), .A2(new_n799), .A3(new_n770), .A4(new_n750), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n279), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n279), .A2(G900), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(KEYINPUT125), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n984), .A2(new_n989), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n496), .A2(new_n497), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n988), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n708), .B1(new_n842), .B2(new_n726), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n996), .A2(new_n770), .A3(new_n785), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT123), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(KEYINPUT124), .B1(new_n999), .B2(new_n801), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT124), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n998), .B(new_n1001), .C1(new_n800), .C2(new_n788), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n808), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n716), .A2(new_n978), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT62), .ZN(new_n1005));
  AOI21_X1  g819(.A(G953), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n1006), .A2(new_n993), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n994), .A2(new_n995), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n995), .B1(new_n994), .B2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n976), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n994), .A2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(KEYINPUT126), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n994), .A2(new_n995), .A3(new_n1007), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n975), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1010), .A2(new_n1014), .ZN(G72));
  OR2_X1    g829(.A1(new_n983), .A2(new_n969), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  AND2_X1   g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n943), .B1(new_n1019), .B2(new_n514), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n514), .A2(new_n1018), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n908), .A2(new_n700), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1018), .B1(new_n1023), .B2(new_n969), .ZN(new_n1024));
  AOI211_X1 g838(.A(new_n1020), .B(new_n1022), .C1(new_n700), .C2(new_n1024), .ZN(G57));
endmodule


