//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1214, new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n470), .B2(new_n465), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n468), .B1(new_n471), .B2(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n476), .A2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n465), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n466), .A2(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n464), .A2(new_n487), .A3(new_n465), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n489), .B2(G136), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n473), .A2(new_n475), .A3(G138), .A4(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  OAI211_X1 g069(.A(KEYINPUT70), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n473), .A2(new_n475), .A3(G126), .A4(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  AND4_X1   g076(.A1(G138), .A2(new_n473), .A3(new_n475), .A4(new_n465), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT71), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT4), .B1(new_n493), .B2(KEYINPUT70), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n495), .B(new_n500), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  INV_X1    g095(.A(G88), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n508), .A2(new_n510), .A3(new_n515), .A4(new_n517), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n514), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND3_X1  g100(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n526), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n515), .A2(new_n517), .A3(G51), .A4(G543), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n522), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G168));
  NAND3_X1  g110(.A1(new_n508), .A2(new_n510), .A3(G64), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n511), .A2(new_n518), .A3(G90), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n515), .A2(new_n517), .A3(G52), .A4(G543), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n539), .A2(KEYINPUT72), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n541), .B1(new_n522), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n513), .B1(new_n536), .B2(new_n537), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n542), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n508), .A2(new_n510), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n553), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n554), .A2(G651), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n519), .ZN(new_n557));
  INV_X1    g132(.A(new_n522), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n557), .A2(G43), .B1(G81), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  AND3_X1   g137(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  XNOR2_X1  g142(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n557), .A2(KEYINPUT75), .A3(G53), .A4(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n518), .A2(G53), .A3(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT9), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n573), .B1(new_n571), .B2(new_n568), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n570), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n576), .A2(G65), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n558), .A2(G91), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n575), .A2(new_n581), .A3(new_n582), .ZN(G299));
  INV_X1    g158(.A(G171), .ZN(G301));
  OR2_X1    g159(.A1(new_n531), .A2(new_n534), .ZN(G286));
  NAND2_X1  g160(.A1(new_n557), .A2(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n558), .A2(G87), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  INV_X1    g164(.A(G48), .ZN(new_n590));
  INV_X1    g165(.A(G86), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n519), .A2(new_n590), .B1(new_n591), .B2(new_n522), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n550), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT77), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n592), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n513), .ZN(new_n604));
  XNOR2_X1  g179(.A(KEYINPUT78), .B(G47), .ZN(new_n605));
  INV_X1    g180(.A(G85), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n519), .A2(new_n605), .B1(new_n606), .B2(new_n522), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT79), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n576), .A2(G66), .A3(new_n577), .ZN(new_n612));
  AND2_X1   g187(.A1(G79), .A2(G543), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(new_n513), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n614), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(KEYINPUT79), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n558), .A2(KEYINPUT10), .A3(G92), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT10), .ZN(new_n620));
  INV_X1    g195(.A(G92), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n522), .B2(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n619), .A2(new_n622), .B1(new_n557), .B2(G54), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT80), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n610), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n610), .B1(new_n625), .B2(G868), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n575), .A2(new_n581), .A3(new_n582), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G297));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(G868), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  INV_X1    g208(.A(G868), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n560), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n625), .A2(new_n632), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(new_n634), .ZN(G323));
  XNOR2_X1  g212(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g213(.A1(new_n481), .A2(G123), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n465), .A2(G111), .ZN(new_n640));
  OAI21_X1  g215(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(G135), .B2(new_n489), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT82), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n464), .A2(new_n462), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT13), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2100), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n645), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2435), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2443), .B(G2446), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1341), .B(G1348), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XOR2_X1   g243(.A(G2067), .B(G2678), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT84), .ZN(new_n670));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n670), .A2(new_n672), .ZN(new_n675));
  INV_X1    g250(.A(new_n671), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(KEYINPUT17), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n672), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n676), .B1(new_n675), .B2(KEYINPUT17), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G2096), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n683), .A3(new_n684), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  INV_X1    g266(.A(new_n683), .ZN(new_n692));
  INV_X1    g267(.A(new_n684), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(KEYINPUT85), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n683), .A2(new_n684), .A3(KEYINPUT85), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n695), .A2(new_n688), .A3(new_n696), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n689), .B(new_n690), .C1(new_n691), .C2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n691), .B2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT21), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT86), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1981), .B(G1986), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n704), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n702), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n706), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n707), .A2(new_n711), .ZN(G229));
  NOR2_X1   g287(.A1(G16), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(G288), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G22), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n718), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(G1971), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(G6), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n601), .B2(new_n718), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT32), .B(G1981), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n720), .A2(G1971), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n717), .A2(new_n721), .A3(new_n725), .A4(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n723), .A2(new_n724), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n718), .A2(G24), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n608), .B2(new_n718), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1986), .Z(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G25), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n481), .A2(G119), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n465), .A2(G107), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n489), .B2(G131), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n735), .B1(new_n740), .B2(new_n734), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT35), .B(G1991), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n741), .A2(new_n743), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n733), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n730), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT87), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n730), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n749), .A2(KEYINPUT36), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n734), .A2(G27), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n757), .B(new_n758), .C1(new_n505), .C2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  INV_X1    g335(.A(G2078), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT23), .B1(new_n629), .B2(new_n718), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n718), .A2(G20), .ZN(new_n764));
  MUX2_X1   g339(.A(KEYINPUT23), .B(new_n763), .S(new_n764), .Z(new_n765));
  OAI21_X1  g340(.A(new_n762), .B1(new_n765), .B2(G1956), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n734), .A2(G26), .ZN(new_n767));
  OR2_X1    g342(.A1(G104), .A2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n769));
  INV_X1    g344(.A(new_n481), .ZN(new_n770));
  INV_X1    g345(.A(G128), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n489), .B2(G140), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n767), .B1(new_n773), .B2(new_n734), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n767), .B(new_n774), .S(KEYINPUT28), .Z(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G19), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n561), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT88), .B(G1341), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n766), .B(new_n782), .C1(G1956), .C2(new_n765), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n489), .A2(G139), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n462), .A2(G103), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT25), .Z(new_n786));
  AOI22_X1  g361(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n786), .C1(new_n465), .C2(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G33), .B(new_n788), .S(G29), .Z(new_n789));
  NOR2_X1   g364(.A1(new_n789), .A2(G2072), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n789), .A2(G2072), .ZN(new_n791));
  AOI211_X1 g366(.A(new_n790), .B(new_n791), .C1(G29), .C2(new_n644), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n734), .B1(KEYINPUT24), .B2(G34), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(KEYINPUT24), .B2(G34), .ZN(new_n794));
  INV_X1    g369(.A(G160), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G29), .ZN(new_n796));
  INV_X1    g371(.A(G2084), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(G168), .A2(G16), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G16), .B2(G21), .ZN(new_n800));
  INV_X1    g375(.A(G1966), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G28), .ZN(new_n803));
  AOI21_X1  g378(.A(G29), .B1(new_n803), .B2(KEYINPUT30), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(KEYINPUT30), .B2(new_n803), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT90), .B(KEYINPUT31), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G11), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n802), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n796), .A2(new_n797), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n800), .A2(new_n801), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G5), .A2(G16), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G171), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(G1961), .Z(new_n814));
  NAND4_X1  g389(.A1(new_n792), .A2(new_n798), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n734), .A2(G32), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n462), .A2(G105), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT89), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n481), .A2(G129), .ZN(new_n819));
  NAND3_X1  g394(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT26), .Z(new_n821));
  NAND3_X1  g396(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G141), .B2(new_n489), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n816), .B1(new_n823), .B2(new_n734), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT27), .ZN(new_n825));
  INV_X1    g400(.A(G1996), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n734), .A2(G35), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G162), .B2(new_n734), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT29), .B(G2090), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n815), .A2(new_n827), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(G4), .A2(G16), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n625), .B2(G16), .ZN(new_n834));
  INV_X1    g409(.A(G1348), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n783), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT92), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n756), .A2(new_n839), .ZN(G311));
  XNOR2_X1  g415(.A(new_n837), .B(KEYINPUT92), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n841), .A2(new_n755), .A3(new_n754), .ZN(G150));
  NAND3_X1  g417(.A1(new_n518), .A2(G55), .A3(G543), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n558), .A2(G93), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n513), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n625), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n556), .A2(new_n846), .A3(new_n559), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n846), .B1(new_n556), .B2(new_n559), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n851), .A2(new_n855), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n848), .B1(new_n857), .B2(new_n858), .ZN(G145));
  XNOR2_X1  g434(.A(new_n773), .B(G164), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n788), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(new_n823), .Z(new_n862));
  INV_X1    g437(.A(KEYINPUT96), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n481), .A2(G130), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n465), .A2(G118), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n489), .B2(G142), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n648), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n740), .ZN(new_n870));
  XNOR2_X1  g445(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT93), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n870), .B(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n862), .A2(new_n863), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G162), .B(G160), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n644), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n861), .B(new_n823), .ZN(new_n877));
  INV_X1    g452(.A(new_n872), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n870), .B(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n877), .B1(new_n879), .B2(KEYINPUT96), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n874), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n877), .B(new_n873), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(new_n876), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(G395));
  INV_X1    g463(.A(KEYINPUT99), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n854), .B(KEYINPUT97), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n636), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n618), .A2(G299), .A3(new_n623), .ZN(new_n892));
  AOI21_X1  g467(.A(G299), .B1(new_n618), .B2(new_n623), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n625), .A2(new_n632), .ZN(new_n896));
  INV_X1    g471(.A(new_n890), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n891), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n892), .B2(new_n893), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n624), .A2(new_n629), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n618), .A2(G299), .A3(new_n623), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n891), .B2(new_n898), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n889), .B(KEYINPUT42), .C1(new_n899), .C2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(G166), .B(new_n601), .ZN(new_n909));
  NAND2_X1  g484(.A1(G290), .A2(new_n714), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n608), .A2(G288), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT98), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n912), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT98), .B1(new_n910), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n913), .B1(new_n916), .B2(new_n909), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(KEYINPUT99), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n891), .A2(new_n895), .A3(new_n898), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n891), .A2(new_n898), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n921), .B(new_n922), .C1(new_n923), .C2(new_n906), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n908), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n920), .B1(new_n908), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n846), .A2(new_n634), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT101), .B1(G171), .B2(G286), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n933));
  NAND4_X1  g508(.A1(G168), .A2(new_n933), .A3(new_n542), .A4(new_n547), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(G171), .A2(G286), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(KEYINPUT102), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(G171), .B2(G286), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n854), .B(new_n935), .C1(new_n937), .C2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n936), .B(KEYINPUT102), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n854), .B1(new_n943), .B2(new_n935), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n941), .B(new_n854), .C1(new_n943), .C2(new_n935), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n937), .A2(new_n939), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n932), .A2(new_n934), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n855), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n940), .ZN(new_n952));
  OAI211_X1 g527(.A(KEYINPUT103), .B(new_n855), .C1(new_n948), .C2(new_n949), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n894), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n905), .A2(new_n947), .B1(new_n954), .B2(KEYINPUT106), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n954), .A2(KEYINPUT106), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n917), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n895), .B1(new_n945), .B2(new_n946), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n905), .A2(new_n952), .A3(new_n953), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n917), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n882), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT43), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n905), .A2(new_n952), .A3(new_n953), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n942), .A2(new_n944), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n950), .A2(new_n941), .A3(new_n940), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n894), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n918), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n882), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n917), .B1(new_n958), .B2(new_n959), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT105), .B1(new_n970), .B2(G37), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT100), .B(KEYINPUT43), .Z(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n969), .A2(new_n971), .A3(new_n960), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n931), .B1(new_n962), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n957), .A2(new_n961), .A3(new_n972), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n969), .A2(new_n971), .A3(new_n960), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n975), .B1(new_n978), .B2(new_n931), .ZN(G397));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n464), .A2(KEYINPUT71), .A3(G138), .A4(new_n465), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n504), .B1(KEYINPUT70), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n495), .A2(new_n500), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n468), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n470), .A2(new_n469), .A3(new_n465), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT67), .B1(new_n478), .B2(G2105), .ZN(new_n989));
  OAI211_X1 g564(.A(G40), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n986), .A2(G1996), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT107), .B1(new_n991), .B2(new_n823), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n986), .A2(new_n990), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n773), .B(G2067), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n826), .B2(new_n823), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n740), .B(new_n743), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n993), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(KEYINPUT107), .A3(new_n823), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n608), .B(G1986), .Z(new_n1001));
  AOI21_X1  g576(.A(new_n1000), .B1(new_n993), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT109), .B(G8), .Z(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G40), .ZN(new_n1005));
  AOI211_X1 g580(.A(new_n1005), .B(new_n468), .C1(new_n471), .C2(new_n479), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n495), .A2(new_n500), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT70), .B1(new_n493), .B2(new_n494), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(KEYINPUT4), .C1(KEYINPUT70), .C2(new_n493), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1384), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1004), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n601), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(G1981), .B1(new_n597), .B2(new_n592), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(KEYINPUT110), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(KEYINPUT110), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1014), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1011), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n714), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1013), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1011), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  XOR2_X1   g600(.A(new_n1025), .B(KEYINPUT55), .Z(new_n1026));
  NAND3_X1  g601(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT108), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n986), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n984), .A2(KEYINPUT108), .A3(new_n985), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1006), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1971), .ZN(new_n1032));
  AND2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n505), .A2(new_n1035), .A3(new_n980), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1006), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(G2090), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1026), .C1(new_n1033), .C2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n714), .A2(G1976), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n1021), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1011), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1011), .A2(new_n1040), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1020), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1024), .B1(new_n1039), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1045), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1047), .A2(new_n1039), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT113), .B(G2084), .Z(new_n1049));
  AND4_X1   g624(.A1(new_n1006), .A2(new_n1034), .A3(new_n1036), .A4(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n505), .B2(new_n980), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT112), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1027), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1010), .A2(KEYINPUT112), .A3(KEYINPUT45), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1006), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1055), .B2(new_n801), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(G168), .A3(new_n1003), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT63), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1061));
  INV_X1    g636(.A(G8), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1048), .B(new_n1060), .C1(new_n1063), .C2(new_n1026), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1035), .B1(new_n505), .B2(new_n980), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT111), .B1(new_n1065), .B2(new_n990), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1006), .B(new_n1067), .C1(new_n1010), .C2(new_n1035), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1036), .A3(new_n1068), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1069), .A2(G2090), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1004), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1047), .B(new_n1039), .C1(new_n1026), .C2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1059), .B1(new_n1073), .B2(new_n1058), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1046), .B1(new_n1064), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(G2078), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n987), .A2(G40), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(G2105), .B2(new_n478), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n986), .A2(new_n1079), .A3(new_n1027), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT122), .B(G1961), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1037), .A2(KEYINPUT123), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT123), .B1(new_n1037), .B2(new_n1081), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1080), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1029), .A2(new_n761), .A3(new_n1006), .A4(new_n1030), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1086), .A2(new_n1076), .ZN(new_n1087));
  OAI21_X1  g662(.A(G171), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1076), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1037), .A2(new_n1081), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT112), .B1(new_n1010), .B2(KEYINPUT45), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n990), .B1(new_n1091), .B2(new_n1027), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(new_n1054), .A3(new_n1077), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1089), .A2(G301), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1088), .A2(KEYINPUT54), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1090), .ZN(new_n1096));
  OAI21_X1  g671(.A(G171), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1084), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1082), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1099), .A2(G301), .A3(new_n1089), .A4(new_n1080), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT54), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1095), .A2(new_n1073), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G168), .A2(new_n1004), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1966), .B1(new_n1092), .B2(new_n1054), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1003), .B1(new_n1106), .B2(new_n1050), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1103), .A2(KEYINPUT51), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1105), .A2(KEYINPUT51), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1056), .A2(new_n1104), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT121), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1110), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  OAI21_X1  g689(.A(G8), .B1(new_n1106), .B2(new_n1050), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n1104), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1108), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1117), .B1(new_n1057), .B2(new_n1003), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1112), .B(new_n1113), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1111), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1102), .A2(new_n1120), .ZN(new_n1121));
  XOR2_X1   g696(.A(KEYINPUT114), .B(G1956), .Z(new_n1122));
  NAND2_X1  g697(.A1(new_n1069), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n629), .B(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT56), .B(G2072), .Z(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT116), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1029), .A2(new_n1006), .A3(new_n1030), .A4(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1037), .A2(new_n835), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1006), .A2(new_n1010), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(G2067), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n624), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1123), .A2(new_n1128), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1125), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT117), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1135), .A2(new_n1141), .A3(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1138), .A2(KEYINPUT61), .A3(new_n1129), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT61), .B1(new_n1138), .B2(new_n1129), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n624), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1130), .A2(new_n1133), .A3(KEYINPUT60), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1130), .A2(new_n1133), .A3(KEYINPUT60), .A4(new_n624), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1144), .A2(new_n1145), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT58), .B(G1341), .Z(new_n1155));
  AOI21_X1  g730(.A(new_n1154), .B1(new_n1131), .B2(new_n1155), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1154), .B(new_n1155), .C1(new_n984), .C2(new_n990), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1029), .A2(new_n826), .A3(new_n1006), .A4(new_n1030), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT120), .B1(new_n1161), .B2(new_n561), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n1163));
  AOI211_X1 g738(.A(new_n1163), .B(new_n560), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT119), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1162), .A2(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1161), .A2(new_n561), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1163), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1161), .A2(KEYINPUT120), .A3(new_n561), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1143), .B1(new_n1153), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1075), .B1(new_n1121), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1111), .A2(new_n1176), .A3(new_n1119), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1073), .A2(new_n1097), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1176), .B1(new_n1111), .B2(new_n1119), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1002), .B1(new_n1175), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n773), .A2(new_n776), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n996), .A2(new_n999), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n740), .A2(new_n743), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n993), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1186), .A2(KEYINPUT124), .A3(new_n993), .ZN(new_n1190));
  NOR4_X1   g765(.A1(new_n986), .A2(G1986), .A3(G290), .A4(new_n990), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT48), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n1000), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n994), .A2(new_n823), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT125), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT46), .ZN(new_n1196));
  AOI22_X1  g771(.A1(new_n1194), .A2(new_n993), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n991), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n991), .A2(KEYINPUT125), .A3(KEYINPUT46), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  XOR2_X1   g776(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1202));
  XNOR2_X1  g777(.A(new_n1201), .B(new_n1202), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1189), .A2(new_n1190), .A3(new_n1193), .A4(new_n1203), .ZN(new_n1204));
  XNOR2_X1  g779(.A(new_n1204), .B(KEYINPUT127), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1182), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(G319), .ZN(new_n1208));
  NOR2_X1   g782(.A1(G227), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n667), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n707), .B2(new_n711), .ZN(new_n1211));
  OAI21_X1  g785(.A(new_n1211), .B1(new_n885), .B2(new_n883), .ZN(new_n1212));
  NOR2_X1   g786(.A1(new_n1212), .A2(new_n978), .ZN(G308));
  INV_X1    g787(.A(new_n886), .ZN(new_n1214));
  AND2_X1   g788(.A1(new_n977), .A2(new_n972), .ZN(new_n1215));
  OAI211_X1 g789(.A(new_n1214), .B(new_n1211), .C1(new_n1215), .C2(new_n976), .ZN(G225));
endmodule


