//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  OR2_X1    g032(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n458), .A2(KEYINPUT3), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n460), .A2(new_n462), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n462), .A2(new_n465), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n471), .A2(KEYINPUT67), .A3(new_n460), .A4(new_n467), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n464), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n458), .B2(new_n459), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G2105), .B1(G101), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT68), .Z(G160));
  NAND4_X1  g058(.A1(new_n460), .A2(G2105), .A3(new_n462), .A4(new_n465), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n471), .A2(KEYINPUT69), .A3(G2105), .A4(new_n460), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT70), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G112), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n459), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n494), .A2(new_n495), .A3(new_n464), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n462), .A2(new_n465), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n496), .A2(new_n497), .A3(G2105), .ZN(new_n498));
  AND2_X1   g073(.A1(new_n498), .A2(G136), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n490), .A2(new_n493), .A3(new_n499), .ZN(G162));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G126), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n484), .B2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G138), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n508), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(new_n513), .B2(new_n477), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n466), .A2(G138), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT3), .B(G2104), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n510), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n460), .A2(new_n462), .A3(new_n465), .A4(new_n508), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT4), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n506), .B1(new_n521), .B2(new_n523), .ZN(G164));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT5), .B(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n525), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G651), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n531), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  XNOR2_X1  g111(.A(KEYINPUT73), .B(G89), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n527), .A2(new_n537), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n539), .A2(new_n543), .ZN(G168));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n527), .A2(new_n545), .B1(new_n529), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n533), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n547), .A2(new_n549), .ZN(G171));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  INV_X1    g126(.A(G43), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n527), .A2(new_n551), .B1(new_n529), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n533), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  XOR2_X1   g136(.A(KEYINPUT75), .B(G65), .Z(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(new_n526), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n533), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n526), .A2(new_n525), .A3(G91), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n568), .B1(KEYINPUT74), .B2(KEYINPUT9), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT74), .B(KEYINPUT9), .Z(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n567), .A2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  OAI21_X1  g149(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI221_X1 g152(.A(new_n575), .B1(new_n529), .B2(new_n576), .C1(new_n577), .C2(new_n527), .ZN(G288));
  AOI21_X1  g153(.A(KEYINPUT76), .B1(new_n526), .B2(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(G73), .B2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n526), .A2(KEYINPUT76), .A3(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n533), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  INV_X1    g158(.A(G48), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n527), .A2(new_n583), .B1(new_n529), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n527), .A2(new_n588), .B1(new_n529), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n533), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n526), .A2(new_n525), .A3(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT10), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n526), .A2(G66), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n533), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n529), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(G54), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n595), .B1(new_n604), .B2(G868), .ZN(G321));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  XNOR2_X1  g184(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  INV_X1    g187(.A(new_n556), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n603), .A2(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(new_n614), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT78), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n480), .A2(new_n519), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(KEYINPUT79), .B2(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(KEYINPUT79), .A2(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n488), .A2(G123), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(KEYINPUT80), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n627), .A2(KEYINPUT80), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n498), .A2(G135), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n622), .A2(KEYINPUT79), .A3(G2100), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(G2096), .ZN(new_n635));
  NAND4_X1  g210(.A1(new_n625), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT81), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n641), .B(new_n647), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(G14), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT82), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n656), .B(KEYINPUT17), .Z(new_n659));
  INV_X1    g234(.A(new_n657), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n654), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n654), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n657), .A2(new_n654), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT83), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(new_n678), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n681), .B(new_n682), .Z(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT84), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  NOR2_X1   g264(.A1(G29), .A2(G35), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G162), .B2(G29), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT29), .B(G2090), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n604), .A2(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G4), .B2(G16), .ZN(new_n695));
  INV_X1    g270(.A(G1348), .ZN(new_n696));
  NAND2_X1  g271(.A1(G168), .A2(G16), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(KEYINPUT93), .C1(G16), .C2(G21), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(KEYINPUT93), .B2(new_n697), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n695), .A2(new_n696), .B1(new_n699), .B2(G1966), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n696), .B2(new_n695), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n699), .A2(G1966), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT95), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G20), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT23), .Z(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G299), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1956), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT31), .B(G11), .Z(new_n712));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G28), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n713), .B2(G28), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(new_n716), .ZN(new_n719));
  NOR2_X1   g294(.A1(G5), .A2(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT96), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(KEYINPUT96), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n721), .B(new_n722), .C1(G301), .C2(new_n706), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n712), .B(new_n719), .C1(new_n724), .C2(G1961), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n724), .A2(G1961), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G19), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n556), .B2(G16), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(G1341), .Z(new_n729));
  INV_X1    g304(.A(new_n632), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n725), .A2(new_n726), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  NOR4_X1   g307(.A1(new_n701), .A2(new_n704), .A3(new_n711), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G160), .A2(G29), .ZN(new_n734));
  AND2_X1   g309(.A1(KEYINPUT24), .A2(G34), .ZN(new_n735));
  NOR2_X1   g310(.A1(KEYINPUT24), .A2(G34), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n715), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT92), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2084), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n715), .A2(G33), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n498), .A2(G139), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n519), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(new_n466), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT25), .Z(new_n746));
  NAND3_X1  g321(.A1(new_n742), .A2(new_n744), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(new_n715), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT91), .ZN(new_n750));
  INV_X1    g325(.A(G2072), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n715), .A2(G32), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n486), .A2(G129), .A3(new_n487), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n480), .A2(G105), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n471), .A2(new_n466), .A3(new_n460), .ZN(new_n759));
  INV_X1    g334(.A(G141), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n752), .B1(new_n763), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n750), .A2(new_n751), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(G27), .A2(G29), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G164), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2078), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n715), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT28), .Z(new_n771));
  OAI21_X1  g346(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n772));
  INV_X1    g347(.A(G116), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G2105), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n498), .B2(G140), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n486), .A2(new_n487), .ZN(new_n776));
  INV_X1    g351(.A(G128), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT90), .B(G2067), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n769), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n766), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n764), .A2(new_n765), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n779), .A2(new_n780), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n750), .A2(new_n751), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n782), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n693), .A2(new_n733), .A3(new_n740), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n706), .A2(G22), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n706), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n706), .A2(G6), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n586), .B2(new_n706), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT88), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT32), .B(G1981), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n795), .A2(new_n797), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n706), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(G288), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n706), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT33), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1976), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n792), .A2(new_n798), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT87), .B(KEYINPUT34), .Z(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n486), .A2(G119), .A3(new_n487), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(G107), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n498), .B2(G131), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n809), .A2(new_n813), .A3(KEYINPUT85), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(KEYINPUT85), .B1(new_n809), .B2(new_n813), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G29), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G25), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  AND2_X1   g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NOR2_X1   g397(.A1(G16), .A2(G24), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n593), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT86), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1986), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n807), .A2(new_n808), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n787), .B1(new_n829), .B2(new_n830), .ZN(G311));
  XNOR2_X1  g406(.A(G311), .B(KEYINPUT97), .ZN(G150));
  NAND2_X1  g407(.A1(new_n604), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n526), .A2(new_n525), .A3(G93), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT98), .B(G55), .Z(new_n837));
  OAI221_X1 g412(.A(new_n835), .B1(new_n533), .B2(new_n836), .C1(new_n529), .C2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n613), .B(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n834), .B(new_n839), .Z(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n841), .A2(new_n842), .A3(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n838), .A2(G860), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(G162), .B(G160), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n730), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n775), .B1(new_n777), .B2(new_n776), .C1(new_n753), .C2(new_n761), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n754), .A2(new_n778), .A3(new_n762), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n523), .A2(new_n514), .A3(new_n520), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n496), .A2(new_n497), .A3(new_n466), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n503), .B1(new_n854), .B2(G126), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT99), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n858));
  NAND2_X1  g433(.A1(G164), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n850), .A2(new_n851), .B1(new_n857), .B2(new_n859), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n861), .A2(new_n747), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT100), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(new_n860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(new_n850), .A3(new_n851), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n852), .A2(new_n860), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n748), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n863), .B1(new_n870), .B2(KEYINPUT101), .ZN(new_n871));
  INV_X1    g446(.A(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n466), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI22_X1  g449(.A1(new_n759), .A2(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G130), .ZN(new_n876));
  OR3_X1    g451(.A1(new_n776), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT102), .B1(new_n776), .B2(new_n876), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n816), .ZN(new_n880));
  INV_X1    g455(.A(new_n621), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n814), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n621), .B1(new_n815), .B2(new_n816), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n879), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n883), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n861), .A2(KEYINPUT100), .A3(new_n862), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n747), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT101), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n871), .A2(new_n889), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n889), .B1(new_n871), .B2(new_n894), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n849), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n871), .A2(new_n889), .A3(new_n894), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n871), .A2(new_n894), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n848), .B(new_n898), .C1(new_n899), .C2(new_n887), .ZN(new_n900));
  INV_X1    g475(.A(G37), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT104), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n897), .A2(new_n900), .A3(new_n904), .A4(new_n901), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n903), .A2(KEYINPUT40), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT40), .B1(new_n903), .B2(new_n905), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n907), .ZN(G395));
  NAND2_X1  g483(.A1(new_n838), .A2(new_n614), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n593), .B(G288), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(G303), .B2(G305), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G303), .B2(G305), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT106), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT42), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n839), .B(new_n616), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n608), .B(new_n603), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n920), .B(KEYINPUT41), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n919), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n918), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n909), .B1(new_n924), .B2(new_n614), .ZN(G295));
  OAI21_X1  g500(.A(new_n909), .B1(new_n924), .B2(new_n614), .ZN(G331));
  XNOR2_X1  g501(.A(new_n839), .B(G301), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(G168), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(new_n922), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n920), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G37), .B1(new_n931), .B2(new_n916), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n929), .A2(new_n915), .A3(new_n930), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n936), .A3(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(KEYINPUT107), .B2(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n935), .A2(new_n937), .A3(new_n940), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(G397));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n865), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n473), .A2(G40), .A3(new_n481), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n473), .A2(G40), .A3(new_n481), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(KEYINPUT108), .A3(new_n948), .A4(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n778), .B(G2067), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT109), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n763), .B(G1996), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n957), .A2(new_n959), .B1(new_n954), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n817), .A2(new_n820), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n817), .A2(new_n820), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n593), .B(G1986), .Z(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n954), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1966), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n853), .B2(new_n855), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n969), .B(new_n952), .C1(new_n970), .C2(KEYINPUT45), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n948), .B1(G164), .B2(G1384), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n969), .B1(new_n974), .B2(new_n952), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n968), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(G2084), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n950), .B1(new_n970), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n856), .A2(new_n946), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT110), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n970), .A2(new_n982), .A3(new_n978), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n977), .B(new_n979), .C1(new_n981), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n976), .A2(KEYINPUT117), .A3(new_n984), .ZN(new_n988));
  AOI21_X1  g563(.A(G286), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(KEYINPUT51), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  NOR2_X1   g566(.A1(G168), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n992), .A2(KEYINPUT51), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n991), .B1(new_n976), .B2(new_n984), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT119), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI211_X1 g571(.A(KEYINPUT119), .B(new_n991), .C1(new_n976), .C2(new_n984), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n989), .A2(new_n990), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT62), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n987), .A2(new_n992), .A3(new_n988), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n987), .A2(KEYINPUT118), .A3(new_n988), .A4(new_n992), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT124), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n857), .A2(new_n859), .A3(KEYINPUT45), .A4(new_n946), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n950), .B1(new_n980), .B2(new_n948), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n790), .ZN(new_n1009));
  OAI21_X1  g584(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n979), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(G2090), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(G303), .A2(G8), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n952), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1010), .A2(new_n982), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n980), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2090), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n991), .B1(new_n1022), .B2(new_n1009), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1015), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G305), .A2(G1981), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n582), .A2(G1981), .A3(new_n585), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n980), .A2(new_n950), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n991), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1027), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n801), .A2(G1976), .ZN(new_n1035));
  INV_X1    g610(.A(G1976), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1034), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1016), .A2(new_n1025), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n952), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT111), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(G2078), .ZN(new_n1046));
  AND4_X1   g621(.A1(new_n1044), .A2(new_n971), .A3(new_n972), .A4(new_n1046), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT120), .B(G1961), .Z(new_n1048));
  NAND2_X1  g623(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1049), .B2(new_n979), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT121), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1044), .A2(new_n971), .A3(new_n972), .A4(new_n1046), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(new_n1053), .C1(new_n1020), .C2(new_n1048), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1008), .A2(G2078), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1056));
  AOI22_X1  g631(.A1(new_n1051), .A2(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1042), .A2(G301), .A3(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1004), .A2(new_n1005), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1005), .B1(new_n1004), .B2(new_n1058), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n999), .B1(new_n1061), .B2(new_n998), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT113), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1065), .A2(KEYINPUT63), .A3(new_n1025), .A4(new_n1041), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n994), .A2(G168), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1064), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1065), .A2(KEYINPUT63), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1067), .B(KEYINPUT112), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1025), .A2(new_n1041), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(KEYINPUT113), .A4(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1069), .B2(new_n1042), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1070), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1025), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1034), .A2(new_n1036), .A3(new_n801), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1027), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1078), .A2(new_n1041), .B1(new_n1080), .B2(new_n1032), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n949), .A2(new_n952), .A3(new_n1006), .A4(new_n1046), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1050), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(G301), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1085), .B1(new_n1057), .B2(G301), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1086), .A2(KEYINPUT123), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT123), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT114), .B1(new_n565), .B2(new_n566), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n571), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n565), .A2(KEYINPUT114), .A3(new_n566), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n608), .A2(KEYINPUT57), .ZN(new_n1098));
  OAI211_X1 g673(.A(KEYINPUT115), .B(new_n1091), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1011), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1006), .A2(new_n1007), .A3(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1100), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT116), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT61), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT116), .B(new_n1109), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1031), .ZN(new_n1112));
  OAI221_X1 g687(.A(KEYINPUT60), .B1(G2067), .B2(new_n1112), .C1(new_n1020), .C2(G1348), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT60), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1348), .B1(new_n1049), .B2(new_n979), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1112), .A2(G2067), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1113), .A2(new_n1117), .A3(new_n604), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT58), .B(G1341), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1008), .A2(G1996), .B1(new_n1031), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(KEYINPUT59), .A3(new_n556), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT60), .A3(new_n603), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n556), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1118), .A2(new_n1121), .A3(new_n1123), .A4(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1122), .A2(new_n603), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(new_n1106), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1111), .A2(new_n1127), .B1(new_n1129), .B2(new_n1105), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1057), .A2(G301), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1087), .B1(new_n1133), .B2(G171), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1042), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1077), .B(new_n1081), .C1(new_n1090), .C2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n967), .B1(new_n1063), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n955), .A2(new_n763), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n954), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(KEYINPUT125), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n951), .A2(new_n953), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1142), .A2(G1996), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1143), .A2(KEYINPUT46), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1140), .A2(KEYINPUT125), .B1(new_n1143), .B2(KEYINPUT46), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1142), .A2(G1986), .A3(G290), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT48), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n1149), .A2(new_n1150), .B1(new_n965), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n961), .A2(new_n962), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n778), .A2(G2067), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1142), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1138), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g733(.A1(new_n903), .A2(new_n905), .ZN(new_n1160));
  OAI21_X1  g734(.A(G319), .B1(new_n651), .B2(new_n652), .ZN(new_n1161));
  NOR2_X1   g735(.A1(G227), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n688), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g737(.A(new_n1163), .B(KEYINPUT127), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n1160), .A2(new_n938), .A3(new_n1164), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


