

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783;

  NOR2_X1 U369 ( .A1(n715), .A2(n378), .ZN(n375) );
  XNOR2_X1 U370 ( .A(n616), .B(n346), .ZN(n379) );
  XNOR2_X1 U371 ( .A(n380), .B(KEYINPUT90), .ZN(n346) );
  XNOR2_X1 U372 ( .A(n596), .B(KEYINPUT101), .ZN(n698) );
  NAND2_X1 U373 ( .A1(n412), .A2(n410), .ZN(n606) );
  OR2_X1 U374 ( .A1(n583), .A2(n639), .ZN(n575) );
  XNOR2_X1 U375 ( .A(n528), .B(n527), .ZN(n563) );
  OR2_X1 U376 ( .A1(n600), .A2(n601), .ZN(n430) );
  XNOR2_X1 U377 ( .A(n548), .B(n547), .ZN(n772) );
  XNOR2_X1 U378 ( .A(G116), .B(G122), .ZN(n513) );
  XNOR2_X1 U379 ( .A(G104), .B(G122), .ZN(n439) );
  NAND2_X2 U380 ( .A1(n372), .A2(n371), .ZN(n445) );
  XNOR2_X2 U381 ( .A(n529), .B(n530), .ZN(n773) );
  XNOR2_X2 U382 ( .A(n510), .B(n509), .ZN(n529) );
  XNOR2_X1 U383 ( .A(n725), .B(KEYINPUT86), .ZN(n627) );
  INV_X2 U384 ( .A(G125), .ZN(n460) );
  XNOR2_X1 U385 ( .A(G119), .B(G128), .ZN(n549) );
  XNOR2_X1 U386 ( .A(KEYINPUT16), .B(G122), .ZN(n488) );
  NOR2_X1 U387 ( .A1(n386), .A2(n751), .ZN(n588) );
  XNOR2_X1 U388 ( .A(n641), .B(n640), .ZN(n782) );
  XNOR2_X2 U389 ( .A(n449), .B(n352), .ZN(n614) );
  BUF_X1 U390 ( .A(n511), .Z(n777) );
  NOR2_X1 U391 ( .A1(n608), .A2(n607), .ZN(n609) );
  AND2_X1 U392 ( .A1(n414), .A2(n413), .ZN(n412) );
  NAND2_X1 U393 ( .A1(n422), .A2(n442), .ZN(n596) );
  XNOR2_X1 U394 ( .A(n645), .B(n454), .ZN(n783) );
  AND2_X1 U395 ( .A1(n379), .A2(n732), .ZN(n715) );
  NAND2_X1 U396 ( .A1(n408), .A2(n407), .ZN(n635) );
  XNOR2_X1 U397 ( .A(n638), .B(KEYINPUT38), .ZN(n720) );
  NAND2_X1 U398 ( .A1(n434), .A2(n431), .ZN(n713) );
  NAND2_X1 U399 ( .A1(n430), .A2(n435), .ZN(n434) );
  XNOR2_X1 U400 ( .A(n673), .B(n676), .ZN(n677) );
  OR2_X1 U401 ( .A1(n666), .A2(G902), .ZN(n389) );
  INV_X4 U402 ( .A(G953), .ZN(n511) );
  XNOR2_X1 U403 ( .A(G104), .B(G107), .ZN(n478) );
  AND2_X1 U404 ( .A1(n582), .A2(n731), .ZN(n347) );
  INV_X1 U405 ( .A(n638), .ZN(n348) );
  AND2_X1 U406 ( .A1(n620), .A2(n577), .ZN(n615) );
  XNOR2_X2 U407 ( .A(n613), .B(n612), .ZN(n758) );
  NOR2_X1 U408 ( .A1(n397), .A2(n394), .ZN(n381) );
  NAND2_X1 U409 ( .A1(n393), .A2(n452), .ZN(n392) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n537) );
  INV_X1 U411 ( .A(G469), .ZN(n427) );
  OR2_X1 U412 ( .A1(n693), .A2(G902), .ZN(n428) );
  XNOR2_X1 U413 ( .A(n459), .B(n505), .ZN(n548) );
  XOR2_X1 U414 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n505) );
  XNOR2_X1 U415 ( .A(n504), .B(G140), .ZN(n459) );
  OR2_X1 U416 ( .A1(n712), .A2(n419), .ZN(n416) );
  INV_X1 U417 ( .A(KEYINPUT68), .ZN(n461) );
  NAND2_X1 U418 ( .A1(n630), .A2(n629), .ZN(n401) );
  OR2_X1 U419 ( .A1(n783), .A2(KEYINPUT46), .ZN(n452) );
  AND2_X1 U420 ( .A1(n698), .A2(n355), .ZN(n358) );
  NAND2_X1 U421 ( .A1(n627), .A2(KEYINPUT108), .ZN(n417) );
  XNOR2_X1 U422 ( .A(KEYINPUT4), .B(G131), .ZN(n530) );
  XNOR2_X1 U423 ( .A(n593), .B(n533), .ZN(n582) );
  AND2_X1 U424 ( .A1(n441), .A2(n597), .ZN(n440) );
  NAND2_X1 U425 ( .A1(n594), .A2(n595), .ZN(n441) );
  NAND2_X1 U426 ( .A1(n444), .A2(KEYINPUT99), .ZN(n443) );
  XNOR2_X1 U427 ( .A(n354), .B(n503), .ZN(n436) );
  AND2_X1 U428 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U429 ( .A1(n715), .A2(n378), .ZN(n373) );
  AND2_X1 U430 ( .A1(n604), .A2(n471), .ZN(n611) );
  INV_X1 U431 ( .A(KEYINPUT112), .ZN(n426) );
  XNOR2_X1 U432 ( .A(n458), .B(n457), .ZN(n750) );
  INV_X1 U433 ( .A(KEYINPUT41), .ZN(n457) );
  NOR2_X1 U434 ( .A1(n723), .A2(n456), .ZN(n455) );
  XNOR2_X1 U435 ( .A(n405), .B(n468), .ZN(n647) );
  NOR2_X1 U436 ( .A1(n635), .A2(n406), .ZN(n405) );
  NAND2_X1 U437 ( .A1(n720), .A2(n446), .ZN(n406) );
  NAND2_X1 U438 ( .A1(n567), .A2(KEYINPUT32), .ZN(n413) );
  XOR2_X1 U439 ( .A(KEYINPUT93), .B(KEYINPUT0), .Z(n467) );
  AND2_X1 U440 ( .A1(n623), .A2(n631), .ZN(n643) );
  XNOR2_X1 U441 ( .A(KEYINPUT28), .B(KEYINPUT113), .ZN(n621) );
  NAND2_X1 U442 ( .A1(n398), .A2(n400), .ZN(n397) );
  NAND2_X1 U443 ( .A1(n401), .A2(KEYINPUT76), .ZN(n400) );
  AND2_X1 U444 ( .A1(n403), .A2(n402), .ZN(n399) );
  INV_X1 U445 ( .A(KEYINPUT108), .ZN(n419) );
  INV_X1 U446 ( .A(G237), .ZN(n489) );
  XOR2_X1 U447 ( .A(G137), .B(KEYINPUT100), .Z(n539) );
  XNOR2_X1 U448 ( .A(n439), .B(n438), .ZN(n437) );
  XNOR2_X1 U449 ( .A(KEYINPUT102), .B(KEYINPUT11), .ZN(n438) );
  XOR2_X1 U450 ( .A(G137), .B(KEYINPUT71), .Z(n547) );
  XNOR2_X1 U451 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n475) );
  XNOR2_X1 U452 ( .A(G902), .B(KEYINPUT15), .ZN(n654) );
  NAND2_X1 U453 ( .A1(G234), .A2(G237), .ZN(n496) );
  INV_X1 U454 ( .A(KEYINPUT48), .ZN(n378) );
  XNOR2_X1 U455 ( .A(n463), .B(n560), .ZN(n581) );
  XNOR2_X1 U456 ( .A(KEYINPUT94), .B(KEYINPUT3), .ZN(n486) );
  XOR2_X1 U457 ( .A(KEYINPUT24), .B(KEYINPUT88), .Z(n552) );
  XOR2_X1 U458 ( .A(KEYINPUT23), .B(G110), .Z(n550) );
  XNOR2_X1 U459 ( .A(n421), .B(n420), .ZN(n551) );
  INV_X1 U460 ( .A(KEYINPUT8), .ZN(n420) );
  NAND2_X1 U461 ( .A1(n511), .A2(G234), .ZN(n421) );
  XNOR2_X1 U462 ( .A(KEYINPUT9), .B(KEYINPUT105), .ZN(n515) );
  XOR2_X1 U463 ( .A(KEYINPUT103), .B(KEYINPUT7), .Z(n516) );
  XOR2_X1 U464 ( .A(KEYINPUT104), .B(G107), .Z(n514) );
  INV_X1 U465 ( .A(G134), .ZN(n509) );
  XNOR2_X1 U466 ( .A(n773), .B(G146), .ZN(n536) );
  XNOR2_X1 U467 ( .A(n713), .B(KEYINPUT107), .ZN(n646) );
  AND2_X1 U468 ( .A1(n631), .A2(n731), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n633), .B(n409), .ZN(n408) );
  INV_X1 U470 ( .A(KEYINPUT30), .ZN(n409) );
  INV_X1 U471 ( .A(KEYINPUT106), .ZN(n435) );
  INV_X1 U472 ( .A(G475), .ZN(n507) );
  AND2_X1 U473 ( .A1(n415), .A2(n440), .ZN(n422) );
  XOR2_X1 U474 ( .A(KEYINPUT62), .B(n658), .Z(n659) );
  XNOR2_X1 U475 ( .A(n465), .B(n390), .ZN(n778) );
  INV_X1 U476 ( .A(n776), .ZN(n390) );
  XNOR2_X1 U477 ( .A(n541), .B(n488), .ZN(n766) );
  XNOR2_X1 U478 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U479 ( .A(n536), .B(n383), .ZN(n693) );
  XNOR2_X1 U480 ( .A(n384), .B(n532), .ZN(n383) );
  XNOR2_X1 U481 ( .A(n531), .B(n385), .ZN(n384) );
  XNOR2_X1 U482 ( .A(n429), .B(KEYINPUT80), .ZN(n385) );
  NOR2_X1 U483 ( .A1(n777), .A2(G952), .ZN(n696) );
  INV_X1 U484 ( .A(KEYINPUT79), .ZN(n650) );
  NAND2_X1 U485 ( .A1(n580), .A2(n638), .ZN(n649) );
  XNOR2_X1 U486 ( .A(n579), .B(n425), .ZN(n580) );
  XNOR2_X1 U487 ( .A(n426), .B(KEYINPUT43), .ZN(n425) );
  INV_X1 U488 ( .A(KEYINPUT42), .ZN(n454) );
  XNOR2_X1 U489 ( .A(KEYINPUT40), .B(KEYINPUT114), .ZN(n640) );
  INV_X1 U490 ( .A(KEYINPUT36), .ZN(n380) );
  NOR2_X1 U491 ( .A1(n567), .A2(KEYINPUT32), .ZN(n411) );
  INV_X1 U492 ( .A(KEYINPUT31), .ZN(n356) );
  AND2_X1 U493 ( .A1(n649), .A2(n781), .ZN(n349) );
  AND2_X1 U494 ( .A1(n349), .A2(KEYINPUT2), .ZN(n350) );
  AND2_X1 U495 ( .A1(n643), .A2(n370), .ZN(n351) );
  XOR2_X1 U496 ( .A(n492), .B(n491), .Z(n352) );
  XOR2_X1 U497 ( .A(n508), .B(n507), .Z(n353) );
  BUF_X1 U498 ( .A(n582), .Z(n732) );
  AND2_X1 U499 ( .A1(G214), .A2(n537), .ZN(n354) );
  AND2_X1 U500 ( .A1(n602), .A2(n419), .ZN(n355) );
  INV_X1 U501 ( .A(KEYINPUT76), .ZN(n402) );
  XNOR2_X1 U502 ( .A(n586), .B(n585), .ZN(n751) );
  XNOR2_X1 U503 ( .A(n632), .B(KEYINPUT6), .ZN(n583) );
  XNOR2_X1 U504 ( .A(n357), .B(n356), .ZN(n712) );
  AND2_X1 U505 ( .A1(n599), .A2(n740), .ZN(n357) );
  XNOR2_X1 U506 ( .A(n495), .B(n494), .ZN(n387) );
  NAND2_X1 U507 ( .A1(n563), .A2(n583), .ZN(n568) );
  NOR2_X1 U508 ( .A1(n358), .A2(n359), .ZN(n368) );
  NAND2_X1 U509 ( .A1(n418), .A2(n417), .ZN(n359) );
  XNOR2_X1 U510 ( .A(n592), .B(KEYINPUT35), .ZN(n360) );
  BUF_X1 U511 ( .A(n632), .Z(n738) );
  AND2_X1 U512 ( .A1(n729), .A2(n632), .ZN(n619) );
  AND2_X1 U513 ( .A1(n563), .A2(n583), .ZN(n361) );
  NAND2_X1 U514 ( .A1(n653), .A2(n652), .ZN(n362) );
  NAND2_X1 U515 ( .A1(n653), .A2(n652), .ZN(n448) );
  BUF_X1 U516 ( .A(n681), .Z(n690) );
  NOR2_X1 U517 ( .A1(n608), .A2(n360), .ZN(n363) );
  NAND2_X1 U518 ( .A1(n363), .A2(n469), .ZN(n366) );
  NAND2_X1 U519 ( .A1(n364), .A2(n365), .ZN(n367) );
  NAND2_X1 U520 ( .A1(n367), .A2(n366), .ZN(n610) );
  INV_X1 U521 ( .A(n609), .ZN(n364) );
  INV_X1 U522 ( .A(n469), .ZN(n365) );
  XNOR2_X1 U523 ( .A(n592), .B(KEYINPUT35), .ZN(n607) );
  NAND2_X1 U524 ( .A1(n368), .A2(n369), .ZN(n604) );
  OR2_X1 U525 ( .A1(n698), .A2(n416), .ZN(n369) );
  NAND2_X1 U526 ( .A1(n361), .A2(n411), .ZN(n410) );
  INV_X1 U527 ( .A(n387), .ZN(n370) );
  NAND2_X1 U528 ( .A1(n377), .A2(n378), .ZN(n371) );
  NAND2_X1 U529 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U530 ( .A(n377), .ZN(n376) );
  NAND2_X1 U531 ( .A1(n382), .A2(n381), .ZN(n377) );
  NAND2_X1 U532 ( .A1(n392), .A2(n391), .ZN(n382) );
  NAND2_X1 U533 ( .A1(n386), .A2(n595), .ZN(n415) );
  OR2_X1 U534 ( .A1(n386), .A2(n443), .ZN(n442) );
  XNOR2_X2 U535 ( .A(n599), .B(KEYINPUT97), .ZN(n386) );
  NOR2_X2 U536 ( .A1(n387), .A2(n500), .ZN(n501) );
  INV_X1 U537 ( .A(n758), .ZN(n424) );
  NAND2_X1 U538 ( .A1(n395), .A2(n451), .ZN(n394) );
  XNOR2_X1 U539 ( .A(n707), .B(KEYINPUT87), .ZN(n403) );
  NAND2_X1 U540 ( .A1(n606), .A2(n605), .ZN(n608) );
  XNOR2_X1 U541 ( .A(n436), .B(n388), .ZN(n506) );
  XNOR2_X1 U542 ( .A(n437), .B(n502), .ZN(n388) );
  NOR2_X1 U543 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X2 U544 ( .A(n389), .B(n353), .ZN(n600) );
  AND2_X2 U545 ( .A1(n445), .A2(n349), .ZN(n465) );
  INV_X1 U546 ( .A(n401), .ZN(n404) );
  NAND2_X1 U547 ( .A1(n782), .A2(n453), .ZN(n391) );
  INV_X1 U548 ( .A(n782), .ZN(n393) );
  NAND2_X1 U549 ( .A1(n396), .A2(KEYINPUT76), .ZN(n395) );
  INV_X1 U550 ( .A(n403), .ZN(n396) );
  NAND2_X1 U551 ( .A1(n404), .A2(n399), .ZN(n398) );
  NAND2_X1 U552 ( .A1(n568), .A2(KEYINPUT32), .ZN(n414) );
  NAND2_X1 U553 ( .A1(n712), .A2(n355), .ZN(n418) );
  NAND2_X1 U554 ( .A1(n582), .A2(n731), .ZN(n598) );
  NAND2_X1 U555 ( .A1(n610), .A2(n611), .ZN(n613) );
  NOR2_X2 U556 ( .A1(n718), .A2(n656), .ZN(n423) );
  XNOR2_X1 U557 ( .A(n651), .B(n650), .ZN(n718) );
  XNOR2_X2 U558 ( .A(n423), .B(KEYINPUT64), .ZN(n681) );
  NAND2_X1 U559 ( .A1(n424), .A2(n465), .ZN(n653) );
  NOR2_X1 U560 ( .A1(n758), .A2(n464), .ZN(n651) );
  XNOR2_X2 U561 ( .A(n428), .B(n427), .ZN(n593) );
  INV_X1 U562 ( .A(G140), .ZN(n429) );
  NAND2_X1 U563 ( .A1(n433), .A2(n432), .ZN(n431) );
  NOR2_X1 U564 ( .A1(n601), .A2(n435), .ZN(n432) );
  INV_X1 U565 ( .A(n600), .ZN(n433) );
  NAND2_X1 U566 ( .A1(n646), .A2(n639), .ZN(n624) );
  INV_X1 U567 ( .A(n594), .ZN(n444) );
  NAND2_X1 U568 ( .A1(n350), .A2(n445), .ZN(n464) );
  NOR2_X1 U569 ( .A1(n635), .A2(n634), .ZN(n447) );
  INV_X1 U570 ( .A(n634), .ZN(n446) );
  AND2_X1 U571 ( .A1(n447), .A2(n637), .ZN(n707) );
  XNOR2_X2 U572 ( .A(G143), .B(G128), .ZN(n510) );
  NAND2_X1 U573 ( .A1(n448), .A2(n655), .ZN(n656) );
  XNOR2_X1 U574 ( .A(n362), .B(KEYINPUT85), .ZN(n717) );
  NAND2_X1 U575 ( .A1(n672), .A2(n654), .ZN(n449) );
  XNOR2_X1 U576 ( .A(n450), .B(n766), .ZN(n672) );
  XNOR2_X1 U577 ( .A(n482), .B(n532), .ZN(n450) );
  NAND2_X1 U578 ( .A1(n783), .A2(KEYINPUT46), .ZN(n451) );
  INV_X1 U579 ( .A(KEYINPUT46), .ZN(n453) );
  NAND2_X1 U580 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U581 ( .A1(n720), .A2(n455), .ZN(n458) );
  INV_X1 U582 ( .A(n719), .ZN(n456) );
  INV_X1 U583 ( .A(n750), .ZN(n644) );
  XNOR2_X2 U584 ( .A(n460), .B(G146), .ZN(n504) );
  XNOR2_X2 U585 ( .A(n462), .B(n461), .ZN(n731) );
  NAND2_X1 U586 ( .A1(n581), .A2(n729), .ZN(n462) );
  NAND2_X1 U587 ( .A1(n682), .A2(n557), .ZN(n463) );
  BUF_X1 U588 ( .A(n581), .Z(n574) );
  AND2_X1 U589 ( .A1(G227), .A2(n777), .ZN(n466) );
  XNOR2_X1 U590 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n468) );
  OR2_X1 U591 ( .A1(KEYINPUT44), .A2(KEYINPUT73), .ZN(n469) );
  AND2_X1 U592 ( .A1(KEYINPUT44), .A2(KEYINPUT73), .ZN(n470) );
  NOR2_X1 U593 ( .A1(n603), .A2(n470), .ZN(n471) );
  XNOR2_X1 U594 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U595 ( .A(n547), .B(n466), .ZN(n531) );
  BUF_X1 U596 ( .A(n657), .Z(n658) );
  XNOR2_X2 U597 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n473) );
  NAND2_X1 U598 ( .A1(n511), .A2(G224), .ZN(n472) );
  XNOR2_X1 U599 ( .A(n472), .B(n473), .ZN(n474) );
  XNOR2_X1 U600 ( .A(n474), .B(n504), .ZN(n477) );
  XNOR2_X1 U601 ( .A(n510), .B(n475), .ZN(n476) );
  XNOR2_X1 U602 ( .A(n477), .B(n476), .ZN(n482) );
  INV_X1 U603 ( .A(n478), .ZN(n480) );
  XNOR2_X1 U604 ( .A(KEYINPUT78), .B(G110), .ZN(n479) );
  XNOR2_X1 U605 ( .A(n480), .B(n479), .ZN(n765) );
  XOR2_X1 U606 ( .A(KEYINPUT67), .B(G101), .Z(n535) );
  INV_X1 U607 ( .A(n535), .ZN(n481) );
  XNOR2_X1 U608 ( .A(n765), .B(n481), .ZN(n532) );
  INV_X1 U609 ( .A(KEYINPUT72), .ZN(n483) );
  XNOR2_X1 U610 ( .A(n483), .B(G113), .ZN(n485) );
  XNOR2_X1 U611 ( .A(G119), .B(G116), .ZN(n484) );
  XNOR2_X1 U612 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U613 ( .A(n487), .B(n486), .ZN(n541) );
  INV_X1 U614 ( .A(G902), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n557), .A2(n489), .ZN(n493) );
  NAND2_X1 U616 ( .A1(n493), .A2(G210), .ZN(n492) );
  INV_X1 U617 ( .A(KEYINPUT84), .ZN(n490) );
  XNOR2_X1 U618 ( .A(n490), .B(KEYINPUT95), .ZN(n491) );
  NAND2_X1 U619 ( .A1(n493), .A2(G214), .ZN(n719) );
  NAND2_X1 U620 ( .A1(n614), .A2(n719), .ZN(n495) );
  INV_X1 U621 ( .A(KEYINPUT19), .ZN(n494) );
  XOR2_X1 U622 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n497) );
  XNOR2_X1 U623 ( .A(n497), .B(n496), .ZN(n498) );
  NAND2_X1 U624 ( .A1(G952), .A2(n498), .ZN(n749) );
  NOR2_X1 U625 ( .A1(n749), .A2(G953), .ZN(n573) );
  NAND2_X1 U626 ( .A1(G902), .A2(n498), .ZN(n569) );
  XOR2_X1 U627 ( .A(G898), .B(KEYINPUT96), .Z(n762) );
  NAND2_X1 U628 ( .A1(G953), .A2(n762), .ZN(n769) );
  NOR2_X1 U629 ( .A1(n569), .A2(n769), .ZN(n499) );
  NOR2_X1 U630 ( .A1(n573), .A2(n499), .ZN(n500) );
  XNOR2_X2 U631 ( .A(n501), .B(n467), .ZN(n599) );
  XNOR2_X1 U632 ( .A(G113), .B(G143), .ZN(n502) );
  XNOR2_X1 U633 ( .A(G131), .B(KEYINPUT12), .ZN(n503) );
  XNOR2_X1 U634 ( .A(n506), .B(n548), .ZN(n666) );
  INV_X1 U635 ( .A(KEYINPUT13), .ZN(n508) );
  AND2_X1 U636 ( .A1(G217), .A2(n551), .ZN(n512) );
  XNOR2_X1 U637 ( .A(n529), .B(n512), .ZN(n520) );
  XNOR2_X1 U638 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U639 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U640 ( .A(n518), .B(n517), .Z(n519) );
  XNOR2_X1 U641 ( .A(n520), .B(n519), .ZN(n686) );
  NAND2_X1 U642 ( .A1(n686), .A2(n557), .ZN(n522) );
  INV_X1 U643 ( .A(G478), .ZN(n521) );
  XNOR2_X1 U644 ( .A(n522), .B(n521), .ZN(n601) );
  INV_X1 U645 ( .A(n601), .ZN(n589) );
  NOR2_X1 U646 ( .A1(n600), .A2(n589), .ZN(n642) );
  NAND2_X1 U647 ( .A1(G234), .A2(n654), .ZN(n523) );
  XNOR2_X1 U648 ( .A(KEYINPUT20), .B(n523), .ZN(n558) );
  AND2_X1 U649 ( .A1(n558), .A2(G221), .ZN(n525) );
  XNOR2_X1 U650 ( .A(KEYINPUT98), .B(KEYINPUT21), .ZN(n524) );
  XNOR2_X1 U651 ( .A(n525), .B(n524), .ZN(n729) );
  AND2_X1 U652 ( .A1(n642), .A2(n729), .ZN(n526) );
  NAND2_X1 U653 ( .A1(n599), .A2(n526), .ZN(n528) );
  XNOR2_X1 U654 ( .A(KEYINPUT75), .B(KEYINPUT22), .ZN(n527) );
  XNOR2_X1 U655 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n533) );
  INV_X1 U656 ( .A(n732), .ZN(n618) );
  NAND2_X1 U657 ( .A1(n563), .A2(n618), .ZN(n534) );
  XNOR2_X1 U658 ( .A(n534), .B(KEYINPUT109), .ZN(n562) );
  XNOR2_X1 U659 ( .A(n536), .B(n535), .ZN(n545) );
  NAND2_X1 U660 ( .A1(n537), .A2(G210), .ZN(n538) );
  XNOR2_X1 U661 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U662 ( .A(n540), .B(KEYINPUT5), .Z(n543) );
  INV_X1 U663 ( .A(n541), .ZN(n542) );
  XNOR2_X1 U664 ( .A(n545), .B(n544), .ZN(n657) );
  NAND2_X1 U665 ( .A1(n657), .A2(n557), .ZN(n546) );
  XNOR2_X2 U666 ( .A(n546), .B(G472), .ZN(n632) );
  XNOR2_X1 U667 ( .A(n550), .B(n549), .ZN(n555) );
  NAND2_X1 U668 ( .A1(n551), .A2(G221), .ZN(n553) );
  XNOR2_X1 U669 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U670 ( .A(n555), .B(n554), .Z(n556) );
  XNOR2_X1 U671 ( .A(n772), .B(n556), .ZN(n682) );
  NAND2_X1 U672 ( .A1(n558), .A2(G217), .ZN(n559) );
  XOR2_X1 U673 ( .A(n559), .B(KEYINPUT25), .Z(n560) );
  INV_X1 U674 ( .A(n574), .ZN(n566) );
  NOR2_X1 U675 ( .A1(n738), .A2(n574), .ZN(n561) );
  NAND2_X1 U676 ( .A1(n562), .A2(n561), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(G110), .ZN(G12) );
  XOR2_X1 U678 ( .A(n568), .B(KEYINPUT89), .Z(n565) );
  NAND2_X1 U679 ( .A1(n574), .A2(n618), .ZN(n564) );
  NOR2_X1 U680 ( .A1(n565), .A2(n564), .ZN(n603) );
  XOR2_X1 U681 ( .A(G101), .B(n603), .Z(G3) );
  NAND2_X1 U682 ( .A1(n566), .A2(n732), .ZN(n567) );
  XNOR2_X1 U683 ( .A(n606), .B(G119), .ZN(G21) );
  NOR2_X1 U684 ( .A1(G900), .A2(n569), .ZN(n570) );
  NAND2_X1 U685 ( .A1(G953), .A2(n570), .ZN(n571) );
  XOR2_X1 U686 ( .A(KEYINPUT110), .B(n571), .Z(n572) );
  NOR2_X1 U687 ( .A1(n573), .A2(n572), .ZN(n634) );
  NOR2_X1 U688 ( .A1(n634), .A2(n574), .ZN(n620) );
  NAND2_X1 U689 ( .A1(n729), .A2(n719), .ZN(n576) );
  AND2_X1 U690 ( .A1(n600), .A2(n601), .ZN(n710) );
  INV_X1 U691 ( .A(n710), .ZN(n639) );
  NOR2_X1 U692 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U693 ( .A(n615), .B(KEYINPUT111), .ZN(n578) );
  NOR2_X1 U694 ( .A1(n732), .A2(n578), .ZN(n579) );
  INV_X1 U695 ( .A(n614), .ZN(n638) );
  XNOR2_X1 U696 ( .A(n649), .B(G140), .ZN(G42) );
  INV_X1 U697 ( .A(n583), .ZN(n584) );
  NAND2_X1 U698 ( .A1(n347), .A2(n584), .ZN(n586) );
  INV_X1 U699 ( .A(KEYINPUT33), .ZN(n585) );
  XOR2_X1 U700 ( .A(KEYINPUT83), .B(KEYINPUT34), .Z(n587) );
  XNOR2_X1 U701 ( .A(n588), .B(n587), .ZN(n591) );
  NAND2_X1 U702 ( .A1(n600), .A2(n589), .ZN(n636) );
  XOR2_X1 U703 ( .A(KEYINPUT82), .B(n636), .Z(n590) );
  NAND2_X1 U704 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U705 ( .A(n360), .B(G122), .Z(G24) );
  INV_X1 U706 ( .A(n593), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n731), .A2(n631), .ZN(n594) );
  INV_X1 U708 ( .A(KEYINPUT99), .ZN(n595) );
  INV_X1 U709 ( .A(n738), .ZN(n597) );
  NOR2_X1 U710 ( .A1(n598), .A2(n597), .ZN(n740) );
  INV_X1 U711 ( .A(n624), .ZN(n725) );
  INV_X1 U712 ( .A(n627), .ZN(n602) );
  INV_X1 U713 ( .A(KEYINPUT45), .ZN(n612) );
  NAND2_X1 U714 ( .A1(n615), .A2(n348), .ZN(n616) );
  NAND2_X1 U715 ( .A1(n620), .A2(n619), .ZN(n622) );
  XNOR2_X1 U716 ( .A(n622), .B(n621), .ZN(n623) );
  NAND2_X1 U717 ( .A1(n351), .A2(n624), .ZN(n625) );
  NAND2_X1 U718 ( .A1(n625), .A2(KEYINPUT47), .ZN(n630) );
  XOR2_X1 U719 ( .A(KEYINPUT47), .B(KEYINPUT69), .Z(n626) );
  NAND2_X1 U720 ( .A1(n351), .A2(n628), .ZN(n629) );
  NAND2_X1 U721 ( .A1(n632), .A2(n719), .ZN(n633) );
  NOR2_X1 U722 ( .A1(n638), .A2(n636), .ZN(n637) );
  NOR2_X1 U723 ( .A1(n647), .A2(n639), .ZN(n641) );
  INV_X1 U724 ( .A(n642), .ZN(n723) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U727 ( .A(n648), .B(KEYINPUT115), .ZN(n781) );
  INV_X1 U728 ( .A(KEYINPUT2), .ZN(n652) );
  INV_X1 U729 ( .A(n654), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n681), .A2(G472), .ZN(n660) );
  XNOR2_X1 U731 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X2 U732 ( .A1(n661), .A2(n696), .ZN(n663) );
  XNOR2_X1 U733 ( .A(KEYINPUT91), .B(KEYINPUT63), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(G57) );
  NAND2_X1 U735 ( .A1(n681), .A2(G475), .ZN(n668) );
  XOR2_X1 U736 ( .A(KEYINPUT66), .B(KEYINPUT124), .Z(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(KEYINPUT59), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n668), .B(n667), .ZN(n669) );
  NOR2_X2 U739 ( .A1(n669), .A2(n696), .ZN(n671) );
  XOR2_X1 U740 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(G60) );
  NAND2_X1 U742 ( .A1(n681), .A2(G210), .ZN(n678) );
  BUF_X1 U743 ( .A(n672), .Z(n673) );
  XOR2_X1 U744 ( .A(KEYINPUT55), .B(KEYINPUT92), .Z(n675) );
  XNOR2_X1 U745 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n674) );
  XOR2_X1 U746 ( .A(n675), .B(n674), .Z(n676) );
  XNOR2_X1 U747 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U748 ( .A1(n679), .A2(n696), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n680), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U750 ( .A1(n690), .A2(G217), .ZN(n684) );
  XNOR2_X1 U751 ( .A(n682), .B(KEYINPUT127), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n684), .B(n683), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n685), .A2(n696), .ZN(G66) );
  NAND2_X1 U754 ( .A1(n690), .A2(G478), .ZN(n688) );
  XOR2_X1 U755 ( .A(n686), .B(KEYINPUT126), .Z(n687) );
  XNOR2_X1 U756 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n689), .A2(n696), .ZN(G63) );
  NAND2_X1 U758 ( .A1(n690), .A2(G469), .ZN(n695) );
  XNOR2_X1 U759 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT58), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n695), .B(n694), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(G54) );
  BUF_X1 U764 ( .A(n698), .Z(n701) );
  NAND2_X1 U765 ( .A1(n701), .A2(n710), .ZN(n699) );
  XNOR2_X1 U766 ( .A(n699), .B(KEYINPUT116), .ZN(n700) );
  XNOR2_X1 U767 ( .A(G104), .B(n700), .ZN(G6) );
  XOR2_X1 U768 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U769 ( .A1(n701), .A2(n713), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U771 ( .A(G107), .B(n704), .ZN(G9) );
  XOR2_X1 U772 ( .A(G128), .B(KEYINPUT29), .Z(n706) );
  NAND2_X1 U773 ( .A1(n351), .A2(n713), .ZN(n705) );
  XNOR2_X1 U774 ( .A(n706), .B(n705), .ZN(G30) );
  XOR2_X1 U775 ( .A(G143), .B(n707), .Z(G45) );
  XOR2_X1 U776 ( .A(G146), .B(KEYINPUT117), .Z(n709) );
  NAND2_X1 U777 ( .A1(n351), .A2(n710), .ZN(n708) );
  XNOR2_X1 U778 ( .A(n709), .B(n708), .ZN(G48) );
  NAND2_X1 U779 ( .A1(n712), .A2(n710), .ZN(n711) );
  XNOR2_X1 U780 ( .A(n711), .B(G113), .ZN(G15) );
  NAND2_X1 U781 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U782 ( .A(n714), .B(G116), .ZN(G18) );
  XNOR2_X1 U783 ( .A(G125), .B(n715), .ZN(n716) );
  XNOR2_X1 U784 ( .A(n716), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n756) );
  NOR2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U787 ( .A(n721), .B(KEYINPUT120), .ZN(n722) );
  NOR2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U789 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U791 ( .A1(n751), .A2(n728), .ZN(n745) );
  NOR2_X1 U792 ( .A1(n729), .A2(n574), .ZN(n730) );
  XNOR2_X1 U793 ( .A(KEYINPUT49), .B(n730), .ZN(n736) );
  OR2_X1 U794 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U795 ( .A(n733), .B(KEYINPUT118), .ZN(n734) );
  XNOR2_X1 U796 ( .A(KEYINPUT50), .B(n734), .ZN(n735) );
  NAND2_X1 U797 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U798 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U799 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U800 ( .A(n741), .B(KEYINPUT51), .ZN(n742) );
  XNOR2_X1 U801 ( .A(n742), .B(KEYINPUT119), .ZN(n743) );
  NOR2_X1 U802 ( .A1(n743), .A2(n750), .ZN(n744) );
  NOR2_X1 U803 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U804 ( .A(n746), .B(KEYINPUT121), .Z(n747) );
  XNOR2_X1 U805 ( .A(KEYINPUT52), .B(n747), .ZN(n748) );
  NOR2_X1 U806 ( .A1(n749), .A2(n748), .ZN(n753) );
  NOR2_X1 U807 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U808 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U809 ( .A1(n754), .A2(n777), .ZN(n755) );
  NOR2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n757), .B(KEYINPUT53), .ZN(G75) );
  BUF_X1 U812 ( .A(n758), .Z(n759) );
  NOR2_X1 U813 ( .A1(n759), .A2(G953), .ZN(n764) );
  NAND2_X1 U814 ( .A1(G953), .A2(G224), .ZN(n760) );
  XOR2_X1 U815 ( .A(KEYINPUT61), .B(n760), .Z(n761) );
  NOR2_X1 U816 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U817 ( .A1(n764), .A2(n763), .ZN(n771) );
  XNOR2_X1 U818 ( .A(n765), .B(G101), .ZN(n767) );
  XOR2_X1 U819 ( .A(n767), .B(n766), .Z(n768) );
  NAND2_X1 U820 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(G69) );
  XNOR2_X1 U822 ( .A(n773), .B(n772), .ZN(n776) );
  XNOR2_X1 U823 ( .A(G227), .B(n776), .ZN(n774) );
  NAND2_X1 U824 ( .A1(G900), .A2(n774), .ZN(n775) );
  NAND2_X1 U825 ( .A1(n775), .A2(G953), .ZN(n780) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n780), .A2(n779), .ZN(G72) );
  XNOR2_X1 U828 ( .A(G134), .B(n781), .ZN(G36) );
  XOR2_X1 U829 ( .A(n782), .B(G131), .Z(G33) );
  XOR2_X1 U830 ( .A(G137), .B(n783), .Z(G39) );
endmodule

