//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n220), .B1(new_n212), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n207), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n210), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n234), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT66), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  NAND2_X1  g0049(.A1(G20), .A2(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n217), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n217), .A2(G33), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT15), .B(G87), .ZN(new_n255));
  OAI221_X1 g0055(.A(new_n250), .B1(new_n251), .B2(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n216), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n260), .A2(new_n217), .A3(G1), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n256), .A2(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n258), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(G77), .A3(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n263), .A2(KEYINPUT68), .A3(G77), .A4(new_n265), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n278), .B1(G244), .B2(new_n281), .ZN(new_n282));
  XNOR2_X1  g0082(.A(KEYINPUT3), .B(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G232), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G238), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n283), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n287), .B(new_n288), .C1(G107), .C2(new_n283), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G169), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n271), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  INV_X1    g0094(.A(new_n290), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n293), .A2(KEYINPUT71), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n271), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n204), .A2(G20), .ZN(new_n301));
  INV_X1    g0101(.A(G150), .ZN(new_n302));
  OAI221_X1 g0102(.A(new_n301), .B1(new_n302), .B2(new_n253), .C1(new_n251), .C2(new_n254), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n258), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n263), .A2(G50), .A3(new_n265), .ZN(new_n305));
  INV_X1    g0105(.A(new_n261), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(G50), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT67), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n307), .B(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n283), .A2(G223), .A3(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n283), .A2(new_n285), .ZN(new_n312));
  INV_X1    g0112(.A(G222), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n311), .B1(new_n259), .B2(new_n283), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n288), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n278), .B1(G226), .B2(new_n281), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n294), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n310), .B(new_n319), .C1(G169), .C2(new_n318), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(G226), .A2(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n236), .A2(G1698), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n283), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n288), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n277), .B1(new_n221), .B2(new_n280), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n276), .B1(new_n324), .B2(new_n325), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT13), .B1(new_n332), .B2(new_n328), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  NOR2_X1   g0135(.A1(G20), .A2(G33), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(G50), .B1(G20), .B2(new_n212), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n259), .B2(new_n254), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n258), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT11), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n261), .A2(new_n212), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT12), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n263), .A2(G68), .A3(new_n265), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n341), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n335), .B(new_n347), .C1(new_n348), .C2(new_n334), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n300), .A2(new_n321), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT69), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n262), .A2(new_n270), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n290), .A2(G200), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n352), .B1(new_n262), .B2(new_n270), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT70), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n356), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT70), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n358), .A2(new_n359), .A3(new_n353), .A4(new_n354), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n295), .A2(G190), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n330), .B1(new_n327), .B2(new_n329), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n332), .A2(new_n328), .A3(KEYINPUT13), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n363), .B(G169), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n331), .A2(G179), .A3(new_n333), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n363), .B1(new_n334), .B2(G169), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n346), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n351), .A2(new_n362), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n310), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n373), .B(KEYINPUT72), .ZN(new_n374));
  INV_X1    g0174(.A(new_n310), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT9), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n318), .A2(G190), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n317), .A2(G200), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(KEYINPUT10), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT72), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n373), .B(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT10), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(KEYINPUT75), .A2(KEYINPUT18), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n251), .B1(new_n264), .B2(G20), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n388), .A2(new_n263), .B1(new_n261), .B2(new_n251), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n258), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT3), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G33), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n395), .B2(new_n217), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n397), .B(G20), .C1(new_n392), .C2(new_n394), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT73), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n217), .B1(new_n213), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n336), .A2(G159), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n400), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n406), .B2(new_n201), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n403), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n399), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n391), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n399), .A2(new_n409), .A3(KEYINPUT16), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n390), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n392), .A2(new_n394), .A3(G223), .A4(new_n285), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT74), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n283), .A2(KEYINPUT74), .A3(G223), .A4(new_n285), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n283), .A2(G226), .A3(G1698), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n288), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n277), .B1(new_n280), .B2(new_n236), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n291), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g0225(.A(new_n294), .B(new_n423), .C1(new_n421), .C2(new_n288), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n387), .B1(new_n414), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT17), .ZN(new_n429));
  AND3_X1   g0229(.A1(new_n407), .A2(KEYINPUT73), .A3(new_n403), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT73), .B1(new_n407), .B2(new_n403), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n397), .B1(new_n283), .B2(G20), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n395), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n212), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n411), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n413), .A3(new_n258), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n389), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n422), .A2(G190), .A3(new_n424), .ZN(new_n439));
  INV_X1    g0239(.A(G200), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n423), .B1(new_n421), .B2(new_n288), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n429), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n441), .A2(new_n440), .ZN(new_n444));
  AOI211_X1 g0244(.A(new_n348), .B(new_n423), .C1(new_n421), .C2(new_n288), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n414), .A2(new_n446), .A3(KEYINPUT17), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n428), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n414), .A2(new_n427), .A3(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n441), .A2(G179), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n291), .B2(new_n441), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n438), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT75), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n371), .A2(new_n386), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n264), .A2(G33), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n263), .A2(G116), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G116), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n261), .A2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n257), .A2(new_n216), .B1(G20), .B2(new_n460), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n463), .B(new_n217), .C1(G33), .C2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n462), .B2(new_n465), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n459), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT21), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n272), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n273), .A2(G1), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT5), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT77), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G41), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n472), .A2(G274), .A3(new_n276), .A4(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n475), .A2(new_n471), .A3(new_n470), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G270), .A3(new_n276), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n392), .A2(new_n394), .A3(G264), .A4(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n392), .A2(new_n394), .A3(G257), .A4(new_n285), .ZN(new_n481));
  INV_X1    g0281(.A(G303), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n481), .C1(new_n482), .C2(new_n283), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n288), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n469), .B(new_n291), .C1(new_n479), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(new_n476), .A3(new_n478), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n294), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n468), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n468), .B1(new_n486), .B2(G200), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n348), .B2(new_n486), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(G169), .A3(new_n468), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n491), .A2(new_n492), .A3(new_n469), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n491), .B2(new_n469), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n488), .B(new_n490), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n283), .A2(new_n217), .A3(G87), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT81), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT81), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n283), .A2(new_n498), .A3(new_n217), .A4(G87), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(KEYINPUT22), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(KEYINPUT23), .B1(new_n217), .B2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT23), .ZN(new_n502));
  INV_X1    g0302(.A(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(G20), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n217), .A2(G33), .A3(G116), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT82), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT22), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n496), .A2(KEYINPUT81), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n500), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT83), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n500), .A2(new_n507), .A3(KEYINPUT83), .A4(new_n509), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(KEYINPUT24), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n510), .A2(new_n511), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n258), .A3(new_n516), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n263), .A2(new_n458), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT25), .B1(new_n261), .B2(new_n503), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n261), .A2(KEYINPUT25), .A3(new_n503), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n518), .A2(G107), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n283), .A2(G257), .A3(G1698), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G294), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n523), .B(new_n524), .C1(new_n312), .C2(new_n223), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n477), .A2(new_n276), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n525), .A2(new_n288), .B1(G264), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n476), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n440), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(G190), .B2(new_n528), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n517), .A2(new_n522), .A3(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n522), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n516), .A2(new_n258), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n532), .B1(new_n534), .B2(new_n514), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n291), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G179), .B2(new_n528), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n531), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT78), .B1(new_n273), .B2(G1), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT78), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(new_n264), .A3(G45), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n276), .A2(new_n539), .A3(new_n541), .A4(G250), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n276), .A2(G274), .A3(new_n471), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n283), .A2(G238), .A3(new_n285), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n283), .A2(G244), .A3(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n548), .B2(new_n288), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n549), .A2(new_n440), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(G190), .B2(new_n549), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n217), .B1(new_n325), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n222), .A2(new_n464), .A3(new_n503), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n392), .A2(new_n394), .A3(new_n217), .A4(G68), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n552), .B1(new_n254), .B2(new_n464), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT79), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n391), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT79), .A4(new_n557), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(new_n261), .B2(new_n255), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n518), .A2(G87), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n549), .A2(G169), .ZN(new_n566));
  AOI211_X1 g0366(.A(G179), .B(new_n544), .C1(new_n548), .C2(new_n288), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n255), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n518), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n562), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n551), .A2(new_n565), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT6), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n573), .A2(new_n464), .A3(G107), .ZN(new_n574));
  XNOR2_X1  g0374(.A(G97), .B(G107), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n574), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n576), .A2(new_n217), .B1(new_n259), .B2(new_n253), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n503), .B1(new_n433), .B2(new_n434), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n258), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n306), .A2(G97), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n518), .B2(G97), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(G274), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n477), .A2(new_n583), .A3(new_n288), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(G257), .B2(new_n526), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n392), .A2(new_n394), .A3(G244), .A4(new_n285), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n392), .A2(new_n394), .A3(G250), .A4(G1698), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n463), .B(new_n590), .C1(new_n586), .C2(new_n587), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n288), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(new_n592), .A3(G190), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n526), .A2(G257), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n476), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT76), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n283), .A2(KEYINPUT4), .A3(G244), .A4(new_n285), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n588), .A2(new_n598), .A3(new_n463), .A4(new_n590), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(KEYINPUT76), .A3(new_n288), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n595), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n582), .B(new_n593), .C1(new_n601), .C2(new_n440), .ZN(new_n602));
  INV_X1    g0402(.A(new_n600), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT76), .B1(new_n599), .B2(new_n288), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n294), .B(new_n585), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n585), .A2(new_n592), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n291), .B1(new_n579), .B2(new_n581), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n572), .A2(new_n602), .A3(new_n608), .ZN(new_n609));
  NOR4_X1   g0409(.A1(new_n457), .A2(new_n495), .A3(new_n538), .A4(new_n609), .ZN(G372));
  OAI21_X1  g0410(.A(KEYINPUT18), .B1(new_n414), .B2(new_n427), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n438), .A2(new_n452), .A3(new_n450), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n370), .B1(new_n299), .B2(new_n350), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n443), .A2(new_n447), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n321), .B1(new_n386), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n566), .A2(KEYINPUT84), .ZN(new_n620));
  INV_X1    g0420(.A(new_n567), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n549), .B2(G169), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n620), .A2(new_n571), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n537), .B1(new_n517), .B2(new_n522), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT86), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n491), .A2(new_n469), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT80), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n491), .A2(new_n492), .A3(new_n469), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n628), .B1(new_n632), .B2(new_n488), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n488), .B(new_n628), .C1(new_n493), .C2(new_n494), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n627), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n517), .A2(new_n522), .A3(new_n530), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n602), .A2(new_n608), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT85), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n562), .A2(new_n639), .A3(new_n563), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n562), .B2(new_n563), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n551), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n624), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n637), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n625), .B1(new_n636), .B2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n605), .A2(new_n607), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n642), .A3(new_n624), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT87), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n572), .A2(new_n646), .A3(KEYINPUT26), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n647), .A2(KEYINPUT87), .A3(new_n648), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n619), .B1(new_n656), .B2(new_n457), .ZN(G369));
  INV_X1    g0457(.A(new_n495), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n264), .A2(new_n217), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n468), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n488), .B1(new_n493), .B2(new_n494), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT86), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n634), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n666), .B1(new_n669), .B2(new_n665), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n664), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n535), .A2(new_n673), .ZN(new_n674));
  OAI22_X1  g0474(.A1(new_n538), .A2(new_n674), .B1(new_n627), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n637), .A2(new_n626), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n667), .A2(new_n673), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n626), .A2(new_n673), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n676), .A2(new_n683), .ZN(G399));
  NOR2_X1   g0484(.A1(new_n554), .A2(G116), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n208), .A2(new_n272), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(new_n686), .A3(G1), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n214), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT30), .ZN(new_n690));
  INV_X1    g0490(.A(new_n487), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n527), .A2(new_n549), .A3(new_n585), .A4(new_n592), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n549), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n528), .A2(new_n294), .A3(new_n486), .A4(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n601), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT88), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n527), .A2(new_n549), .ZN(new_n698));
  INV_X1    g0498(.A(new_n606), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(KEYINPUT30), .A4(new_n487), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n696), .A2(KEYINPUT88), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT31), .B(new_n664), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n693), .B(new_n700), .C1(new_n601), .C2(new_n695), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n664), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR4_X1   g0508(.A1(new_n538), .A2(new_n609), .A3(new_n495), .A4(new_n664), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n488), .B(new_n632), .C1(new_n535), .C2(new_n537), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n602), .A2(new_n608), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n642), .A2(new_n624), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n715), .A2(new_n531), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n568), .A2(new_n571), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n549), .A2(G190), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n440), .B2(new_n549), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n719), .B1(new_n564), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n648), .B1(new_n722), .B2(new_n608), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n646), .A2(new_n642), .A3(KEYINPUT26), .A4(new_n624), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(KEYINPUT89), .A3(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n724), .A2(KEYINPUT89), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n718), .A2(new_n725), .A3(new_n624), .A4(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n714), .B1(new_n727), .B2(new_n673), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n664), .B1(new_n645), .B2(new_n654), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n728), .B1(new_n714), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n713), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n689), .B1(new_n732), .B2(G1), .ZN(G364));
  NOR2_X1   g0533(.A1(new_n260), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n264), .B1(new_n734), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n686), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n672), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G330), .B2(new_n670), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n283), .A2(new_n208), .ZN(new_n741));
  INV_X1    g0541(.A(G355), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n741), .A2(new_n742), .B1(G116), .B2(new_n208), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n248), .A2(G45), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n395), .A2(new_n208), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n745), .B1(new_n273), .B2(new_n215), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n743), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n216), .B1(G20), .B2(new_n291), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n738), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(G20), .B1(new_n756), .B2(new_n348), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT93), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n757), .A2(new_n758), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G294), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  NAND3_X1  g0564(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n348), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n762), .A2(new_n763), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT94), .Z(new_n769));
  NOR2_X1   g0569(.A1(new_n217), .A2(new_n348), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n294), .A2(G200), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n771), .A3(G322), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n217), .A2(G190), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n440), .A2(G179), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G283), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n770), .A2(new_n774), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n772), .B1(new_n775), .B2(new_n776), .C1(new_n482), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n773), .A2(new_n771), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n765), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT33), .B(G317), .Z(new_n783));
  OAI221_X1 g0583(.A(new_n395), .B1(new_n779), .B2(new_n780), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n773), .A2(new_n755), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT92), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT92), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n778), .B(new_n784), .C1(new_n789), .C2(G329), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n769), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n770), .A2(new_n771), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT90), .Z(new_n793));
  OAI22_X1  g0593(.A1(new_n793), .A2(new_n211), .B1(new_n259), .B2(new_n779), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT91), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n789), .A2(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(KEYINPUT32), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n283), .B1(new_n775), .B2(new_n503), .C1(new_n222), .C2(new_n777), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n782), .A2(new_n212), .B1(new_n767), .B2(new_n202), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n762), .ZN(new_n801));
  AOI22_X1  g0601(.A1(KEYINPUT32), .A2(new_n796), .B1(new_n801), .B2(G97), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n795), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n754), .B1(new_n804), .B2(new_n751), .ZN(new_n805));
  INV_X1    g0605(.A(new_n750), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n670), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g0607(.A1(new_n740), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(G396));
  INV_X1    g0609(.A(new_n729), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n673), .B1(new_n262), .B2(new_n270), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n296), .B2(new_n298), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n362), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n300), .A2(new_n811), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n362), .A2(new_n812), .A3(KEYINPUT97), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n810), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT98), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n664), .B1(new_n815), .B2(new_n817), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n653), .A2(new_n652), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT87), .B1(new_n647), .B2(new_n648), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n626), .B1(new_n668), .B2(new_n634), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n717), .A2(new_n716), .A3(new_n531), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n624), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n822), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n821), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n738), .B1(new_n830), .B2(new_n713), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n713), .B2(new_n830), .ZN(new_n832));
  INV_X1    g0632(.A(new_n751), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n749), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n738), .B1(G77), .B2(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n782), .A2(new_n776), .B1(new_n767), .B2(new_n482), .ZN(new_n836));
  INV_X1    g0636(.A(new_n775), .ZN(new_n837));
  INV_X1    g0637(.A(new_n779), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G87), .A2(new_n837), .B1(new_n838), .B2(G116), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n763), .B2(new_n792), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n836), .B(new_n840), .C1(G97), .C2(new_n801), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT95), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n395), .B1(new_n777), .B2(new_n503), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n789), .A2(G311), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n841), .B(new_n844), .C1(new_n842), .C2(new_n843), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n838), .A2(G159), .B1(G137), .B2(new_n766), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n302), .B2(new_n782), .ZN(new_n847));
  INV_X1    g0647(.A(new_n793), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(G143), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n283), .B1(new_n775), .B2(new_n212), .C1(new_n202), .C2(new_n777), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n789), .B2(G132), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n851), .B(new_n853), .C1(new_n211), .C2(new_n762), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n845), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n855), .A2(KEYINPUT96), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n833), .B1(new_n855), .B2(KEYINPUT96), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n835), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n749), .B2(new_n818), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n832), .A2(new_n859), .ZN(G384));
  XNOR2_X1  g0660(.A(new_n576), .B(KEYINPUT99), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT35), .ZN(new_n862));
  OAI211_X1 g0662(.A(G116), .B(new_n218), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT36), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n215), .A2(G77), .A3(new_n401), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n202), .A2(G68), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n264), .B(G13), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n370), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(KEYINPUT101), .B(new_n346), .C1(new_n368), .C2(new_n369), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n346), .A2(new_n664), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n349), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n368), .A2(new_n369), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n346), .B(new_n664), .C1(new_n876), .C2(new_n350), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT102), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n875), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  INV_X1    g0683(.A(new_n662), .ZN(new_n884));
  AND3_X1   g0684(.A1(new_n437), .A2(KEYINPUT103), .A3(new_n389), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT103), .B1(new_n437), .B2(new_n389), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n452), .B1(new_n885), .B2(new_n886), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n414), .A2(new_n446), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n438), .A2(new_n452), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n438), .A2(new_n884), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n889), .A2(new_n892), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n883), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT104), .ZN(new_n897));
  INV_X1    g0697(.A(new_n887), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n455), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT75), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n611), .B2(new_n612), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n428), .A2(new_n443), .A3(new_n447), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n897), .B(new_n898), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n896), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT104), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n907), .A2(new_n903), .B1(new_n895), .B2(new_n891), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n908), .B2(KEYINPUT38), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n362), .A2(new_n812), .A3(KEYINPUT97), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT97), .B1(new_n362), .B2(new_n812), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n673), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n645), .B2(new_n654), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT100), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n299), .A2(new_n664), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n915), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT100), .B1(new_n829), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n882), .B(new_n909), .C1(new_n916), .C2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n613), .A2(new_n662), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n438), .B(new_n884), .C1(new_n613), .C2(new_n615), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n895), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT38), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n905), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT105), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n905), .A2(new_n926), .A3(KEYINPUT105), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n929), .A2(new_n930), .B1(KEYINPUT39), .B2(new_n909), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n871), .A2(new_n872), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n673), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n919), .B(new_n920), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT106), .ZN(new_n935));
  INV_X1    g0735(.A(new_n920), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n905), .A2(KEYINPUT105), .A3(new_n926), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT105), .B1(new_n905), .B2(new_n926), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n891), .A2(new_n895), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n899), .B2(new_n904), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n907), .A2(new_n903), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n940), .A2(new_n883), .B1(new_n941), .B2(new_n896), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT39), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n937), .A2(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n933), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT106), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(new_n919), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n935), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n619), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n727), .A2(new_n673), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT29), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n810), .B2(KEYINPUT29), .ZN(new_n953));
  INV_X1    g0753(.A(new_n457), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n949), .B(new_n955), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n875), .A2(new_n880), .A3(new_n877), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n880), .B1(new_n875), .B2(new_n877), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n818), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n707), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n709), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT40), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n959), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n925), .B1(new_n941), .B2(new_n896), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(KEYINPUT107), .A3(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT107), .ZN(new_n968));
  INV_X1    g0768(.A(new_n609), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n677), .A2(new_n658), .A3(new_n969), .A4(new_n673), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT31), .B1(new_n704), .B2(new_n664), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n974), .A4(new_n818), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n968), .B1(new_n975), .B2(new_n965), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n882), .A2(new_n818), .A3(new_n974), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n963), .B1(new_n942), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n954), .A2(new_n974), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(G330), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n956), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n264), .B2(new_n734), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n956), .A2(new_n984), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n869), .B1(new_n986), .B2(new_n987), .ZN(G367));
  AND3_X1   g0788(.A1(new_n234), .A2(new_n208), .A3(new_n395), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n752), .B1(new_n208), .B2(new_n255), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n738), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(G159), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n782), .A2(new_n992), .B1(new_n779), .B2(new_n202), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT113), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n801), .A2(G68), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n283), .B1(new_n775), .B2(new_n259), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n211), .A2(new_n777), .B1(new_n792), .B2(new_n302), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n997), .B(new_n998), .C1(G143), .C2(new_n766), .ZN(new_n999));
  INV_X1    g0799(.A(G137), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n999), .B1(new_n1000), .B2(new_n788), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n395), .B1(new_n775), .B2(new_n464), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G283), .B2(new_n838), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1003), .B1(new_n788), .B2(new_n1004), .C1(new_n793), .C2(new_n482), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n777), .A2(new_n460), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(KEYINPUT46), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G294), .B2(new_n781), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT112), .B(G311), .Z(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1006), .A2(KEYINPUT46), .B1(new_n1010), .B2(new_n766), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1008), .B(new_n1011), .C1(new_n503), .C2(new_n762), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n996), .A2(new_n1001), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT47), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n991), .B1(new_n1014), .B2(new_n751), .ZN(new_n1015));
  OR3_X1    g0815(.A1(new_n640), .A2(new_n641), .A3(new_n673), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n717), .A2(new_n1016), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n624), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1015), .B1(new_n806), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n582), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n638), .B1(new_n1021), .B2(new_n664), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT109), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n608), .A2(new_n673), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1025), .A2(KEYINPUT42), .A3(new_n680), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT42), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n680), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1023), .A2(new_n626), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n664), .B1(new_n1031), .B2(new_n608), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1026), .B1(new_n1033), .B2(KEYINPUT110), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT110), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1019), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(KEYINPUT108), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT108), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT43), .B1(new_n1019), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1034), .A2(new_n1036), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT43), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1041), .B1(new_n1045), .B2(new_n1037), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1044), .A2(new_n1047), .B1(new_n676), .B2(new_n1025), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n676), .A2(new_n1025), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1043), .C1(new_n1050), .C2(new_n1046), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n1025), .A2(KEYINPUT44), .A3(new_n682), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT44), .B1(new_n1025), .B2(new_n682), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n1056));
  NAND3_X1  g0856(.A1(new_n1028), .A2(new_n683), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1056), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n1025), .B2(new_n682), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n676), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1055), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1061), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n680), .B1(new_n675), .B2(new_n679), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(new_n671), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n731), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n732), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n686), .B(KEYINPUT41), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n736), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1020), .B1(new_n1052), .B2(new_n1071), .ZN(G387));
  INV_X1    g0872(.A(new_n1066), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n731), .A2(new_n1065), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n1074), .A3(new_n737), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1065), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n741), .A2(new_n685), .B1(G107), .B2(new_n208), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n239), .A2(G45), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n685), .ZN(new_n1079));
  AOI211_X1 g0879(.A(G45), .B(new_n1079), .C1(G68), .C2(G77), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n251), .A2(G50), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT50), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n745), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1077), .B1(new_n1078), .B2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n738), .B1(new_n1084), .B2(new_n753), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n801), .A2(new_n569), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n283), .B1(new_n775), .B2(new_n464), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n782), .A2(new_n251), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(G159), .C2(new_n766), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n789), .A2(G150), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n202), .A2(new_n792), .B1(new_n777), .B2(new_n259), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G68), .B2(new_n838), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1086), .A2(new_n1089), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n838), .A2(G303), .B1(G322), .B2(new_n766), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n782), .B2(new_n1009), .C1(new_n793), .C2(new_n1004), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT48), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n777), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n801), .A2(G283), .B1(G294), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT49), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(KEYINPUT114), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n283), .B1(new_n837), .B2(G116), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n764), .C2(new_n788), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1102), .A2(KEYINPUT114), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1093), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1085), .B1(new_n1107), .B2(new_n751), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n675), .A2(new_n806), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n736), .A2(new_n1076), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1075), .A2(new_n1110), .ZN(G393));
  NAND3_X1  g0911(.A1(new_n1062), .A2(new_n1063), .A3(new_n736), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n752), .B1(new_n464), .B2(new_n208), .C1(new_n243), .C2(new_n745), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n738), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n767), .A2(new_n302), .B1(new_n792), .B2(new_n992), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT51), .Z(new_n1116));
  NAND2_X1  g0916(.A1(new_n801), .A2(G77), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n789), .A2(G143), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n283), .B1(new_n775), .B2(new_n222), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n777), .A2(new_n212), .B1(new_n779), .B2(new_n251), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(G50), .C2(new_n781), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n395), .B1(new_n775), .B2(new_n503), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n777), .A2(new_n776), .B1(new_n779), .B2(new_n763), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G303), .C2(new_n781), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n789), .A2(G322), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n460), .C2(new_n762), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n767), .A2(new_n1004), .B1(new_n792), .B2(new_n780), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT52), .Z(new_n1129));
  OAI22_X1  g0929(.A1(new_n1116), .A2(new_n1122), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1114), .B1(new_n1130), .B2(new_n751), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n1028), .B2(new_n806), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1112), .A2(new_n1132), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1067), .A2(new_n737), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1073), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(G390));
  NAND3_X1  g0938(.A1(new_n727), .A2(new_n673), .A3(new_n818), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n917), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n882), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n966), .B(new_n933), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(G330), .B(new_n818), .C1(new_n708), .C2(new_n709), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1144), .A2(new_n1142), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n829), .A2(KEYINPUT100), .A3(new_n917), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n945), .B1(new_n1148), .B2(new_n882), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1143), .B(new_n1145), .C1(new_n1149), .C2(new_n944), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n965), .B(new_n945), .C1(new_n1140), .C2(new_n882), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n882), .B1(new_n916), .B2(new_n918), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n933), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1151), .B1(new_n1153), .B2(new_n931), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n974), .A2(G330), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1155), .A2(new_n959), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n736), .B(new_n1150), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n251), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n738), .B1(new_n1158), .B2(new_n834), .ZN(new_n1159));
  INV_X1    g0959(.A(G132), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n283), .B1(new_n775), .B2(new_n202), .C1(new_n1160), .C2(new_n792), .ZN(new_n1161));
  OR3_X1    g0961(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n302), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT53), .B1(new_n777), .B2(new_n302), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(new_n1163), .C1(new_n767), .C2(new_n1164), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1161), .B(new_n1165), .C1(G125), .C2(new_n789), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT54), .B(G143), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n782), .A2(new_n1000), .B1(new_n779), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n801), .B2(G159), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1169), .A2(KEYINPUT115), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(KEYINPUT115), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1166), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT116), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n395), .B1(new_n777), .B2(new_n222), .C1(new_n503), .C2(new_n782), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G283), .B2(new_n766), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n789), .A2(G294), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n792), .A2(new_n460), .B1(new_n775), .B2(new_n212), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G97), .B2(new_n838), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1117), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1174), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1159), .B1(new_n1182), .B2(new_n751), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n944), .B2(new_n749), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1157), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT117), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT117), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n457), .A2(new_n1155), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n619), .B(new_n1190), .C1(new_n730), .C2(new_n457), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1144), .A2(new_n1142), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1156), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1148), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1142), .B1(new_n1155), .B2(new_n819), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1145), .A2(new_n1141), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1197), .B(new_n1150), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1150), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1197), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n686), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1187), .A2(new_n1189), .B1(new_n1198), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(G378));
  AOI21_X1  g1003(.A(KEYINPUT107), .B1(new_n964), .B2(new_n966), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n975), .A2(new_n965), .A3(new_n968), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G330), .B(new_n979), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n386), .A2(new_n320), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n375), .A2(new_n662), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1208), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n1207), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1206), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1219), .A2(new_n977), .A3(G330), .A4(new_n979), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n934), .A2(KEYINPUT106), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n947), .B1(new_n946), .B2(new_n919), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n935), .A2(new_n948), .A3(new_n1220), .A4(new_n1218), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT120), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1224), .A2(KEYINPUT120), .A3(new_n1225), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1217), .A2(new_n748), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n738), .B1(G50), .B2(new_n834), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n788), .A2(new_n776), .ZN(new_n1233));
  AOI211_X1 g1033(.A(G41), .B(new_n283), .C1(new_n1099), .C2(G77), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n837), .A2(G58), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n1235), .C1(new_n503), .C2(new_n792), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1233), .B(new_n1236), .C1(G116), .C2(new_n766), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n801), .A2(G68), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n838), .A2(new_n569), .B1(G97), .B2(new_n781), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1239), .A2(KEYINPUT118), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT118), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT58), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n252), .A2(new_n272), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n202), .B(new_n1244), .C1(new_n283), .C2(G41), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n1164), .A2(new_n792), .B1(new_n777), .B2(new_n1167), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(G137), .B2(new_n838), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n781), .A2(G132), .B1(new_n766), .B2(G125), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n762), .C2(new_n302), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n789), .A2(G124), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1244), .B1(new_n837), .B2(G159), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1251), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1253), .B(new_n1254), .C1(new_n1249), .C2(new_n1255), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1243), .B(new_n1245), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1232), .B1(new_n1257), .B2(new_n751), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1230), .A2(new_n736), .B1(new_n1231), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1191), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1198), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT57), .B1(new_n1230), .B2(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(KEYINPUT57), .A3(new_n1225), .A4(new_n1224), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n737), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1259), .B1(new_n1262), .B2(new_n1264), .ZN(G375));
  NAND2_X1  g1065(.A1(new_n1196), .A2(new_n1194), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(KEYINPUT121), .A3(new_n736), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n793), .A2(new_n1000), .B1(new_n788), .B2(new_n1164), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G159), .A2(new_n1099), .B1(new_n838), .B2(G150), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1270), .A2(new_n283), .A3(new_n1235), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n1160), .B2(new_n767), .C1(new_n782), .C2(new_n1167), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1269), .B(new_n1272), .C1(G50), .C2(new_n801), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1086), .B1(new_n776), .B2(new_n792), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT124), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(KEYINPUT124), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n788), .A2(new_n482), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n395), .B1(new_n775), .B2(new_n259), .C1(new_n464), .C2(new_n777), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n782), .A2(new_n460), .B1(new_n779), .B2(new_n503), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1280), .A2(KEYINPUT122), .B1(G294), .B2(new_n766), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(KEYINPUT122), .B2(new_n1280), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(KEYINPUT123), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1273), .B1(new_n1279), .B2(new_n1283), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n738), .B1(G68), .B2(new_n834), .C1(new_n1284), .C2(new_n833), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n1142), .B2(new_n748), .ZN(new_n1286));
  AOI21_X1  g1086(.A(KEYINPUT121), .B1(new_n1266), .B2(new_n736), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1268), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1266), .A2(new_n1260), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1070), .A3(new_n1200), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(G381));
  NAND3_X1  g1092(.A1(new_n1075), .A2(new_n808), .A3(new_n1110), .ZN(new_n1293));
  OR4_X1    g1093(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1185), .B1(new_n1201), .B2(new_n1198), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  OR4_X1    g1096(.A1(G375), .A2(new_n1294), .A3(G381), .A4(new_n1296), .ZN(G407));
  NAND2_X1  g1097(.A1(new_n663), .A2(G213), .ZN(new_n1298));
  OR3_X1    g1098(.A1(G375), .A2(new_n1296), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G407), .A2(G213), .A3(new_n1299), .ZN(G409));
  NAND2_X1  g1100(.A1(new_n1200), .A2(KEYINPUT60), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1290), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1301), .A2(KEYINPUT125), .A3(new_n1290), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n686), .B1(new_n1289), .B2(KEYINPUT60), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1307), .A2(G384), .A3(new_n1288), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G384), .B1(new_n1307), .B2(new_n1288), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AND3_X1   g1110(.A1(new_n1224), .A2(KEYINPUT120), .A3(new_n1225), .ZN(new_n1311));
  AOI21_X1  g1111(.A(KEYINPUT120), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1261), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT57), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1264), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n736), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1231), .A2(new_n1258), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1315), .A2(new_n1318), .A3(new_n1202), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1230), .A2(new_n1070), .A3(new_n1261), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1226), .A2(new_n735), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1321), .B1(new_n1231), .B2(new_n1258), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1296), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1298), .B(new_n1310), .C1(new_n1319), .C2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT62), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1298), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n663), .A2(G213), .A3(G2897), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1328), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1307), .A2(new_n1288), .ZN(new_n1330));
  INV_X1    g1130(.A(G384), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1307), .A2(G384), .A3(new_n1288), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1327), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1329), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1326), .A2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT61), .ZN(new_n1337));
  OAI211_X1 g1137(.A(G378), .B(new_n1259), .C1(new_n1262), .C2(new_n1264), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1295), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1338), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT62), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1341), .A2(new_n1342), .A3(new_n1298), .A4(new_n1310), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1325), .A2(new_n1336), .A3(new_n1337), .A4(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(G393), .A2(G396), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1345), .A2(new_n1293), .ZN(new_n1346));
  OAI211_X1 g1146(.A(G390), .B(new_n1020), .C1(new_n1071), .C2(new_n1052), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(G387), .A2(new_n1137), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1346), .B1(new_n1349), .B2(KEYINPUT126), .ZN(new_n1350));
  AOI21_X1  g1150(.A(KEYINPUT126), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1346), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1350), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1344), .A2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT63), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1354), .B1(new_n1324), .B2(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(KEYINPUT61), .B1(new_n1326), .B2(new_n1335), .ZN(new_n1358));
  OAI211_X1 g1158(.A(new_n1357), .B(new_n1358), .C1(new_n1356), .C2(new_n1324), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1355), .A2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1362));
  AOI211_X1 g1162(.A(KEYINPUT126), .B(new_n1346), .C1(new_n1347), .C2(new_n1348), .ZN(new_n1363));
  OAI211_X1 g1163(.A(KEYINPUT127), .B(new_n1361), .C1(new_n1362), .C2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1361), .A2(KEYINPUT127), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1350), .A2(new_n1365), .A3(new_n1353), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1338), .B1(KEYINPUT127), .B2(new_n1361), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1368), .B1(G375), .B2(new_n1295), .ZN(new_n1369));
  XNOR2_X1  g1169(.A(new_n1367), .B(new_n1369), .ZN(G402));
endmodule


