//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n552,
    new_n554, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT68), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n459), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n459), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND3_X1  g049(.A1(new_n462), .A2(G2105), .A3(new_n464), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n466), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND3_X1   g057(.A1(new_n459), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n461), .B2(new_n460), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n484), .A2(new_n485), .A3(G126), .A4(G2105), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n462), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n459), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n491), .A2(KEYINPUT70), .A3(new_n492), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n468), .A2(G138), .A3(new_n463), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n466), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n489), .A2(KEYINPUT71), .A3(new_n497), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n486), .A2(new_n488), .A3(new_n497), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n500), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n465), .B2(new_n498), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n520), .A2(new_n522), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n514), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(new_n525), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n518), .A2(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(new_n524), .A2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n518), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n514), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n523), .B2(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n518), .A2(G43), .B1(G651), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n524), .A2(G81), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT73), .Z(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n518), .A2(G53), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n559), .A2(KEYINPUT76), .ZN(new_n561));
  AOI211_X1 g136(.A(new_n558), .B(new_n560), .C1(new_n561), .C2(KEYINPUT75), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n563));
  INV_X1    g138(.A(G78), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n523), .B(KEYINPUT77), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI221_X1 g141(.A(new_n563), .B1(new_n564), .B2(new_n517), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n523), .A2(KEYINPUT77), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n523), .A2(KEYINPUT77), .ZN(new_n569));
  NOR3_X1   g144(.A1(new_n568), .A2(new_n569), .A3(new_n566), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n564), .A2(new_n517), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT78), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n567), .A2(new_n572), .A3(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n524), .A2(G91), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n567), .A2(new_n572), .A3(new_n576), .A4(G651), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT75), .B(new_n558), .C1(new_n559), .C2(KEYINPUT76), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n574), .A2(new_n575), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n562), .A2(new_n579), .ZN(G299));
  NAND2_X1  g155(.A1(new_n518), .A2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n524), .A2(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n523), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n524), .A2(G86), .B1(G651), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  INV_X1    g164(.A(new_n518), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n524), .A2(G85), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n518), .A2(G47), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n514), .C2(new_n594), .ZN(G290));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NOR2_X1   g171(.A1(G171), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n524), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n603), .A2(G54), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n565), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g182(.A1(G79), .A2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n602), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n605), .A2(new_n602), .A3(new_n609), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n598), .B1(new_n613), .B2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(KEYINPUT80), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(KEYINPUT80), .B2(new_n597), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(KEYINPUT80), .B2(new_n597), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n562), .A2(new_n579), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n613), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n547), .A2(new_n548), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(new_n596), .ZN(new_n625));
  INV_X1    g200(.A(new_n612), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n600), .B1(new_n626), .B2(new_n610), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n627), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n625), .B1(new_n628), .B2(new_n596), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n476), .A2(G123), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n466), .A2(G135), .ZN(new_n632));
  NOR2_X1   g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n637), .B(new_n644), .C1(new_n642), .C2(new_n640), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2435), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2438), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2443), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1341), .B(G1348), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT86), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n656), .B(new_n658), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n663), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT87), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n662), .A3(new_n663), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  INV_X1    g246(.A(new_n664), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n662), .A3(new_n665), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(G2096), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT88), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(new_n641), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n680), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n681), .A2(new_n682), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n684), .A2(KEYINPUT20), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n688), .A2(new_n680), .A3(new_n683), .ZN(new_n689));
  OAI211_X1 g264(.A(new_n687), .B(new_n689), .C1(KEYINPUT20), .C2(new_n684), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT89), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n476), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n466), .A2(G131), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n463), .A2(G107), .ZN(new_n703));
  OR3_X1    g278(.A1(KEYINPUT90), .A2(G95), .A3(G2105), .ZN(new_n704));
  OAI21_X1  g279(.A(KEYINPUT90), .B1(G95), .B2(G2105), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n704), .A2(G2104), .A3(new_n705), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n700), .B1(new_n708), .B2(new_n699), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT35), .B(G1991), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G24), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G290), .B2(G16), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n712), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(G22), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G166), .B2(new_n714), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(G1971), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n714), .A2(G23), .ZN(new_n721));
  INV_X1    g296(.A(G288), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n714), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT33), .Z(new_n724));
  AOI21_X1  g299(.A(new_n720), .B1(new_n724), .B2(G1976), .ZN(new_n725));
  MUX2_X1   g300(.A(G6), .B(G305), .S(G16), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT32), .B(G1981), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n725), .B(new_n728), .C1(G1976), .C2(new_n724), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n717), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n730), .B2(new_n729), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n713), .B2(new_n716), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT36), .Z(new_n734));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n735));
  INV_X1    g310(.A(G26), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G29), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n476), .A2(G128), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n466), .A2(G140), .ZN(new_n740));
  NOR2_X1   g315(.A1(G104), .A2(G2105), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n738), .B1(new_n743), .B2(G29), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n737), .B1(new_n744), .B2(new_n735), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(G2067), .ZN(new_n746));
  NOR2_X1   g321(.A1(G29), .A2(G33), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n471), .A2(G103), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT25), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n463), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n749), .B(new_n751), .C1(G139), .C2(new_n466), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n747), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT92), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G2072), .ZN(new_n755));
  OR2_X1    g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  NAND2_X1  g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n756), .A2(new_n699), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G160), .B2(new_n699), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G2084), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT96), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n714), .A2(G5), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G171), .B2(new_n714), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n699), .B1(new_n766), .B2(G28), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(G28), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n635), .B2(new_n699), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n759), .B2(G2084), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n755), .A2(new_n761), .A3(new_n765), .A4(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G32), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n476), .A2(G129), .B1(G105), .B2(new_n471), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT26), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n466), .A2(G141), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT93), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n779), .B1(new_n785), .B2(G29), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT27), .B(G1996), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G27), .A2(G29), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G164), .B2(G29), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G2078), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT94), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G16), .B2(G21), .ZN(new_n793));
  NOR2_X1   g368(.A1(G286), .A2(new_n714), .ZN(new_n794));
  MUX2_X1   g369(.A(new_n793), .B(new_n792), .S(new_n794), .Z(new_n795));
  INV_X1    g370(.A(G1966), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n778), .A2(new_n788), .A3(new_n791), .A4(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(KEYINPUT97), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n714), .A2(G20), .ZN(new_n800));
  OAI211_X1 g375(.A(KEYINPUT23), .B(new_n800), .C1(new_n619), .C2(new_n714), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT23), .B2(new_n800), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n714), .A2(G4), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n613), .B2(new_n714), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(G1348), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n699), .A2(G35), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G162), .B2(new_n699), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT98), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT29), .ZN(new_n812));
  INV_X1    g387(.A(G2090), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n549), .A2(new_n714), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n714), .B2(G19), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G1341), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n817), .A2(G1341), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n814), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n807), .A2(G1348), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n812), .A2(new_n813), .B1(G2067), .B2(new_n745), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n808), .B(new_n823), .C1(new_n798), .C2(KEYINPUT97), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n734), .A2(new_n746), .A3(new_n805), .A4(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  NAND2_X1  g401(.A1(G80), .A2(G543), .ZN(new_n827));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n523), .B2(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n518), .A2(G55), .B1(G651), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n524), .A2(G93), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT100), .B(G860), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n613), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n549), .A2(new_n832), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n624), .A2(new_n831), .A3(new_n830), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n835), .B1(new_n843), .B2(new_n833), .ZN(G145));
  XNOR2_X1  g419(.A(new_n785), .B(new_n743), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n505), .A2(KEYINPUT101), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n486), .A2(new_n488), .A3(new_n848), .A4(new_n497), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n846), .B1(new_n850), .B2(new_n502), .ZN(new_n851));
  AOI211_X1 g426(.A(KEYINPUT102), .B(new_n507), .C1(new_n847), .C2(new_n849), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n845), .B(new_n853), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n752), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n466), .A2(G142), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n856), .A2(KEYINPUT103), .B1(G130), .B2(new_n476), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n463), .A2(G118), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n459), .B1(new_n858), .B2(KEYINPUT104), .ZN(new_n859));
  OAI221_X1 g434(.A(new_n859), .B1(KEYINPUT104), .B2(new_n858), .C1(G106), .C2(G2105), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n860), .C1(KEYINPUT103), .C2(new_n856), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n639), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n707), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT105), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n855), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n635), .B(new_n473), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n481), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n855), .B2(new_n863), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n864), .B2(new_n855), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g447(.A1(new_n832), .A2(new_n596), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n628), .B(new_n840), .ZN(new_n874));
  NAND2_X1  g449(.A1(G299), .A2(new_n613), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n627), .A2(new_n619), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n878), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G288), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(G166), .B(G305), .ZN(new_n890));
  MUX2_X1   g465(.A(new_n887), .B(new_n889), .S(new_n890), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n884), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n873), .B1(new_n892), .B2(new_n596), .ZN(G295));
  OAI21_X1  g468(.A(new_n873), .B1(new_n892), .B2(new_n596), .ZN(G331));
  NAND2_X1  g469(.A1(new_n840), .A2(G171), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n840), .A2(G171), .ZN(new_n897));
  OAI21_X1  g472(.A(G286), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n897), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(G168), .A3(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n880), .B2(new_n881), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n898), .A2(new_n900), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n877), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n904), .A3(new_n891), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT109), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n902), .A2(new_n904), .A3(new_n907), .A4(new_n891), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n906), .B2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n891), .B(KEYINPUT108), .Z(new_n910));
  NOR2_X1   g485(.A1(new_n877), .A2(KEYINPUT41), .ZN(new_n911));
  AOI211_X1 g486(.A(new_n903), .B(new_n911), .C1(new_n877), .C2(new_n879), .ZN(new_n912));
  INV_X1    g487(.A(new_n904), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n914), .A3(KEYINPUT43), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n902), .A2(new_n904), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT43), .B1(new_n909), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n909), .A2(new_n914), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n922), .B1(new_n909), .B2(new_n918), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n920), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n920), .B2(new_n926), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(G397));
  XNOR2_X1  g505(.A(new_n785), .B(G1996), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n743), .B(G2067), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT111), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(new_n711), .B2(new_n708), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n711), .B2(new_n708), .ZN(new_n936));
  NOR2_X1   g511(.A1(G290), .A2(G1986), .ZN(new_n937));
  AND2_X1   g512(.A1(G290), .A2(G1986), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n853), .B2(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(G160), .A2(G40), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT54), .ZN(new_n947));
  INV_X1    g522(.A(G1384), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT45), .B(new_n948), .C1(new_n851), .C2(new_n852), .ZN(new_n949));
  INV_X1    g524(.A(G2078), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n503), .A2(new_n508), .A3(new_n948), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n942), .B1(new_n951), .B2(new_n940), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT124), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n951), .A2(KEYINPUT50), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT112), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n951), .A2(new_n959), .A3(KEYINPUT50), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n942), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G1384), .B1(new_n850), .B2(new_n502), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G1961), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n955), .A2(new_n956), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n507), .B1(new_n847), .B2(new_n849), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n940), .B1(new_n967), .B2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n969));
  INV_X1    g544(.A(new_n942), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n969), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n951), .A2(new_n940), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n954), .A2(G2078), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(G301), .B1(new_n966), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n953), .A2(new_n954), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT124), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n954), .ZN(new_n981));
  INV_X1    g556(.A(new_n960), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n959), .B1(new_n951), .B2(KEYINPUT50), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n970), .B(new_n964), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n764), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n941), .A2(new_n949), .A3(new_n970), .A4(new_n975), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n980), .A2(new_n981), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(G171), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n947), .B1(new_n977), .B2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n980), .A2(new_n976), .A3(new_n985), .A4(new_n981), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT125), .B1(new_n990), .B2(G171), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT125), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n966), .A2(new_n992), .A3(G301), .A4(new_n976), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n947), .B1(new_n987), .B2(G171), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n958), .A2(new_n960), .ZN(new_n996));
  INV_X1    g571(.A(G2084), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n970), .A4(new_n964), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n998), .B1(new_n974), .B2(G1966), .ZN(new_n999));
  NAND2_X1  g574(.A1(G286), .A2(G8), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(G8), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n1000), .B(KEYINPUT123), .Z(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G8), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n968), .A2(new_n970), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT117), .ZN(new_n1009));
  INV_X1    g584(.A(new_n973), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n796), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1007), .B1(new_n1013), .B2(new_n998), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1001), .A2(KEYINPUT51), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1002), .B1(new_n1006), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n949), .A2(new_n952), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(G2090), .B2(new_n984), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G303), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT113), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1022), .B(G8), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G288), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT114), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n962), .A2(new_n970), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1030), .A2(KEYINPUT114), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1031), .A2(G8), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n722), .A2(G1976), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n1034), .A2(KEYINPUT52), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G305), .A2(G1981), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n588), .B(new_n1039), .C1(new_n589), .C2(new_n590), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1043), .A2(G8), .A3(new_n1032), .A4(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1036), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1027), .A2(new_n1025), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT50), .B1(new_n967), .B2(G1384), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(new_n970), .C1(KEYINPUT50), .C2(new_n951), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1051), .B2(new_n1007), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1028), .A2(new_n1046), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n989), .A2(new_n995), .A3(new_n1018), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT126), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT120), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1032), .B(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2067), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1348), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n984), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT60), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1057), .B1(new_n1066), .B2(new_n613), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT60), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1068), .A2(KEYINPUT121), .A3(new_n627), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1067), .A2(new_n1069), .B1(new_n1065), .B2(new_n1064), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n574), .A2(new_n1071), .A3(new_n575), .A4(new_n577), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n619), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1073), .B(new_n1072), .C1(new_n562), .C2(new_n579), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1049), .A2(new_n803), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT56), .B(G2072), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n949), .A2(new_n952), .A3(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1082), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n1084), .B(KEYINPUT61), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1066), .A2(new_n1057), .A3(new_n613), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT121), .B1(new_n1068), .B2(new_n627), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1064), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(KEYINPUT60), .A4(new_n1088), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT58), .B(G1341), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n1059), .A2(new_n1090), .B1(new_n1019), .B2(G1996), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n549), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT59), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1070), .A2(new_n1085), .A3(new_n1089), .A4(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1083), .B1(new_n1088), .B2(new_n627), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1081), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1002), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1003), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1005), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1014), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1004), .A2(new_n1015), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1098), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(new_n1053), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(new_n1105), .A3(new_n989), .A4(new_n995), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1056), .A2(new_n1097), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1045), .A2(new_n1029), .A3(new_n722), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1040), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT115), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1032), .A2(G8), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1109), .A2(new_n1114), .A3(new_n1040), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1036), .A2(new_n1037), .A3(new_n1045), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1028), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1108), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1120));
  OAI221_X1 g695(.A(KEYINPUT116), .B1(new_n1028), .B2(new_n1117), .C1(new_n1120), .C2(new_n1112), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(KEYINPUT118), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1014), .A2(G168), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1124), .B(new_n1125), .C1(new_n1053), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1022), .A2(G8), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1123), .B1(new_n1129), .B2(new_n1047), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1128), .A2(new_n1130), .A3(new_n1028), .A4(new_n1046), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1054), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT62), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n977), .B1(new_n1103), .B2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1122), .B(new_n1132), .C1(new_n1133), .C2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n946), .B1(new_n1107), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n944), .A2(G1996), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT46), .Z(new_n1139));
  AND2_X1   g714(.A1(new_n933), .A2(new_n785), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1139), .B1(new_n944), .B2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT47), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n936), .A2(new_n943), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n943), .A2(new_n937), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT48), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1144), .A2(KEYINPUT48), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1143), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n934), .A2(new_n710), .A3(new_n707), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n743), .A2(G2067), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n943), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1142), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1137), .A2(KEYINPUT127), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1056), .A2(new_n1097), .A3(new_n1106), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1136), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n945), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1154), .B1(new_n1157), .B2(new_n1151), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1153), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g734(.A1(G319), .A2(new_n871), .A3(new_n660), .A4(new_n677), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n909), .A2(new_n918), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n1162), .A2(KEYINPUT43), .ZN(new_n1163));
  NAND2_X1  g737(.A1(new_n1163), .A2(new_n923), .ZN(new_n1164));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n697), .A3(new_n1164), .ZN(G225));
  INV_X1    g739(.A(G225), .ZN(G308));
endmodule


