//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G20), .ZN(new_n214));
  AND2_X1   g0014(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n219), .A2(G50), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  INV_X1    g0027(.A(G250), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n230));
  INV_X1    g0030(.A(G77), .ZN(new_n231));
  INV_X1    g0031(.A(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G107), .ZN(new_n233));
  INV_X1    g0033(.A(G264), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n230), .B1(new_n231), .B2(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n207), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  INV_X1    g0037(.A(KEYINPUT1), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT68), .ZN(new_n240));
  AOI211_X1 g0040(.A(new_n223), .B(new_n240), .C1(new_n238), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  INV_X1    g0042(.A(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(KEYINPUT2), .B(G226), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G358));
  XNOR2_X1  g0050(.A(G50), .B(G68), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G58), .B(G77), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n251), .B(new_n252), .Z(new_n253));
  XOR2_X1   g0053(.A(G87), .B(G97), .Z(new_n254));
  XOR2_X1   g0054(.A(G107), .B(G116), .Z(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n253), .B(new_n256), .Z(G351));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n216), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n215), .A2(G33), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n263));
  INV_X1    g0063(.A(G150), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n259), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(new_n259), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n211), .A2(G1), .ZN(new_n273));
  INV_X1    g0073(.A(G50), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n272), .A2(new_n275), .B1(new_n274), .B2(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n268), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT9), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(G1), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n280), .A2(G274), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  NOR3_X1   g0085(.A1(new_n279), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT3), .B(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(G222), .ZN(new_n291));
  INV_X1    g0091(.A(G223), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(G1698), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n291), .B1(new_n231), .B2(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n284), .B(new_n286), .C1(new_n294), .C2(new_n279), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G190), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n278), .B(new_n296), .C1(new_n297), .C2(new_n295), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n277), .C1(G169), .C2(new_n295), .ZN(new_n302));
  XOR2_X1   g0102(.A(new_n302), .B(KEYINPUT70), .Z(new_n303));
  XOR2_X1   g0103(.A(KEYINPUT15), .B(G87), .Z(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n260), .A2(new_n305), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n215), .A2(new_n231), .B1(new_n266), .B2(new_n261), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n259), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n272), .ZN(new_n309));
  OAI21_X1  g0109(.A(G77), .B1(new_n211), .B2(G1), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n308), .B1(G77), .B2(new_n270), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n279), .A2(new_n283), .A3(new_n232), .ZN(new_n312));
  INV_X1    g0112(.A(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G107), .ZN(new_n318));
  OR2_X1    g0118(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n319));
  NAND2_X1  g0119(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n319), .A2(new_n314), .A3(new_n316), .A4(new_n320), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n318), .B1(new_n321), .B2(new_n243), .C1(new_n226), .C2(new_n293), .ZN(new_n322));
  AOI211_X1 g0122(.A(new_n284), .B(new_n312), .C1(new_n322), .C2(new_n279), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n297), .ZN(new_n324));
  AOI211_X1 g0124(.A(new_n311), .B(new_n324), .C1(G190), .C2(new_n323), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n311), .B1(new_n323), .B2(G169), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n323), .A2(new_n300), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n299), .A2(new_n303), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n261), .A2(new_n273), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n272), .B1(new_n271), .B2(new_n261), .ZN(new_n332));
  INV_X1    g0132(.A(G58), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(new_n225), .ZN(new_n334));
  OAI21_X1  g0134(.A(G20), .B1(new_n334), .B2(new_n201), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n265), .A2(G159), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n317), .A2(new_n211), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n225), .B1(new_n338), .B2(KEYINPUT7), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n215), .A2(new_n340), .A3(new_n317), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n337), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n259), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n212), .A2(new_n214), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(new_n340), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT73), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n314), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n313), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n348), .A2(new_n316), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT7), .B1(new_n317), .B2(new_n211), .ZN(new_n352));
  OAI21_X1  g0152(.A(G68), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n337), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT16), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n332), .B1(new_n344), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT76), .ZN(new_n357));
  INV_X1    g0157(.A(G274), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n279), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n283), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n279), .A2(new_n283), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G232), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n314), .A2(new_n316), .A3(G226), .A4(G1698), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n364), .B(new_n365), .C1(new_n321), .C2(new_n292), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n280), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n289), .A2(new_n290), .A3(G223), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n369), .A2(KEYINPUT74), .A3(new_n364), .A4(new_n365), .ZN(new_n370));
  AOI211_X1 g0170(.A(G190), .B(new_n363), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n289), .A2(new_n290), .A3(G223), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n364), .A2(new_n365), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n367), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n374), .A2(new_n370), .A3(new_n279), .ZN(new_n375));
  INV_X1    g0175(.A(new_n363), .ZN(new_n376));
  AOI21_X1  g0176(.A(G200), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n357), .B1(new_n371), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G190), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n375), .A2(new_n379), .A3(new_n376), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n363), .B1(new_n368), .B2(new_n370), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(KEYINPUT76), .C1(G200), .C2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n356), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT17), .ZN(new_n384));
  AOI211_X1 g0184(.A(G179), .B(new_n363), .C1(new_n368), .C2(new_n370), .ZN(new_n385));
  AOI21_X1  g0185(.A(G169), .B1(new_n375), .B2(new_n376), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT75), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n375), .A2(new_n300), .A3(new_n376), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n388), .B(new_n389), .C1(G169), .C2(new_n381), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n356), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT18), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n387), .A2(new_n356), .A3(new_n390), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n265), .A2(G50), .B1(G20), .B2(new_n225), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n260), .B2(new_n231), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n259), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT11), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n309), .A2(new_n225), .A3(new_n273), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n271), .A2(new_n225), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT12), .B1(new_n402), .B2(KEYINPUT72), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(KEYINPUT72), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(KEYINPUT72), .A3(KEYINPUT12), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n284), .B1(G238), .B2(new_n361), .ZN(new_n409));
  INV_X1    g0209(.A(G97), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n321), .A2(new_n285), .B1(new_n313), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT71), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n293), .B2(new_n243), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n290), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n409), .B1(new_n415), .B2(new_n280), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT13), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT13), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n409), .B(new_n418), .C1(new_n415), .C2(new_n280), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(G169), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n300), .B2(new_n420), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n420), .B2(G169), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n408), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n407), .B(new_n400), .C1(new_n420), .C2(new_n379), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n297), .B1(new_n417), .B2(new_n419), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n330), .A2(new_n396), .A3(new_n425), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n259), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT19), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n433), .A2(new_n313), .A3(new_n410), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n434), .A2(new_n345), .B1(G87), .B2(new_n205), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n215), .A2(G68), .A3(new_n290), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n212), .A2(new_n214), .A3(G33), .A4(G97), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n433), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT82), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT82), .A4(new_n438), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n441), .A2(new_n442), .B1(new_n271), .B2(new_n305), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n269), .A2(G33), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n270), .A2(new_n444), .A3(new_n216), .A4(new_n258), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G87), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n282), .A2(G1), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n358), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n228), .B1(new_n282), .B2(G1), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n280), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT79), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n321), .B2(new_n226), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT79), .A4(G238), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G116), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n314), .A2(new_n316), .A3(G244), .A4(G1698), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n454), .B1(new_n460), .B2(new_n279), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G190), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n462), .A2(KEYINPUT83), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n279), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n453), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G200), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(KEYINPUT83), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n449), .A2(new_n463), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(G169), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n459), .A2(new_n458), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n289), .A2(new_n290), .A3(G238), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n471), .B1(new_n455), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n280), .B1(new_n473), .B2(new_n457), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n470), .B1(new_n474), .B2(new_n454), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n461), .A2(new_n300), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g0277(.A(G179), .B(new_n454), .C1(new_n460), .C2(new_n279), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(KEYINPUT80), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT81), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n461), .A2(G169), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT80), .B1(new_n481), .B2(new_n478), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n476), .A2(new_n469), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n441), .A2(new_n442), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n305), .A2(new_n271), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n446), .A2(new_n304), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT4), .A4(G244), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT77), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n321), .B2(new_n232), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n290), .A2(G250), .A3(G1698), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n280), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n269), .B(G45), .C1(new_n281), .C2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT78), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n500), .A2(new_n501), .B1(KEYINPUT5), .B2(new_n281), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n450), .B(KEYINPUT78), .C1(KEYINPUT5), .C2(new_n281), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n279), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G257), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n500), .A2(new_n501), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n359), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  OR3_X1    g0310(.A1(new_n499), .A2(G179), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n270), .A2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n445), .B2(new_n410), .ZN(new_n514));
  OAI21_X1  g0314(.A(G107), .B1(new_n351), .B2(new_n352), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n233), .A2(KEYINPUT6), .A3(G97), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n410), .A2(new_n233), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n204), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(KEYINPUT6), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n345), .B1(G77), .B2(new_n265), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n514), .B1(new_n521), .B2(new_n259), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n470), .B1(new_n499), .B2(new_n510), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n511), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n290), .A2(G257), .A3(G1698), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G294), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n228), .C2(new_n321), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n279), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n502), .A2(new_n503), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G264), .A3(new_n280), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n509), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n297), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n279), .A2(new_n528), .B1(new_n504), .B2(G264), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n379), .A3(new_n509), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT85), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n212), .A2(new_n214), .A3(new_n314), .A4(new_n316), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT22), .B1(new_n537), .B2(new_n227), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n215), .A2(new_n539), .A3(G87), .A4(new_n290), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND2_X1  g0342(.A1(KEYINPUT23), .A2(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n544), .B2(G20), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT23), .A2(G107), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n345), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n542), .B1(new_n541), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n259), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n271), .A2(KEYINPUT25), .A3(new_n233), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT25), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n270), .B2(G107), .ZN(new_n553));
  AOI22_X1  g0353(.A1(G107), .A2(new_n446), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT85), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n534), .A2(new_n555), .A3(new_n379), .A4(new_n509), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n536), .A2(new_n550), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(G200), .B1(new_n499), .B2(new_n510), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n491), .A2(new_n492), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n491), .A2(new_n492), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n509), .B(new_n505), .C1(new_n562), .C2(new_n280), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n558), .B(new_n522), .C1(new_n563), .C2(new_n379), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n525), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n289), .A2(new_n290), .A3(G257), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n317), .A2(G303), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n293), .A2(new_n234), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n279), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n504), .A2(G270), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n571), .A2(new_n572), .A3(new_n509), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n313), .A2(G97), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n212), .A2(new_n214), .A3(new_n574), .A4(new_n496), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  AOI22_X1  g0377(.A1(KEYINPUT84), .A2(new_n576), .B1(new_n577), .B2(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n259), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT84), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n270), .A2(new_n577), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n446), .B2(new_n577), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(KEYINPUT20), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n575), .A2(new_n259), .A3(new_n578), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G169), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n566), .B1(new_n573), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(G270), .A2(new_n504), .B1(new_n508), .B2(new_n359), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n589), .A2(new_n586), .A3(G179), .A4(new_n571), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n571), .A2(new_n572), .A3(new_n509), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n591), .A2(KEYINPUT21), .A3(G169), .A4(new_n586), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n550), .A2(new_n554), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n532), .A2(new_n470), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n529), .A2(new_n509), .A3(new_n531), .A4(new_n300), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n586), .B1(new_n591), .B2(G200), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n379), .B2(new_n591), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n593), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n565), .A2(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n431), .A2(new_n468), .A3(new_n490), .A4(new_n601), .ZN(G372));
  INV_X1    g0402(.A(KEYINPUT87), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n395), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n392), .A2(KEYINPUT87), .A3(new_n394), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n424), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(new_n422), .C1(new_n300), .C2(new_n420), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n408), .A2(new_n608), .B1(new_n429), .B2(new_n328), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n606), .B1(new_n609), .B2(new_n384), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n299), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n303), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n525), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n490), .A2(new_n468), .A3(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n615), .A2(KEYINPUT26), .ZN(new_n616));
  INV_X1    g0416(.A(new_n565), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n489), .A2(new_n476), .A3(new_n475), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n466), .A2(new_n447), .A3(new_n443), .A4(new_n462), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT86), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n593), .A2(new_n597), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n595), .A2(new_n596), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n623), .B1(new_n550), .B2(new_n554), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT86), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n617), .A2(new_n620), .A3(new_n622), .A4(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n522), .B1(new_n563), .B2(new_n470), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n628), .A2(new_n511), .A3(new_n618), .A4(new_n619), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n618), .B1(new_n629), .B2(KEYINPUT26), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n431), .B1(new_n616), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n613), .A2(new_n633), .ZN(G369));
  NAND3_X1  g0434(.A1(new_n215), .A2(new_n269), .A3(G13), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(KEYINPUT27), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g0438(.A(KEYINPUT88), .B(G343), .Z(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n586), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n593), .A2(new_n599), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n593), .B2(new_n641), .ZN(new_n643));
  XOR2_X1   g0443(.A(new_n643), .B(KEYINPUT89), .Z(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G330), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n594), .A2(new_n640), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n624), .B1(new_n557), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n597), .A2(new_n640), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n640), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n625), .A2(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n649), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n618), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n525), .A2(new_n564), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT92), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n620), .A2(new_n557), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n597), .B2(new_n593), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT91), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n615), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n614), .A2(new_n620), .A3(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n663), .B1(new_n615), .B2(new_n664), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(KEYINPUT29), .A3(new_n652), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n652), .B1(new_n632), .B2(new_n616), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT29), .ZN(new_n672));
  AOI21_X1  g0472(.A(KEYINPUT93), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n615), .A2(new_n664), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT91), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n666), .A3(new_n665), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n640), .B1(new_n677), .B2(new_n662), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(KEYINPUT93), .A3(KEYINPUT29), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n601), .A2(new_n468), .A3(new_n490), .A4(new_n652), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n573), .A2(G179), .A3(new_n461), .A4(new_n534), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT90), .B1(new_n683), .B2(new_n563), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT30), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT90), .B(new_n686), .C1(new_n683), .C2(new_n563), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n461), .A2(G179), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n563), .A2(new_n532), .A3(new_n591), .A4(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(KEYINPUT31), .B1(new_n690), .B2(new_n640), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n640), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n682), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n681), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n269), .ZN(new_n697));
  INV_X1    g0497(.A(new_n208), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n221), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n697), .A2(new_n704), .ZN(G364));
  NAND2_X1  g0505(.A1(new_n215), .A2(G13), .ZN(new_n706));
  XOR2_X1   g0506(.A(new_n706), .B(KEYINPUT94), .Z(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G45), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G1), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n699), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n646), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G330), .B2(new_n644), .ZN(new_n712));
  INV_X1    g0512(.A(G355), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n290), .A2(new_n208), .ZN(new_n714));
  OAI22_X1  g0514(.A1(new_n713), .A2(new_n714), .B1(G116), .B2(new_n208), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n253), .A2(new_n282), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT95), .Z(new_n717));
  NOR2_X1   g0517(.A1(new_n698), .A2(new_n290), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n221), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n719), .B1(new_n720), .B2(new_n282), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n715), .B1(new_n717), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G13), .A2(G33), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n216), .B1(G20), .B2(new_n470), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n710), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G303), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n297), .A2(G179), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(G20), .A3(G190), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n300), .A2(new_n297), .A3(G190), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n345), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G294), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n317), .B1(new_n730), .B2(new_n732), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n345), .A2(G179), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(new_n379), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G326), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n737), .A2(G190), .ZN(new_n742));
  XNOR2_X1  g0542(.A(KEYINPUT33), .B(G317), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n736), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n345), .A2(new_n379), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT97), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(G179), .A3(new_n297), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n747), .A2(G179), .A3(G200), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G283), .A2(new_n748), .B1(new_n749), .B2(G329), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n345), .A2(G179), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n752));
  AOI21_X1  g0552(.A(G200), .B1(new_n751), .B2(KEYINPUT96), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n379), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(G190), .A3(new_n753), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(G311), .A2(new_n755), .B1(new_n757), .B2(G322), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n744), .A2(new_n750), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n734), .B(KEYINPUT99), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G97), .ZN(new_n761));
  INV_X1    g0561(.A(new_n742), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n761), .B1(new_n762), .B2(new_n225), .C1(new_n274), .C2(new_n739), .ZN(new_n763));
  INV_X1    g0563(.A(new_n749), .ZN(new_n764));
  INV_X1    g0564(.A(G159), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n767), .B2(KEYINPUT32), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT32), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n766), .A2(new_n769), .B1(G58), .B2(new_n757), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n768), .B(new_n770), .C1(new_n231), .C2(new_n754), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n748), .A2(G107), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n772), .B(new_n290), .C1(new_n227), .C2(new_n732), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT98), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n759), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n729), .B1(new_n775), .B2(new_n726), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n725), .B(KEYINPUT100), .Z(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n643), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n712), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(G396));
  NAND2_X1  g0580(.A1(new_n311), .A2(new_n640), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT102), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n325), .A2(new_n782), .B1(new_n327), .B2(new_n326), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n328), .A2(new_n652), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n671), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n785), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n652), .B(new_n787), .C1(new_n632), .C2(new_n616), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(KEYINPUT103), .B1(new_n790), .B2(new_n695), .ZN(new_n791));
  INV_X1    g0591(.A(new_n710), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT103), .ZN(new_n793));
  INV_X1    g0593(.A(G330), .ZN(new_n794));
  INV_X1    g0594(.A(new_n693), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n691), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n794), .B1(new_n796), .B2(new_n682), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n789), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n791), .A2(new_n792), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT104), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(KEYINPUT104), .B1(new_n695), .B2(new_n790), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n726), .A2(new_n723), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n792), .B1(new_n231), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G87), .A2(new_n748), .B1(new_n749), .B2(G311), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n317), .B1(new_n732), .B2(new_n233), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n760), .B2(G97), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G116), .A2(new_n755), .B1(new_n757), .B2(G294), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G283), .A2(new_n742), .B1(new_n738), .B2(G303), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n805), .A2(new_n807), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n290), .B1(new_n274), .B2(new_n732), .C1(new_n734), .C2(new_n333), .ZN(new_n811));
  INV_X1    g0611(.A(new_n748), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n225), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n811), .B(new_n813), .C1(G132), .C2(new_n749), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G137), .A2(new_n738), .B1(new_n742), .B2(G150), .ZN(new_n815));
  INV_X1    g0615(.A(G143), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n754), .B2(new_n765), .C1(new_n816), .C2(new_n756), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(KEYINPUT34), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT34), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n810), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT101), .Z(new_n823));
  INV_X1    g0623(.A(new_n726), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n804), .B1(new_n724), .B2(new_n787), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n802), .A2(new_n825), .ZN(G384));
  OR2_X1    g0626(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n827), .A2(G116), .A3(new_n217), .A4(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT36), .Z(new_n830));
  OR3_X1    g0630(.A1(new_n221), .A2(new_n231), .A3(new_n334), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n274), .A2(G68), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n269), .B(G13), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n608), .A2(new_n408), .A3(new_n652), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT38), .ZN(new_n837));
  INV_X1    g0637(.A(new_n638), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n356), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT17), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n383), .B(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n606), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n378), .A2(new_n382), .ZN(new_n843));
  INV_X1    g0643(.A(new_n356), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n845), .A2(new_n846), .A3(new_n391), .A4(new_n839), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT107), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n391), .A2(new_n839), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT37), .B1(new_n849), .B2(new_n383), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n847), .A2(KEYINPUT107), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n837), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n342), .A2(KEYINPUT16), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n332), .B1(new_n344), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n838), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n384), .B2(new_n395), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n387), .A2(new_n390), .A3(new_n856), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n383), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n858), .B1(new_n861), .B2(KEYINPUT105), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT105), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n860), .B2(new_n383), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n846), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n847), .ZN(new_n866));
  OAI211_X1 g0666(.A(KEYINPUT38), .B(new_n859), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT39), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n387), .A2(new_n390), .A3(new_n856), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n845), .A2(KEYINPUT105), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n864), .A2(new_n871), .A3(new_n857), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n866), .B1(new_n872), .B2(KEYINPUT37), .ZN(new_n873));
  INV_X1    g0673(.A(new_n395), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n857), .B1(new_n841), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n837), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT106), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n867), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT106), .B(new_n837), .C1(new_n873), .C2(new_n875), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n836), .B(new_n869), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n408), .B(new_n640), .C1(new_n608), .C2(new_n428), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n408), .A2(new_n640), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n425), .A2(new_n429), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n788), .B2(new_n784), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n878), .A2(new_n888), .A3(new_n879), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n604), .A2(new_n605), .A3(new_n638), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n612), .B1(new_n680), .B2(new_n431), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n694), .A2(new_n787), .A3(new_n886), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n878), .A2(new_n879), .A3(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT40), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n854), .A2(new_n867), .ZN(new_n900));
  AND4_X1   g0700(.A1(KEYINPUT40), .A2(new_n694), .A3(new_n787), .A4(new_n886), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n431), .A2(new_n694), .ZN(new_n904));
  OAI21_X1  g0704(.A(G330), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n895), .A2(new_n906), .B1(new_n269), .B2(new_n707), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n895), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n834), .B1(new_n907), .B2(new_n908), .ZN(G367));
  OAI221_X1 g0709(.A(new_n727), .B1(new_n208), .B2(new_n305), .C1(new_n249), .C2(new_n719), .ZN(new_n910));
  INV_X1    g0710(.A(new_n732), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(G116), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT46), .Z(new_n913));
  INV_X1    g0713(.A(new_n734), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n290), .B(new_n913), .C1(G107), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n738), .A2(G311), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(new_n735), .C2(new_n762), .ZN(new_n917));
  INV_X1    g0717(.A(G317), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n410), .A2(new_n812), .B1(new_n764), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(G283), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n920), .A2(new_n754), .B1(new_n756), .B2(new_n730), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n917), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n812), .A2(new_n231), .ZN(new_n923));
  XOR2_X1   g0723(.A(KEYINPUT109), .B(G137), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n764), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n760), .A2(G68), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n738), .A2(G143), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n742), .A2(G159), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n317), .B1(new_n911), .B2(G58), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n923), .A2(new_n925), .A3(new_n930), .ZN(new_n931));
  AOI22_X1  g0731(.A1(G50), .A2(new_n755), .B1(new_n757), .B2(G150), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n922), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n710), .B(new_n910), .C1(new_n934), .C2(new_n824), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT110), .Z(new_n936));
  OAI21_X1  g0736(.A(new_n620), .B1(new_n449), .B2(new_n652), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n657), .A2(new_n448), .A3(new_n640), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n936), .B1(new_n777), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n525), .A2(new_n652), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n523), .A2(new_n640), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n941), .B1(new_n659), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n654), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT42), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n659), .A2(new_n624), .A3(new_n942), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n525), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n652), .ZN(new_n950));
  INV_X1    g0750(.A(new_n939), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(KEYINPUT108), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT108), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT43), .B1(new_n939), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n947), .A2(new_n950), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n947), .A2(new_n950), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n954), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n958), .B2(new_n951), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n955), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n651), .A2(new_n943), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n960), .B(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n944), .B2(new_n655), .ZN(new_n965));
  INV_X1    g0765(.A(new_n655), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(new_n943), .A3(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n944), .A2(KEYINPUT45), .A3(new_n655), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n966), .B2(new_n943), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n651), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n651), .A2(new_n968), .A3(new_n972), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n650), .B(new_n653), .Z(new_n978));
  XNOR2_X1  g0778(.A(new_n645), .B(new_n978), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n695), .B(new_n681), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n699), .B(KEYINPUT41), .Z(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n709), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n940), .B1(new_n963), .B2(new_n983), .ZN(G387));
  NAND2_X1  g0784(.A1(new_n696), .A2(new_n979), .ZN(new_n985));
  INV_X1    g0785(.A(new_n979), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n986), .A2(new_n695), .A3(new_n674), .A4(new_n679), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n699), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n246), .A2(G45), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT111), .ZN(new_n990));
  INV_X1    g0790(.A(new_n261), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n274), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT50), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n701), .B(new_n282), .C1(new_n225), .C2(new_n231), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n990), .B(new_n718), .C1(new_n993), .C2(new_n994), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(G107), .B2(new_n208), .C1(new_n701), .C2(new_n714), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n792), .B1(new_n996), .B2(new_n727), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n650), .B2(new_n777), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G311), .A2(new_n742), .B1(new_n738), .B2(G322), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n754), .B2(new_n730), .C1(new_n918), .C2(new_n756), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT113), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT48), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT48), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n914), .A2(G283), .B1(G294), .B2(new_n911), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT49), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n317), .B1(new_n812), .B2(new_n577), .C1(new_n740), .C2(new_n764), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(KEYINPUT49), .B2(new_n1007), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(KEYINPUT112), .B(G150), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G97), .A2(new_n748), .B1(new_n749), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n760), .A2(new_n304), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n317), .B1(new_n911), .B2(G77), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G159), .A2(new_n738), .B1(new_n742), .B2(new_n991), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1013), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n274), .A2(new_n756), .B1(new_n754), .B2(new_n225), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1011), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n998), .B1(new_n1020), .B2(new_n726), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n709), .B2(new_n986), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n988), .A2(new_n1022), .ZN(G393));
  INV_X1    g0823(.A(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n987), .A2(new_n977), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n699), .B1(new_n987), .B2(new_n977), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1024), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n987), .A2(new_n977), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1029), .A2(new_n1025), .A3(KEYINPUT117), .A4(new_n699), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n977), .A2(KEYINPUT114), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n709), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n977), .B2(KEYINPUT114), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n943), .A2(new_n725), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n749), .A2(G322), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n317), .B1(new_n920), .B2(new_n732), .C1(new_n734), .C2(new_n577), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G303), .B2(new_n742), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n772), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n757), .A2(G311), .B1(G317), .B2(new_n738), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT52), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(G294), .C2(new_n755), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT116), .Z(new_n1042));
  OAI22_X1  g0842(.A1(new_n227), .A2(new_n812), .B1(new_n764), .B2(new_n816), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n760), .A2(G77), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n317), .B1(new_n911), .B2(G68), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n274), .C2(new_n762), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n756), .A2(new_n765), .B1(new_n264), .B2(new_n739), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(new_n261), .C2(new_n754), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT115), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n824), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n727), .B1(new_n410), .B2(new_n208), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n256), .B2(new_n718), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1052), .A2(new_n792), .A3(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1031), .A2(new_n1033), .B1(new_n1034), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1028), .A2(new_n1030), .A3(new_n1056), .ZN(G390));
  AOI21_X1  g0857(.A(new_n881), .B1(new_n878), .B2(new_n879), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1058), .A2(new_n868), .B1(new_n836), .B2(new_n888), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n678), .A2(new_n783), .B1(new_n328), .B2(new_n652), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n835), .B(new_n900), .C1(new_n1060), .C2(new_n887), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AND4_X1   g0862(.A1(G330), .A2(new_n694), .A3(new_n787), .A4(new_n886), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n788), .A2(new_n784), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n886), .B1(new_n797), .B2(new_n787), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1065), .B1(new_n1066), .B2(new_n1063), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n887), .B1(new_n695), .B2(new_n785), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n797), .A2(new_n787), .A3(new_n886), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n669), .A2(new_n652), .A3(new_n783), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n784), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT93), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n626), .A2(new_n622), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n618), .A2(new_n619), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n565), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n630), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n615), .A2(KEYINPUT26), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n640), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1079), .B2(KEYINPUT29), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(new_n678), .B2(KEYINPUT29), .ZN(new_n1081));
  AND4_X1   g0881(.A1(KEYINPUT93), .A2(new_n669), .A3(KEYINPUT29), .A4(new_n652), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n431), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n431), .A2(new_n797), .ZN(new_n1084));
  AND4_X1   g0884(.A1(new_n613), .A2(new_n1072), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1059), .A2(new_n1061), .A3(new_n1069), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1064), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n894), .A2(new_n1084), .A3(new_n1072), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n1059), .A2(new_n1061), .A3(new_n1069), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1069), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1087), .A2(new_n1091), .A3(new_n699), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1058), .A2(new_n868), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n724), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n803), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n813), .B1(G294), .B2(new_n749), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n317), .B1(new_n227), .B2(new_n732), .C1(new_n739), .C2(new_n920), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G107), .B2(new_n742), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G97), .B2(new_n755), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1044), .B1(new_n577), .B2(new_n756), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT118), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n749), .A2(G125), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n812), .B2(new_n274), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n911), .A2(new_n1012), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n317), .B1(new_n1105), .B2(KEYINPUT53), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n760), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(KEYINPUT53), .B2(new_n1105), .C1(new_n1107), .C2(new_n765), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n738), .A2(G128), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n762), .B2(new_n924), .ZN(new_n1110));
  NOR3_X1   g0910(.A1(new_n1104), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G132), .A2(new_n757), .B1(new_n755), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1100), .A2(new_n1102), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n710), .B1(new_n991), .B2(new_n1095), .C1(new_n1115), .C2(new_n824), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1094), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n709), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1092), .A2(new_n1119), .ZN(G378));
  AOI21_X1  g0920(.A(new_n794), .B1(new_n900), .B2(new_n901), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n899), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n299), .A2(new_n302), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n838), .A2(new_n277), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1125), .B(new_n1126), .Z(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n899), .A2(new_n1121), .A3(new_n1127), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n893), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n891), .B1(new_n1093), .B2(new_n836), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n899), .A2(new_n1121), .A3(new_n1127), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1127), .B1(new_n899), .B2(new_n1121), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT120), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1131), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n893), .A2(new_n1129), .A3(KEYINPUT120), .A4(new_n1130), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n709), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1127), .A2(new_n723), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n710), .B1(G50), .B2(new_n1095), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n754), .A2(new_n305), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(G58), .A2(new_n748), .B1(new_n749), .B2(G283), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n317), .A2(new_n281), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n911), .B2(G77), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G97), .A2(new_n742), .B1(new_n738), .B2(G116), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n926), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1142), .B(new_n1147), .C1(G107), .C2(new_n757), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n760), .A2(G150), .B1(G125), .B2(new_n738), .ZN(new_n1150));
  INV_X1    g0950(.A(G132), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n762), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G137), .B2(new_n755), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n757), .A2(G128), .B1(new_n911), .B2(new_n1113), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1153), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n749), .A2(G124), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G33), .B(G41), .C1(new_n748), .C2(G159), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1148), .A2(KEYINPUT58), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1144), .B(new_n274), .C1(G33), .C2(G41), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1149), .A2(new_n1163), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1141), .B1(new_n1166), .B2(new_n726), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1140), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1139), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1083), .A2(new_n613), .A3(new_n1084), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT121), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT121), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n894), .A2(new_n1174), .A3(new_n1084), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1118), .B2(new_n1085), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1170), .B1(new_n1171), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1087), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1170), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n700), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1169), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(G375));
  AOI22_X1  g0983(.A1(new_n749), .A2(G128), .B1(G159), .B2(new_n911), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT122), .Z(new_n1185));
  OAI22_X1  g0985(.A1(new_n264), .A2(new_n754), .B1(new_n756), .B2(new_n924), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n317), .B1(new_n738), .B2(G132), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n762), .B2(new_n1112), .C1(new_n1107), .C2(new_n274), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(G58), .C2(new_n748), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n290), .B1(new_n911), .B2(G97), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G116), .A2(new_n742), .B1(new_n738), .B2(G294), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1014), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1192), .B(new_n923), .C1(G303), .C2(new_n749), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G107), .A2(new_n755), .B1(new_n757), .B2(G283), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1185), .A2(new_n1189), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n710), .B1(G68), .B2(new_n1095), .C1(new_n1195), .C2(new_n824), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT123), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n724), .B2(new_n886), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1072), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n1032), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1085), .A2(new_n981), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1172), .A2(new_n1199), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(G381));
  INV_X1    g1004(.A(G384), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n940), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n980), .A2(new_n982), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1032), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n960), .B(new_n961), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1206), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(G393), .A2(G396), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n1205), .A2(new_n1210), .A3(new_n1211), .A4(new_n1203), .ZN(new_n1212));
  AND3_X1   g1012(.A1(new_n1028), .A2(new_n1030), .A3(new_n1056), .ZN(new_n1213));
  INV_X1    g1013(.A(G378), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1212), .A2(new_n1182), .A3(new_n1213), .A4(new_n1214), .ZN(G407));
  NAND2_X1  g1015(.A1(new_n639), .A2(G213), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1182), .A2(new_n1214), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G407), .B(G213), .C1(new_n1216), .C2(new_n1217), .ZN(G409));
  INV_X1    g1018(.A(KEYINPUT63), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1169), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(G378), .A3(new_n1221), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1179), .A2(new_n982), .A3(new_n1138), .A4(new_n1137), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1032), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1140), .B2(new_n1167), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G378), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1216), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1200), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1202), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(KEYINPUT60), .B2(new_n1088), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1172), .A2(KEYINPUT60), .A3(new_n1199), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n699), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1230), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1205), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G384), .B(new_n1230), .C1(new_n1232), .C2(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1219), .B1(new_n1229), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1216), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G2897), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1238), .B(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT61), .B1(new_n1229), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n779), .B1(new_n988), .B2(new_n1022), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1211), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1210), .A2(G390), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1213), .A2(G387), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT124), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1210), .A2(new_n1250), .A3(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1248), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n1210), .B2(G390), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1245), .B(KEYINPUT125), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT124), .B1(new_n1213), .B2(G387), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1251), .A3(new_n1248), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT125), .B1(new_n1257), .B2(new_n1245), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1249), .B1(new_n1255), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1240), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1238), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(KEYINPUT63), .A3(new_n1261), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1239), .A2(new_n1243), .A3(new_n1259), .A4(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1241), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1238), .B(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1266), .B2(new_n1260), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT126), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1269), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1226), .B1(new_n1182), .B2(G378), .ZN(new_n1271));
  XOR2_X1   g1071(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1272));
  NOR4_X1   g1072(.A1(new_n1271), .A2(new_n1240), .A3(new_n1238), .A4(new_n1272), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1267), .A2(new_n1270), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1263), .B1(new_n1274), .B2(new_n1259), .ZN(G405));
  INV_X1    g1075(.A(new_n1249), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1257), .A2(new_n1245), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT125), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1276), .B1(new_n1279), .B2(new_n1254), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT127), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G375), .A2(G378), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1217), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1261), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1217), .A3(new_n1238), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1280), .A2(new_n1281), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1281), .B(new_n1249), .C1(new_n1255), .C2(new_n1258), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1286), .B1(new_n1289), .B2(new_n1290), .ZN(G402));
endmodule


