//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT72), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT73), .B1(new_n190), .B2(G104), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(new_n190), .A3(G104), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT74), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n197), .A2(new_n199), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(new_n203), .A3(new_n196), .A4(new_n195), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n196), .B1(new_n202), .B2(new_n195), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT4), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT0), .B(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n218), .B1(new_n206), .B2(new_n207), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n209), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT10), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  AND4_X1   g036(.A1(new_n222), .A2(new_n211), .A3(new_n213), .A4(G128), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT1), .B1(new_n212), .B2(G146), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n224), .A2(G128), .B1(new_n211), .B2(new_n213), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT75), .B1(new_n193), .B2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n193), .A2(G107), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n193), .A2(KEYINPUT75), .A3(G107), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n196), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AND4_X1   g046(.A1(new_n221), .A2(new_n205), .A3(new_n226), .A4(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n231), .B1(new_n201), .B2(new_n204), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n221), .B1(new_n234), .B2(new_n226), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n220), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT11), .ZN(new_n237));
  INV_X1    g051(.A(G134), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G137), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .A3(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G131), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n239), .A2(new_n241), .A3(new_n245), .A4(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n249), .B(new_n220), .C1(new_n233), .C2(new_n235), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G140), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n253), .A2(G227), .ZN(new_n254));
  XOR2_X1   g068(.A(new_n252), .B(new_n254), .Z(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n205), .A2(new_n226), .A3(new_n232), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT10), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n234), .A2(new_n221), .A3(new_n226), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n258), .A2(new_n259), .B1(new_n209), .B2(new_n219), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n256), .B1(new_n260), .B2(new_n249), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n223), .A2(new_n225), .ZN(new_n262));
  AOI211_X1 g076(.A(new_n231), .B(new_n262), .C1(new_n201), .C2(new_n204), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n226), .B1(new_n205), .B2(new_n232), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n247), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT12), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(KEYINPUT12), .B(new_n247), .C1(new_n263), .C2(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n251), .A2(new_n256), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n270), .A2(G469), .A3(G902), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n248), .A2(new_n250), .A3(new_n255), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n267), .A2(new_n268), .B1(new_n260), .B2(new_n249), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n272), .B(G469), .C1(new_n273), .C2(new_n255), .ZN(new_n274));
  NAND2_X1  g088(.A1(G469), .A2(G902), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n189), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(G475), .A2(G902), .ZN(new_n278));
  OR2_X1    g092(.A1(KEYINPUT68), .A2(G125), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT68), .A2(G125), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(G140), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(G125), .A2(G140), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n281), .A2(G146), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(G125), .B(G140), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n210), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(G237), .A2(G953), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(G143), .A3(G214), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G143), .B1(new_n288), .B2(G214), .ZN(new_n291));
  OAI211_X1 g105(.A(KEYINPUT18), .B(G131), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G237), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n253), .A3(G214), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n212), .ZN(new_n295));
  NAND2_X1  g109(.A1(KEYINPUT18), .A2(G131), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n289), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n287), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT80), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT80), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n287), .A2(new_n292), .A3(new_n300), .A4(new_n297), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n295), .A2(new_n245), .A3(new_n289), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT81), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT17), .ZN(new_n306));
  OAI21_X1  g120(.A(G131), .B1(new_n290), .B2(new_n291), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n295), .A2(KEYINPUT81), .A3(new_n245), .A4(new_n289), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(KEYINPUT16), .A2(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n279), .A2(new_n280), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(KEYINPUT68), .A2(G125), .ZN(new_n314));
  NOR2_X1   g128(.A1(KEYINPUT68), .A2(G125), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT69), .A3(new_n310), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n281), .B2(new_n283), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n210), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n307), .A2(new_n306), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n314), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT16), .B1(new_n324), .B2(new_n282), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n325), .A2(G146), .A3(new_n313), .A4(new_n317), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n309), .A2(new_n321), .A3(new_n322), .A4(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G113), .B(G122), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(new_n193), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n302), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n281), .A2(KEYINPUT19), .A3(new_n283), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT19), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n285), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n331), .B(new_n326), .C1(G146), .C2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n329), .B1(new_n302), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n330), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g153(.A(KEYINPUT82), .B(new_n329), .C1(new_n302), .C2(new_n336), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n278), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT20), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n343), .B(new_n278), .C1(new_n339), .C2(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(G475), .ZN(new_n345));
  INV_X1    g159(.A(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n330), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n329), .B1(new_n302), .B2(new_n327), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT83), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT83), .B(new_n346), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n342), .A2(new_n344), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n212), .B2(G128), .ZN(new_n355));
  INV_X1    g169(.A(G128), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT84), .A3(G143), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n355), .A2(new_n357), .B1(G128), .B2(new_n212), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G134), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G122), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(G116), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(G116), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n190), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n358), .B2(G134), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n361), .A2(G116), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT14), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n363), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(KEYINPUT85), .B(new_n363), .C1(new_n367), .C2(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n368), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G107), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n212), .A2(G128), .ZN(new_n377));
  INV_X1    g191(.A(new_n357), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT84), .B1(new_n356), .B2(G143), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT13), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n378), .B2(new_n379), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n382), .A3(G134), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n362), .A2(new_n363), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n364), .ZN(new_n386));
  OAI221_X1 g200(.A(new_n377), .B1(new_n381), .B2(new_n238), .C1(new_n378), .C2(new_n379), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n187), .A2(new_n390), .A3(G953), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n369), .A2(new_n370), .B1(new_n368), .B2(new_n367), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n190), .B1(new_n394), .B2(new_n372), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n380), .A2(new_n238), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n359), .A3(new_n364), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n388), .B(new_n391), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n346), .ZN(new_n400));
  INV_X1    g214(.A(G478), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT86), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n402), .A2(KEYINPUT15), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(KEYINPUT15), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n400), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n353), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n277), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n262), .B1(new_n315), .B2(new_n314), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n218), .A2(new_n316), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n253), .A2(G224), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT78), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(G110), .B(G122), .Z(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT5), .ZN(new_n420));
  INV_X1    g234(.A(G119), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n421), .A3(G116), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT76), .ZN(new_n423));
  INV_X1    g237(.A(G113), .ZN(new_n424));
  XNOR2_X1  g238(.A(G116), .B(G119), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(KEYINPUT5), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT2), .B(G113), .Z(new_n427));
  AOI22_X1  g241(.A1(new_n423), .A2(new_n426), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n205), .A2(new_n232), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n191), .A2(new_n194), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n197), .A2(new_n199), .ZN(new_n431));
  OAI21_X1  g245(.A(G101), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT4), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n204), .B2(new_n201), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n207), .B(G101), .C1(new_n430), .C2(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n427), .A2(new_n425), .ZN(new_n436));
  XOR2_X1   g250(.A(G116), .B(G119), .Z(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT2), .B(G113), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n429), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n419), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(KEYINPUT77), .B(new_n429), .C1(new_n434), .C2(new_n441), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n419), .B(new_n429), .C1(new_n434), .C2(new_n441), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n444), .A2(new_n445), .B1(KEYINPUT6), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n205), .A2(new_n232), .A3(new_n428), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n441), .B1(new_n205), .B2(new_n208), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n450), .A2(new_n445), .A3(KEYINPUT6), .A4(new_n418), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n417), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G210), .B1(G237), .B2(G902), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n415), .A2(KEYINPUT7), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n413), .A2(new_n455), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n413), .A2(new_n455), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n446), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n418), .B(KEYINPUT8), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n234), .A2(new_n428), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n460), .B2(new_n429), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n346), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n454), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n454), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n450), .A2(new_n418), .A3(new_n445), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n446), .A2(KEYINPUT6), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n416), .B1(new_n468), .B2(new_n451), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n465), .B1(new_n469), .B2(new_n462), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(new_n470), .A3(KEYINPUT79), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT79), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n472), .B(new_n465), .C1(new_n469), .C2(new_n462), .ZN(new_n473));
  NAND2_X1  g287(.A1(G234), .A2(G237), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(G952), .A3(new_n253), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n475), .B(KEYINPUT87), .Z(new_n476));
  XOR2_X1   g290(.A(KEYINPUT21), .B(G898), .Z(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(G902), .A3(G953), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n479), .B(KEYINPUT88), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n471), .A2(new_n473), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n242), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n238), .A2(G137), .ZN(new_n485));
  OAI21_X1  g299(.A(G131), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n486), .A2(new_n246), .ZN(new_n487));
  INV_X1    g301(.A(new_n218), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n226), .A2(new_n487), .B1(new_n247), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT30), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n247), .A2(new_n488), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n246), .B(new_n486), .C1(new_n223), .C2(new_n225), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n490), .A2(new_n495), .A3(new_n440), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n288), .A2(G210), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(G101), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n440), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n491), .A2(new_n502), .A3(new_n492), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT64), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n491), .A2(KEYINPUT64), .A3(new_n502), .A4(new_n492), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT65), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n496), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI211_X1 g323(.A(KEYINPUT65), .B(new_n501), .C1(new_n505), .C2(new_n506), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n511));
  OAI22_X1  g325(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(KEYINPUT31), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n511), .A2(KEYINPUT31), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n503), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n502), .B1(new_n491), .B2(new_n492), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n505), .B2(new_n506), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n517), .B2(new_n514), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n513), .B1(new_n518), .B2(new_n501), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT64), .B1(new_n489), .B2(new_n502), .ZN(new_n520));
  INV_X1    g334(.A(new_n506), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n500), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT65), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n507), .A2(new_n508), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n511), .A2(KEYINPUT31), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .A4(new_n496), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n512), .A2(new_n519), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G472), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n346), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT32), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n527), .A2(KEYINPUT32), .A3(new_n528), .A4(new_n346), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n496), .B1(new_n520), .B2(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n501), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n500), .B(new_n515), .C1(new_n517), .C2(new_n514), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n346), .B1(new_n536), .B2(new_n535), .ZN(new_n538));
  OAI21_X1  g352(.A(G472), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n531), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n390), .B1(G234), .B2(new_n346), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n253), .A2(G221), .A3(G234), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT71), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n326), .A2(new_n286), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n421), .A2(G128), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n356), .A2(G119), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT23), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n551), .A2(new_n356), .A3(G119), .ZN(new_n552));
  AOI211_X1 g366(.A(KEYINPUT70), .B(G110), .C1(new_n550), .C2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT23), .B1(new_n421), .B2(G128), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n356), .A2(G119), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G110), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  OAI21_X1  g374(.A(KEYINPUT67), .B1(new_n356), .B2(G119), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT67), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(new_n421), .A3(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n549), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n553), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n547), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n561), .A2(new_n563), .B1(G119), .B2(new_n356), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n560), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n558), .B2(new_n557), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n321), .B2(new_n326), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n546), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n570), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT69), .B1(new_n316), .B2(new_n310), .ZN(new_n574));
  AND4_X1   g388(.A1(KEYINPUT69), .A2(new_n279), .A3(new_n280), .A4(new_n310), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(G146), .B1(new_n576), .B2(new_n325), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n318), .A2(new_n210), .A3(new_n320), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(G110), .B1(new_n550), .B2(new_n552), .ZN(new_n580));
  OAI22_X1  g394(.A1(new_n580), .A2(new_n554), .B1(new_n568), .B2(new_n560), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n326), .B(new_n286), .C1(new_n581), .C2(new_n553), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n582), .A3(new_n545), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n572), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT25), .B1(new_n584), .B2(new_n346), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n586), .B(G902), .C1(new_n572), .C2(new_n583), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n541), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n541), .A2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n410), .A2(new_n483), .A3(new_n540), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  AOI21_X1  g407(.A(new_n454), .B1(new_n453), .B2(new_n463), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n469), .A2(new_n465), .A3(new_n462), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n482), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n351), .A2(new_n352), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n302), .A2(new_n336), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT82), .B1(new_n598), .B2(new_n329), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n337), .A2(new_n338), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n330), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n343), .B1(new_n601), .B2(new_n278), .ZN(new_n602));
  INV_X1    g416(.A(new_n344), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n399), .A2(KEYINPUT89), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n398), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n391), .B1(new_n376), .B2(new_n388), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT89), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n399), .A2(KEYINPUT90), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT90), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n605), .B1(new_n393), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n606), .A2(new_n611), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n401), .A2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n400), .A2(new_n401), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n604), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT91), .B1(new_n596), .B2(new_n620), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n615), .A2(new_n616), .B1(new_n401), .B2(new_n400), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n353), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT91), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n464), .A2(new_n470), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .A4(new_n482), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n527), .A2(new_n346), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n591), .A3(new_n529), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n277), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n342), .A2(new_n344), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n302), .A2(new_n327), .ZN(new_n636));
  INV_X1    g450(.A(new_n329), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n638), .B2(new_n330), .ZN(new_n639));
  OAI21_X1  g453(.A(G475), .B1(new_n639), .B2(KEYINPUT83), .ZN(new_n640));
  INV_X1    g454(.A(new_n352), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT92), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT92), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n351), .A2(new_n643), .A3(new_n352), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n635), .A2(new_n642), .A3(new_n407), .A4(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n596), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n631), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n190), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  NOR2_X1   g464(.A1(new_n545), .A2(KEYINPUT36), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n567), .A2(new_n571), .A3(KEYINPUT94), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT94), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n579), .B2(new_n582), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n652), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT94), .B1(new_n567), .B2(new_n571), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n579), .A2(new_n654), .A3(new_n582), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n651), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(new_n589), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT95), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n656), .A2(KEYINPUT95), .A3(new_n589), .A4(new_n659), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n588), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n629), .A2(new_n529), .A3(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT96), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n629), .A2(KEYINPUT96), .A3(new_n529), .A4(new_n664), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n667), .A2(new_n483), .A3(new_n410), .A4(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT37), .B(G110), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT97), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n669), .B(new_n671), .ZN(G12));
  OAI211_X1 g486(.A(new_n481), .B(new_n664), .C1(new_n594), .C2(new_n595), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n476), .B1(G900), .B2(new_n478), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n645), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n189), .ZN(new_n678));
  INV_X1    g492(.A(new_n276), .ZN(new_n679));
  INV_X1    g493(.A(G469), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n250), .A2(new_n255), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n268), .B2(new_n267), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n255), .B1(new_n248), .B2(new_n250), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n680), .B(new_n346), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n678), .B1(new_n679), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n674), .A2(new_n540), .A3(new_n677), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  NAND2_X1  g501(.A1(new_n471), .A2(new_n473), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n509), .A2(new_n510), .ZN(new_n691));
  INV_X1    g505(.A(new_n517), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n501), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n531), .A2(new_n532), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n675), .B(KEYINPUT39), .Z(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n685), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT40), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n353), .A2(new_n408), .ZN(new_n702));
  INV_X1    g516(.A(new_n481), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n664), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n697), .B(new_n705), .C1(KEYINPUT40), .C2(new_n700), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G143), .ZN(G45));
  NOR3_X1   g521(.A1(new_n353), .A2(new_n622), .A3(new_n676), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n674), .A2(new_n540), .A3(new_n685), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND2_X1  g524(.A1(new_n540), .A2(new_n591), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n270), .B2(G902), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT99), .A3(new_n684), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT99), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n714), .B(G469), .C1(new_n270), .C2(G902), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n188), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT100), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n188), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n720), .B1(new_n713), .B2(new_n715), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n711), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT101), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n724), .A3(new_n627), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n540), .A2(new_n591), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT100), .B1(new_n716), .B2(new_n188), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n718), .B(new_n720), .C1(new_n713), .C2(new_n715), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n627), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT41), .B(G113), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT102), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n731), .B(new_n733), .ZN(G15));
  OAI211_X1 g548(.A(new_n726), .B(new_n646), .C1(new_n727), .C2(new_n728), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G116), .ZN(G18));
  AND4_X1   g550(.A1(new_n480), .A2(new_n353), .A3(new_n408), .A4(new_n664), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n703), .B1(new_n464), .B2(new_n470), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n721), .A2(new_n540), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  NAND3_X1  g555(.A1(new_n702), .A2(new_n738), .A3(new_n480), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n630), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n727), .B2(new_n728), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  AND3_X1   g559(.A1(new_n629), .A2(new_n529), .A3(new_n664), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n746), .A2(new_n721), .A3(new_n738), .A4(new_n708), .ZN(new_n747));
  XOR2_X1   g561(.A(KEYINPUT104), .B(G125), .Z(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G27));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n711), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n540), .A2(KEYINPUT106), .A3(new_n591), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n720), .B1(new_n679), .B2(new_n684), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT105), .B1(new_n688), .B2(new_n481), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n756), .B(new_n703), .C1(new_n471), .C2(new_n473), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n753), .A2(new_n708), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n688), .A2(new_n481), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n756), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n688), .A2(KEYINPUT105), .A3(new_n481), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n726), .A2(new_n761), .A3(new_n754), .A4(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n708), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(KEYINPUT42), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n759), .A2(KEYINPUT42), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G131), .ZN(G33));
  NAND4_X1  g581(.A1(new_n758), .A2(new_n726), .A3(new_n677), .A4(new_n754), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  OAI21_X1  g583(.A(new_n272), .B1(new_n273), .B2(new_n255), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n680), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n771), .B2(new_n770), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n275), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n271), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(KEYINPUT46), .B2(new_n774), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n188), .A3(new_n699), .ZN(new_n777));
  XNOR2_X1  g591(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT43), .B1(new_n353), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n619), .A2(new_n353), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n629), .A2(new_n529), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n664), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n761), .A2(new_n762), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n786), .B2(new_n787), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n779), .A2(new_n780), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  XOR2_X1   g605(.A(KEYINPUT110), .B(G137), .Z(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G39));
  NAND2_X1  g607(.A1(new_n776), .A2(new_n188), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n764), .A2(new_n540), .A3(new_n591), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n758), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G140), .ZN(G42));
  NOR2_X1   g613(.A1(new_n789), .A2(new_n717), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT116), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n476), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n784), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n753), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n629), .A2(new_n529), .A3(new_n591), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n189), .B1(new_n713), .B2(new_n715), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n758), .B(new_n810), .C1(new_n796), .C2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n803), .A2(new_n746), .A3(new_n805), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n690), .A2(new_n703), .A3(new_n721), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT50), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n812), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n696), .A2(new_n591), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n476), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n803), .A2(KEYINPUT117), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n801), .A2(new_n802), .A3(new_n819), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n820), .A2(new_n353), .A3(new_n622), .A4(new_n823), .ZN(new_n824));
  AND2_X1   g638(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n807), .B1(new_n825), .B2(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n253), .A2(G952), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n721), .A2(new_n738), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n810), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n821), .B(new_n822), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n620), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT118), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n817), .A2(KEYINPUT51), .A3(new_n824), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n834), .B(new_n829), .C1(new_n830), .C2(new_n620), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n826), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT103), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n739), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n735), .A2(new_n744), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n766), .A2(new_n838), .A3(new_n731), .A4(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT114), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n625), .A2(new_n481), .A3(new_n604), .A4(new_n407), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n684), .A2(new_n275), .A3(new_n274), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n588), .A2(new_n662), .A3(new_n663), .A4(new_n675), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n847), .A2(new_n848), .A3(new_n188), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n849), .A3(new_n695), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n747), .A2(new_n686), .A3(new_n709), .A4(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT52), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT112), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n635), .A2(new_n642), .A3(new_n644), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n407), .A2(new_n676), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n758), .B2(new_n857), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n755), .A2(new_n757), .A3(KEYINPUT112), .A4(new_n856), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n540), .A2(new_n685), .A3(new_n664), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n353), .A2(new_n407), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n483), .A2(new_n808), .A3(new_n685), .A4(new_n863), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n669), .A2(new_n592), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n483), .A2(KEYINPUT111), .A3(new_n623), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n623), .A2(new_n471), .A3(new_n473), .A4(new_n482), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n869), .A3(new_n631), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n764), .A2(new_n665), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n758), .A2(new_n871), .A3(new_n754), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n865), .A2(new_n768), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n852), .A2(new_n861), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n735), .A2(new_n744), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n724), .B1(new_n723), .B2(new_n627), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n729), .A2(KEYINPUT101), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n740), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n758), .A2(new_n708), .A3(new_n754), .ZN(new_n879));
  INV_X1    g693(.A(new_n752), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT106), .B1(new_n540), .B2(new_n591), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT42), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n763), .A2(new_n765), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT113), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n844), .A2(new_n845), .A3(new_n874), .A4(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(KEYINPUT53), .A3(new_n874), .A4(new_n843), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT114), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n878), .A2(new_n885), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT53), .B1(new_n890), .B2(new_n874), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n887), .A2(new_n889), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n890), .A2(new_n874), .A3(KEYINPUT53), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OAI22_X1  g713(.A1(new_n837), .A2(new_n899), .B1(G952), .B2(G953), .ZN(new_n900));
  INV_X1    g714(.A(new_n818), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT49), .B1(new_n713), .B2(new_n715), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n902), .A2(new_n703), .A3(new_n678), .A4(new_n783), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n713), .A2(KEYINPUT49), .A3(new_n715), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n901), .A2(new_n903), .A3(new_n690), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n900), .A2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n447), .A2(new_n452), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(new_n417), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT55), .Z(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n887), .A2(new_n889), .A3(new_n892), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(G210), .A3(G902), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n912), .A2(KEYINPUT119), .A3(new_n913), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n910), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n253), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT119), .B1(new_n912), .B2(new_n913), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n909), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n918), .A2(new_n922), .ZN(G51));
  NAND2_X1  g737(.A1(new_n911), .A2(new_n893), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n925), .A3(new_n895), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n911), .A2(KEYINPUT120), .A3(new_n893), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n275), .B(KEYINPUT57), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n270), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n911), .A2(G902), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n932), .A2(new_n773), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n919), .B1(new_n931), .B2(new_n933), .ZN(G54));
  INV_X1    g748(.A(new_n601), .ZN(new_n935));
  NAND2_X1  g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n920), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(G60));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT59), .Z(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n895), .B2(new_n898), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n920), .B1(new_n943), .B2(new_n615), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n926), .A2(new_n927), .ZN(new_n945));
  INV_X1    g759(.A(new_n615), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(new_n942), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n945), .B2(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT121), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n911), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n656), .A2(new_n659), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n920), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n953), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n956), .B(KEYINPUT61), .C1(new_n584), .C2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n584), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n955), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n958), .A2(new_n961), .ZN(G66));
  AOI21_X1  g776(.A(new_n253), .B1(new_n477), .B2(G224), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n842), .A2(new_n731), .A3(new_n870), .A4(new_n865), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT122), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n963), .B1(new_n965), .B2(new_n253), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n907), .B1(G898), .B2(new_n253), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT123), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n966), .B(new_n968), .ZN(G69));
  NAND2_X1  g783(.A1(new_n490), .A2(new_n495), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(new_n335), .Z(new_n971));
  NAND3_X1  g785(.A1(new_n747), .A2(new_n686), .A3(new_n709), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n706), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n620), .A2(new_n862), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(KEYINPUT124), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n685), .B(new_n699), .C1(new_n978), .C2(KEYINPUT124), .ZN(new_n980));
  OR4_X1    g794(.A1(new_n711), .A2(new_n789), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n798), .A2(new_n791), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n971), .B1(new_n983), .B2(G953), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n798), .A2(new_n791), .A3(new_n766), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n779), .A2(new_n780), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n753), .A2(new_n846), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n768), .B(new_n973), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n253), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n253), .A2(G900), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT125), .Z(new_n991));
  AND2_X1   g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n984), .B1(new_n992), .B2(new_n971), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT63), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT126), .ZN(new_n998));
  INV_X1    g812(.A(new_n983), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n965), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n500), .A3(new_n533), .ZN(new_n1001));
  INV_X1    g815(.A(new_n691), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n997), .B1(new_n1002), .B2(new_n534), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n897), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1001), .A2(new_n920), .A3(new_n1004), .ZN(new_n1005));
  OR3_X1    g819(.A1(new_n965), .A2(new_n985), .A3(new_n988), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n1006), .A2(new_n998), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n500), .B(new_n533), .C1(new_n1007), .C2(KEYINPUT127), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1007), .A2(KEYINPUT127), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1005), .B1(new_n1008), .B2(new_n1009), .ZN(G57));
endmodule


