//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034;
  XNOR2_X1  g000(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G183gat), .B(G211gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  OR2_X1    g007(.A1(G71gat), .A2(G78gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT9), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n208), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT100), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n209), .A2(new_n208), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT100), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n214), .B(new_n215), .C1(new_n211), .C2(new_n210), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT101), .ZN(new_n217));
  INV_X1    g016(.A(G64gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G57gat), .ZN(new_n219));
  INV_X1    g018(.A(G57gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(KEYINPUT101), .A3(G64gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n219), .B(new_n221), .C1(new_n220), .C2(G64gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n208), .B1(new_n209), .B2(new_n211), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n213), .A2(new_n216), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n227), .B1(G231gat), .B2(G233gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G231gat), .A2(G233gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n229), .B1(new_n225), .B2(new_n226), .ZN(new_n230));
  OAI21_X1  g029(.A(G127gat), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n228), .A2(G127gat), .A3(new_n230), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n234), .A2(G1gat), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n236), .A2(KEYINPUT94), .A3(KEYINPUT16), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT94), .B1(new_n236), .B2(KEYINPUT16), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT95), .B(G8gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT96), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G8gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT96), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n235), .A2(new_n239), .A3(new_n245), .A4(new_n240), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n225), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(KEYINPUT21), .B2(new_n248), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n232), .A2(new_n233), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  OR3_X1    g050(.A1(new_n228), .A2(G127gat), .A3(new_n230), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n251), .B1(new_n252), .B2(new_n231), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n207), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n249), .B1(new_n232), .B2(new_n233), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n231), .A3(new_n251), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n206), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(G232gat), .A2(G233gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(KEYINPUT41), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(KEYINPUT41), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT90), .B(G36gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G29gat), .ZN(new_n264));
  OR3_X1    g063(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(G43gat), .A2(G50gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(G43gat), .A2(G50gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT15), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(new_n267), .A3(new_n271), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT92), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT91), .B(G50gat), .ZN(new_n275));
  INV_X1    g074(.A(G43gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n269), .A2(KEYINPUT15), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n273), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(KEYINPUT92), .A3(new_n278), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n272), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G85gat), .A2(G92gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT7), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(G99gat), .A2(G106gat), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n287), .A2(KEYINPUT8), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT102), .ZN(new_n289));
  NOR2_X1   g088(.A1(G85gat), .A2(G92gat), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G85gat), .ZN(new_n292));
  INV_X1    g091(.A(G92gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(KEYINPUT8), .A2(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(KEYINPUT102), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n286), .B1(new_n291), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G99gat), .B(G106gat), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(KEYINPUT102), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n297), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n302), .A3(new_n286), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n262), .B1(new_n282), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT103), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n279), .A2(new_n274), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n307), .A2(new_n271), .A3(new_n268), .A4(new_n281), .ZN(new_n308));
  OR2_X1    g107(.A1(new_n268), .A2(new_n271), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT17), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT93), .B(KEYINPUT17), .Z(new_n311));
  OAI211_X1 g110(.A(new_n310), .B(new_n304), .C1(new_n282), .C2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n261), .B1(new_n306), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n305), .A2(KEYINPUT103), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n305), .A2(KEYINPUT103), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n312), .B(new_n261), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G190gat), .B(G218gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(KEYINPUT104), .ZN(new_n319));
  XOR2_X1   g118(.A(G134gat), .B(G162gat), .Z(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n321), .ZN(new_n323));
  INV_X1    g122(.A(new_n317), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n323), .B1(new_n324), .B2(new_n313), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n258), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT105), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT105), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n258), .A2(new_n322), .A3(new_n325), .A4(new_n328), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n212), .A2(KEYINPUT100), .B1(new_n223), .B2(new_n222), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n298), .A2(new_n216), .A3(new_n330), .A4(new_n303), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n302), .B1(new_n301), .B2(new_n286), .ZN(new_n332));
  AOI211_X1 g131(.A(new_n297), .B(new_n285), .C1(new_n299), .C2(new_n300), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n225), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT106), .B(KEYINPUT10), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n331), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n332), .A2(new_n333), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n248), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n331), .A2(new_n334), .ZN(new_n342));
  INV_X1    g141(.A(new_n340), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G120gat), .B(G148gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G176gat), .B(G204gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT107), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT107), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n341), .A2(new_n350), .A3(new_n344), .A4(new_n347), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n343), .B1(new_n336), .B2(new_n338), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n343), .B2(new_n342), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n354), .A2(new_n347), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n327), .A2(new_n329), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n359), .B(new_n310), .C1(new_n282), .C2(new_n311), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n308), .A2(new_n309), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n361), .A2(new_n247), .B1(G229gat), .B2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT18), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n362), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT97), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n359), .A2(new_n282), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n247), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G229gat), .A2(G233gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n371), .B(KEYINPUT13), .Z(new_n372));
  AOI21_X1  g171(.A(new_n367), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  AOI211_X1 g173(.A(KEYINPUT97), .B(new_n374), .C1(new_n368), .C2(new_n369), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n365), .B(new_n366), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(G113gat), .B(G141gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G197gat), .ZN(new_n378));
  XOR2_X1   g177(.A(KEYINPUT11), .B(G169gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT12), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n369), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n361), .A2(new_n247), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n372), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT97), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n367), .A3(new_n372), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n362), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT18), .B1(new_n360), .B2(new_n362), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n392), .A3(new_n381), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n383), .A2(KEYINPUT98), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT98), .B1(new_n383), .B2(new_n393), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XOR2_X1   g195(.A(G155gat), .B(G162gat), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G141gat), .B(G148gat), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT77), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT2), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G141gat), .ZN(new_n402));
  INV_X1    g201(.A(G148gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(KEYINPUT77), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n398), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408));
  INV_X1    g207(.A(G162gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n203), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n413));
  AND2_X1   g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(G141gat), .A2(G148gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n404), .A2(KEYINPUT78), .A3(new_n405), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(new_n407), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT79), .ZN(new_n421));
  XOR2_X1   g220(.A(G127gat), .B(G134gat), .Z(new_n422));
  XNOR2_X1  g221(.A(G113gat), .B(G120gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(KEYINPUT1), .B2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G113gat), .B(G120gat), .Z(new_n425));
  INV_X1    g224(.A(KEYINPUT1), .ZN(new_n426));
  XNOR2_X1  g225(.A(G127gat), .B(G134gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n428), .A3(KEYINPUT80), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n428), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT80), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n420), .A2(new_n421), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n400), .B1(new_n414), .B2(new_n415), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n406), .A3(new_n408), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n397), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n418), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n436), .A2(new_n440), .A3(new_n418), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n418), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n433), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n436), .A2(new_n418), .A3(new_n428), .A4(new_n424), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT4), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n399), .A2(new_n413), .B1(new_n410), .B2(new_n411), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n435), .A2(new_n397), .B1(new_n449), .B2(new_n417), .ZN(new_n450));
  INV_X1    g249(.A(new_n430), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT5), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n445), .A2(new_n446), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT5), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n432), .A2(new_n429), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n443), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n447), .ZN(new_n459));
  INV_X1    g258(.A(new_n446), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n440), .B1(new_n450), .B2(new_n437), .ZN(new_n463));
  INV_X1    g262(.A(new_n441), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n421), .B1(new_n450), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n444), .A3(new_n457), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n446), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT83), .B1(new_n448), .B2(new_n453), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n447), .B2(KEYINPUT4), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n461), .B(new_n462), .C1(new_n469), .C2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n445), .B(new_n446), .C1(new_n472), .C2(new_n470), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n462), .B1(new_n476), .B2(new_n461), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n455), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G1gat), .B(G29gat), .Z(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT0), .ZN(new_n480));
  XNOR2_X1  g279(.A(G57gat), .B(G85gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n478), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n482), .B(new_n455), .C1(new_n475), .C2(new_n477), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n455), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n461), .B1(new_n469), .B2(new_n473), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT84), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n490), .B2(new_n474), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n482), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n484), .B1(new_n487), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(G8gat), .B(G36gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(G64gat), .B(G92gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n494), .B(new_n495), .Z(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT74), .B(G197gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G204gat), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n500), .A2(G204gat), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G211gat), .B(G218gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT75), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n504), .B(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(G226gat), .A2(G233gat), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(KEYINPUT29), .ZN(new_n510));
  AND2_X1   g309(.A1(KEYINPUT69), .A2(G190gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(KEYINPUT69), .A2(G190gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G183gat), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT28), .ZN(new_n515));
  AND2_X1   g314(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(KEYINPUT68), .A2(G183gat), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT27), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g317(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT28), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G183gat), .A2(G190gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(G169gat), .A2(G176gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(G169gat), .A2(G176gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT26), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n524), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT71), .B(new_n524), .C1(new_n528), .C2(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n523), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT68), .B(G183gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT69), .B(G190gat), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n516), .A2(new_n517), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n513), .A3(KEYINPUT70), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT24), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(new_n526), .B2(KEYINPUT23), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT23), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n549), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT25), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n526), .B2(KEYINPUT23), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n551), .A2(new_n525), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT65), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n544), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n557));
  OR2_X1    g356(.A1(G183gat), .A2(G190gat), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n556), .A2(new_n543), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G169gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT66), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT66), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G169gat), .ZN(new_n563));
  INV_X1    g362(.A(G176gat), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT23), .A4(new_n564), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n559), .A2(new_n551), .A3(new_n525), .A4(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n567));
  AOI22_X1  g366(.A1(new_n546), .A2(new_n554), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n535), .A2(new_n568), .A3(KEYINPUT76), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT76), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n546), .A2(new_n554), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n567), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT28), .B1(new_n520), .B2(new_n513), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n532), .B(new_n533), .C1(new_n574), .C2(new_n515), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n510), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n535), .A2(new_n568), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n509), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n508), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT76), .B1(new_n535), .B2(new_n568), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n570), .A3(new_n575), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n509), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n510), .B1(new_n535), .B2(new_n568), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n583), .A2(new_n584), .A3(new_n508), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n497), .B1(new_n580), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n584), .A3(new_n508), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n581), .A2(new_n582), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n588), .A2(new_n510), .B1(new_n509), .B2(new_n578), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n587), .B(new_n496), .C1(new_n589), .C2(new_n508), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(KEYINPUT30), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n580), .A2(new_n585), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n593), .A3(new_n496), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n493), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G78gat), .B(G106gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(KEYINPUT31), .B(G50gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n442), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n508), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT74), .B(G197gat), .Z(new_n605));
  INV_X1    g404(.A(G204gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n498), .B1(new_n607), .B2(new_n501), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n601), .B1(new_n608), .B2(new_n506), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n506), .B(new_n499), .C1(new_n502), .C2(new_n503), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT85), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n504), .A2(new_n505), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT85), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n613), .A2(new_n614), .A3(new_n601), .A4(new_n610), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n437), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n443), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT29), .B1(new_n439), .B2(new_n441), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n608), .B(new_n507), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT86), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G228gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n466), .B1(new_n508), .B2(KEYINPUT29), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n624), .B2(new_n443), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n508), .B1(new_n618), .B2(KEYINPUT87), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n618), .A2(KEYINPUT87), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G22gat), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n623), .B2(new_n628), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n600), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n623), .A2(new_n628), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(G22gat), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n599), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G15gat), .B(G43gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT73), .ZN(new_n639));
  XNOR2_X1  g438(.A(G71gat), .B(G99gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(G227gat), .ZN(new_n642));
  INV_X1    g441(.A(G233gat), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n535), .A2(new_n568), .A3(new_n430), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n451), .B1(new_n573), .B2(new_n575), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n641), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT72), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n647), .A2(new_n650), .A3(KEYINPUT32), .ZN(new_n651));
  INV_X1    g450(.A(new_n644), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n430), .B1(new_n535), .B2(new_n568), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n573), .A2(new_n451), .A3(new_n575), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT32), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT72), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n649), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n647), .B(KEYINPUT32), .C1(new_n648), .C2(new_n641), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(new_n652), .A3(new_n654), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT34), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n658), .A2(new_n662), .A3(new_n659), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n637), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT35), .B1(new_n596), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n666), .B1(new_n636), .B2(new_n632), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n482), .B(KEYINPUT88), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n485), .B(new_n486), .C1(new_n491), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n484), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT35), .B1(new_n591), .B2(new_n594), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n670), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n587), .B1(new_n589), .B2(new_n508), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(KEYINPUT37), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n497), .B1(new_n678), .B2(KEYINPUT37), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT38), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n590), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n497), .A2(KEYINPUT37), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n586), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n583), .A2(new_n584), .A3(new_n619), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n685), .A2(KEYINPUT37), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n577), .A2(new_n579), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n508), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT38), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n682), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n673), .A2(new_n484), .A3(new_n681), .A4(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT89), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n448), .A2(new_n453), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n465), .B2(new_n468), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT39), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n460), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n672), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n446), .B1(new_n445), .B2(new_n693), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n458), .A2(new_n446), .A3(new_n447), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT39), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n697), .A2(new_n701), .A3(KEYINPUT40), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT40), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n671), .B1(new_n698), .B2(new_n695), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n694), .A2(new_n460), .ZN(new_n705));
  INV_X1    g504(.A(new_n700), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  OAI22_X1  g507(.A1(new_n491), .A2(new_n672), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n692), .B1(new_n709), .B2(new_n595), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n591), .A2(new_n594), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT40), .B1(new_n697), .B2(new_n701), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n704), .A2(new_n703), .A3(new_n707), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n478), .A2(new_n671), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n711), .A2(new_n714), .A3(KEYINPUT89), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n691), .A2(new_n710), .A3(new_n715), .A4(new_n637), .ZN(new_n716));
  INV_X1    g515(.A(new_n637), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n596), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT36), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n666), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n664), .A2(KEYINPUT36), .A3(new_n665), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n716), .A2(new_n718), .A3(new_n722), .ZN(new_n723));
  AOI211_X1 g522(.A(KEYINPUT99), .B(new_n396), .C1(new_n677), .C2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT99), .ZN(new_n725));
  AND4_X1   g524(.A1(new_n691), .A2(new_n710), .A3(new_n715), .A4(new_n637), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n478), .A2(new_n483), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n727), .A2(new_n486), .A3(new_n485), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n711), .B1(new_n728), .B2(new_n484), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n722), .B1(new_n729), .B2(new_n637), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT35), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n729), .B2(new_n670), .ZN(new_n732));
  AND4_X1   g531(.A1(new_n674), .A2(new_n637), .A3(new_n667), .A4(new_n675), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n726), .A2(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n396), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n725), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n358), .B1(new_n724), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g538(.A(KEYINPUT108), .B(new_n358), .C1(new_n724), .C2(new_n736), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n493), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(G1gat), .ZN(G1324gat));
  INV_X1    g543(.A(G8gat), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n741), .B2(new_n711), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT16), .B(G8gat), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n595), .B(new_n747), .C1(new_n739), .C2(new_n740), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT42), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n741), .A2(new_n711), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n751), .B2(new_n747), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(G1325gat));
  INV_X1    g552(.A(G15gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n741), .A2(new_n754), .A3(new_n667), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n722), .B1(new_n739), .B2(new_n740), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(new_n754), .ZN(G1326gat));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n717), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT43), .B(G22gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1327gat));
  NOR2_X1   g559(.A1(new_n724), .A2(new_n736), .ZN(new_n761));
  INV_X1    g560(.A(new_n258), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n356), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n322), .A2(new_n325), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(G29gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n769), .A3(new_n742), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n774));
  INV_X1    g573(.A(new_n734), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n765), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n734), .A2(KEYINPUT44), .A3(new_n764), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n376), .A2(new_n382), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n381), .B1(new_n389), .B2(new_n392), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n763), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n778), .A2(new_n742), .A3(new_n782), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n772), .B(new_n773), .C1(new_n769), .C2(new_n783), .ZN(G1328gat));
  NOR2_X1   g583(.A1(new_n595), .A2(new_n263), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n766), .B(new_n785), .C1(new_n724), .C2(new_n736), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n776), .A2(new_n711), .A3(new_n777), .A4(new_n782), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n263), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n787), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(G1329gat));
  INV_X1    g592(.A(new_n722), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n778), .A2(G43gat), .A3(new_n794), .A4(new_n782), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n761), .A2(new_n666), .A3(new_n767), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(G43gat), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g597(.A(new_n275), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n778), .A2(new_n717), .A3(new_n799), .A4(new_n782), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n761), .A2(new_n637), .A3(new_n767), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g602(.A1(new_n352), .A2(new_n355), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n327), .A2(new_n781), .A3(new_n329), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n775), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n493), .B(KEYINPUT110), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g608(.A1(new_n775), .A2(new_n595), .A3(new_n805), .ZN(new_n810));
  NOR2_X1   g609(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n811));
  AND2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n810), .B2(new_n811), .ZN(G1333gat));
  NAND2_X1  g613(.A1(new_n806), .A2(new_n794), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n666), .A2(G71gat), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n815), .A2(G71gat), .B1(new_n806), .B2(new_n816), .ZN(new_n817));
  XOR2_X1   g616(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n818));
  XNOR2_X1  g617(.A(new_n817), .B(new_n818), .ZN(G1334gat));
  NAND2_X1  g618(.A1(new_n806), .A2(new_n717), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G78gat), .ZN(G1335gat));
  INV_X1    g620(.A(new_n781), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(new_n258), .A3(new_n356), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n776), .A2(new_n777), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT112), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n776), .A2(new_n826), .A3(new_n777), .A4(new_n823), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n825), .A2(new_n742), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n734), .A2(new_n781), .A3(new_n762), .A4(new_n764), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n829), .A2(new_n830), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n804), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n742), .A2(new_n292), .ZN(new_n835));
  OAI22_X1  g634(.A1(new_n828), .A2(new_n292), .B1(new_n834), .B2(new_n835), .ZN(G1336gat));
  NOR3_X1   g635(.A1(new_n356), .A2(new_n595), .A3(G92gat), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT113), .ZN(new_n838));
  INV_X1    g637(.A(new_n833), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n831), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  OAI21_X1  g640(.A(G92gat), .B1(new_n824), .B2(new_n595), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n825), .A2(new_n711), .A3(new_n827), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n840), .B1(new_n844), .B2(G92gat), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(G1337gat));
  NAND3_X1  g646(.A1(new_n825), .A2(new_n794), .A3(new_n827), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G99gat), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n666), .A2(G99gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n834), .B2(new_n850), .ZN(G1338gat));
  XNOR2_X1  g650(.A(KEYINPUT114), .B(G106gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(new_n824), .B2(new_n637), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n637), .A2(G106gat), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n853), .B(new_n854), .C1(new_n834), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n834), .A2(new_n856), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n825), .A2(new_n717), .A3(new_n827), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n852), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n857), .B1(new_n860), .B2(new_n854), .ZN(G1339gat));
  NOR2_X1   g660(.A1(new_n357), .A2(new_n822), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n336), .A2(new_n338), .A3(new_n343), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n341), .A2(KEYINPUT54), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n347), .B1(new_n353), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n864), .A2(KEYINPUT55), .A3(new_n866), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n352), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n781), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n370), .A2(new_n372), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n371), .B1(new_n360), .B2(new_n369), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n380), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n393), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n356), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n765), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n352), .A2(new_n869), .A3(new_n870), .ZN(new_n879));
  INV_X1    g678(.A(new_n876), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n764), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n862), .B1(new_n762), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n668), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(new_n742), .A3(new_n595), .ZN(new_n885));
  INV_X1    g684(.A(G113gat), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n885), .A2(new_n886), .A3(new_n396), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n807), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n884), .A2(new_n890), .A3(new_n807), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n711), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n822), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n887), .B1(new_n893), .B2(new_n886), .ZN(G1340gat));
  INV_X1    g693(.A(G120gat), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n885), .A2(new_n895), .A3(new_n356), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n804), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n895), .ZN(G1341gat));
  INV_X1    g697(.A(G127gat), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n885), .A2(new_n899), .A3(new_n762), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT116), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n711), .B(new_n762), .C1(new_n889), .C2(new_n891), .ZN(new_n902));
  OR2_X1    g701(.A1(new_n902), .A2(KEYINPUT117), .ZN(new_n903));
  AOI21_X1  g702(.A(G127gat), .B1(new_n902), .B2(KEYINPUT117), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(G1342gat));
  INV_X1    g704(.A(new_n892), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n765), .A2(G134gat), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n906), .A2(KEYINPUT56), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G134gat), .B1(new_n885), .B2(new_n765), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT56), .B1(new_n906), .B2(new_n908), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G1343gat));
  NAND2_X1  g711(.A1(new_n742), .A2(new_n595), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n794), .ZN(new_n914));
  INV_X1    g713(.A(new_n862), .ZN(new_n915));
  INV_X1    g714(.A(new_n881), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n879), .B1(new_n394), .B2(new_n395), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n880), .A2(new_n804), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n764), .B1(new_n919), .B2(KEYINPUT118), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n917), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n915), .B1(new_n923), .B2(new_n258), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n637), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT119), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT98), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(new_n779), .B2(new_n780), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n383), .A2(new_n393), .A3(KEYINPUT98), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n871), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT118), .B1(new_n931), .B2(new_n877), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n922), .A3(new_n765), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n258), .B1(new_n933), .B2(new_n881), .ZN(new_n934));
  OAI211_X1 g733(.A(KEYINPUT119), .B(new_n926), .C1(new_n934), .C2(new_n862), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n925), .B1(new_n883), .B2(new_n637), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n914), .B1(new_n927), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G141gat), .B1(new_n938), .B2(new_n396), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n883), .A2(new_n637), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n807), .A2(new_n595), .A3(new_n722), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(G141gat), .A3(new_n396), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT58), .ZN(new_n947));
  OAI211_X1 g746(.A(KEYINPUT58), .B(G141gat), .C1(new_n938), .C2(new_n781), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n943), .B1(new_n944), .B2(new_n947), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n946), .A2(new_n947), .B1(new_n948), .B2(new_n949), .ZN(G1344gat));
  NOR2_X1   g749(.A1(new_n357), .A2(new_n735), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n925), .B(new_n717), .C1(new_n934), .C2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(KEYINPUT57), .B1(new_n883), .B2(new_n637), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n913), .A2(new_n794), .A3(new_n356), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT122), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT122), .A4(new_n955), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G148gat), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT59), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n804), .B(new_n914), .C1(new_n927), .C2(new_n937), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n403), .A2(KEYINPUT59), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g764(.A1(new_n940), .A2(new_n403), .A3(new_n804), .A4(new_n941), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1345gat));
  OAI21_X1  g766(.A(G155gat), .B1(new_n938), .B2(new_n762), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n258), .A2(new_n203), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n942), .B2(new_n969), .ZN(G1346gat));
  OAI21_X1  g769(.A(G162gat), .B1(new_n938), .B2(new_n765), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n764), .A2(new_n409), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n942), .B2(new_n972), .ZN(G1347gat));
  NOR2_X1   g772(.A1(new_n883), .A2(new_n742), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n668), .A2(new_n595), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n822), .A2(new_n561), .A3(new_n563), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT123), .Z(new_n978));
  OR3_X1    g777(.A1(new_n807), .A2(new_n595), .A3(new_n666), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n979), .A2(KEYINPUT124), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(KEYINPUT124), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n258), .B1(new_n878), .B2(new_n881), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n637), .B1(new_n982), .B2(new_n862), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n980), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(G169gat), .B1(new_n985), .B2(new_n396), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n978), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n978), .A2(KEYINPUT125), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1348gat));
  OAI21_X1  g790(.A(G176gat), .B1(new_n985), .B2(new_n356), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n975), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n804), .A2(new_n564), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(G1349gat));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n996), .B1(new_n985), .B2(new_n762), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n979), .A2(KEYINPUT124), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n998), .A2(new_n983), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n999), .A2(KEYINPUT126), .A3(new_n258), .A4(new_n981), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n997), .A2(new_n537), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n974), .A2(new_n514), .A3(new_n258), .A4(new_n975), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT60), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1001), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1350gat));
  OAI21_X1  g806(.A(G190gat), .B1(new_n985), .B2(new_n765), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1008), .A2(KEYINPUT61), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n1008), .A2(KEYINPUT61), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n764), .A2(new_n513), .ZN(new_n1011));
  OAI22_X1  g810(.A1(new_n1009), .A2(new_n1010), .B1(new_n993), .B2(new_n1011), .ZN(G1351gat));
  NOR3_X1   g811(.A1(new_n807), .A2(new_n595), .A3(new_n794), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n954), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(G197gat), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n1014), .A2(new_n1015), .A3(new_n396), .ZN(new_n1016));
  NOR3_X1   g815(.A1(new_n794), .A2(new_n595), .A3(new_n637), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n974), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g817(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g818(.A(G197gat), .B1(new_n1019), .B2(new_n822), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1016), .A2(new_n1020), .ZN(G1352gat));
  AOI21_X1  g820(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1019), .A2(new_n804), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g822(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1024));
  XNOR2_X1  g823(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  OAI21_X1  g824(.A(G204gat), .B1(new_n1014), .B2(new_n356), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1025), .A2(new_n1026), .ZN(G1353gat));
  OR3_X1    g826(.A1(new_n1018), .A2(G211gat), .A3(new_n762), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n954), .A2(new_n258), .A3(new_n1013), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n1029), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G1354gat));
  OAI21_X1  g831(.A(G218gat), .B1(new_n1014), .B2(new_n765), .ZN(new_n1033));
  OR2_X1    g832(.A1(new_n765), .A2(G218gat), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1033), .B1(new_n1018), .B2(new_n1034), .ZN(G1355gat));
endmodule


