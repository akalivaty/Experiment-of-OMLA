//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n450, new_n451, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n555, new_n557, new_n558, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1154,
    new_n1156, new_n1157, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  INV_X1    g024(.A(G567), .ZN(new_n450));
  NOR2_X1   g025(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G236), .A3(G237), .A4(G235), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n456), .A2(new_n450), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT68), .A4(G125), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(G2105), .ZN(G160));
  NAND2_X1  g052(.A1(new_n465), .A2(new_n467), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n479), .A2(G102), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n493), .B2(new_n479), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n479), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n492), .A2(KEYINPUT4), .A3(G138), .A4(new_n479), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n488), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n489), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(new_n490), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n501), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n504), .A2(KEYINPUT69), .A3(new_n497), .A4(new_n498), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(G164));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(G651), .A2(new_n514), .B1(new_n516), .B2(G50), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n509), .A3(new_n511), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT70), .ZN(new_n519));
  INV_X1    g094(.A(new_n512), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(new_n515), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n517), .B1(new_n523), .B2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  XNOR2_X1  g101(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n527), .A2(new_n529), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(new_n531), .B1(new_n516), .B2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n519), .A2(new_n522), .A3(G89), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n520), .A2(G63), .A3(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n519), .A2(new_n522), .A3(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n516), .A2(G52), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n540), .A2(KEYINPUT72), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT72), .B1(new_n540), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G56), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n512), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(G651), .A2(new_n548), .B1(new_n516), .B2(G43), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n519), .A2(new_n522), .A3(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n515), .A2(G53), .A3(G543), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n519), .A2(new_n522), .A3(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(KEYINPUT74), .B(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n512), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G651), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(new_n562), .A3(new_n566), .ZN(G299));
  NAND3_X1  g142(.A1(new_n519), .A2(new_n522), .A3(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n516), .A2(G49), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g145(.A(KEYINPUT75), .B(G651), .C1(new_n520), .C2(G74), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  AOI21_X1  g147(.A(G74), .B1(new_n509), .B2(new_n511), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n538), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n570), .A2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT76), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n512), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n516), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n519), .A2(new_n522), .A3(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n516), .A2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT77), .B(G85), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n538), .B2(new_n585), .C1(new_n523), .C2(new_n586), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT78), .Z(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n523), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT10), .A4(G92), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n516), .A2(G54), .ZN(new_n596));
  OR2_X1    g171(.A1(KEYINPUT79), .A2(G66), .ZN(new_n597));
  NAND2_X1  g172(.A1(KEYINPUT79), .A2(G66), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n520), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G79), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n508), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n595), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n590), .B1(new_n604), .B2(G868), .ZN(G321));
  XOR2_X1   g180(.A(G321), .B(KEYINPUT80), .Z(G284));
  NAND2_X1  g181(.A1(G286), .A2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G297));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(G868), .ZN(G280));
  XNOR2_X1  g185(.A(KEYINPUT81), .B(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(G860), .B2(new_n611), .ZN(G148));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g191(.A1(G123), .A2(new_n480), .B1(new_n482), .B2(G135), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n620), .B(new_n621), .C1(G111), .C2(new_n479), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n479), .A2(G2104), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n478), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT13), .B(G2100), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n630), .ZN(G156));
  XOR2_X1   g206(.A(KEYINPUT15), .B(G2435), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n637));
  OR2_X1    g212(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n638));
  NAND4_X1  g213(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2443), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(G14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2072), .B(G2078), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT86), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(KEYINPUT17), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT87), .Z(new_n660));
  NOR3_X1   g235(.A1(new_n657), .A2(new_n653), .A3(new_n651), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n653), .A2(new_n654), .A3(new_n650), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT90), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n673), .A2(new_n675), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n671), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(new_n676), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n677), .B1(new_n676), .B2(new_n670), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT21), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1996), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1991), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n686), .B(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n552), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n693), .B2(G19), .ZN(new_n695));
  INV_X1    g270(.A(G1341), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT25), .Z(new_n700));
  AOI22_X1  g275(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n482), .A2(KEYINPUT96), .A3(G139), .ZN(new_n702));
  AOI21_X1  g277(.A(KEYINPUT96), .B1(new_n482), .B2(G139), .ZN(new_n703));
  OAI221_X1 g278(.A(new_n700), .B1(new_n479), .B2(new_n701), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G33), .B(new_n704), .S(G29), .Z(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(G2072), .Z(new_n706));
  OR2_X1    g281(.A1(KEYINPUT24), .A2(G34), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(KEYINPUT24), .A2(G34), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G160), .B2(new_n708), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G2084), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT27), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT97), .ZN(new_n714));
  AOI22_X1  g289(.A1(G129), .A2(new_n480), .B1(new_n482), .B2(G141), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  INV_X1    g292(.A(G105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n717), .C1(new_n718), .C2(new_n625), .ZN(new_n719));
  MUX2_X1   g294(.A(G32), .B(new_n719), .S(G29), .Z(new_n720));
  OAI211_X1 g295(.A(new_n706), .B(new_n712), .C1(new_n714), .C2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT98), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n693), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n693), .ZN(new_n724));
  INV_X1    g299(.A(G1966), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n708), .A2(G35), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G162), .B2(new_n708), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT29), .B(G2090), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n720), .A2(new_n714), .ZN(new_n731));
  INV_X1    g306(.A(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(KEYINPUT31), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n623), .B2(new_n708), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT99), .B(G28), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n708), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT100), .Z(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n731), .B(new_n740), .C1(KEYINPUT31), .C2(new_n732), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n693), .A2(G4), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n604), .B2(new_n693), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n730), .B(new_n741), .C1(G1348), .C2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G26), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n480), .A2(G128), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n482), .A2(G140), .ZN(new_n748));
  NOR2_X1   g323(.A1(G104), .A2(G2105), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(new_n479), .B2(G116), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n746), .B1(new_n751), .B2(G29), .ZN(new_n752));
  MUX2_X1   g327(.A(new_n746), .B(new_n752), .S(KEYINPUT28), .Z(new_n753));
  INV_X1    g328(.A(G2067), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI22_X1  g330(.A1(new_n695), .A2(new_n696), .B1(G2084), .B2(new_n711), .ZN(new_n756));
  NOR2_X1   g331(.A1(G27), .A2(G29), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G164), .B2(G29), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT102), .B(G2078), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n755), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n743), .A2(G1348), .ZN(new_n762));
  AND4_X1   g337(.A1(new_n726), .A2(new_n744), .A3(new_n761), .A4(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT101), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G5), .B2(G16), .ZN(new_n765));
  OR3_X1    g340(.A1(new_n764), .A2(G5), .A3(G16), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n765), .B(new_n766), .C1(G301), .C2(new_n693), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1961), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n693), .A2(G20), .ZN(new_n769));
  OAI211_X1 g344(.A(KEYINPUT23), .B(new_n769), .C1(new_n608), .C2(new_n693), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(KEYINPUT23), .B2(new_n769), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1956), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n722), .A2(new_n763), .A3(new_n768), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n588), .A2(new_n693), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n693), .B2(G24), .ZN(new_n775));
  INV_X1    g350(.A(G1986), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n480), .A2(G119), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n482), .A2(G131), .ZN(new_n779));
  NOR2_X1   g354(.A1(G95), .A2(G2105), .ZN(new_n780));
  OAI21_X1  g355(.A(G2104), .B1(new_n479), .B2(G107), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  MUX2_X1   g357(.A(G25), .B(new_n782), .S(G29), .Z(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT35), .B(G1991), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT93), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n783), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n775), .B2(new_n776), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n693), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(G288), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n693), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT33), .B(G1976), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT94), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n791), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n693), .A2(G22), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n693), .ZN(new_n796));
  INV_X1    g371(.A(G1971), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n693), .A2(G6), .ZN(new_n799));
  INV_X1    g374(.A(G305), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n693), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n794), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n788), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT95), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(KEYINPUT95), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n777), .B(new_n807), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT36), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n808), .B(KEYINPUT95), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n814), .A2(new_n815), .A3(new_n777), .A4(new_n807), .ZN(new_n816));
  AOI211_X1 g391(.A(new_n698), .B(new_n773), .C1(new_n813), .C2(new_n816), .ZN(G311));
  AOI21_X1  g392(.A(new_n773), .B1(new_n813), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(new_n697), .ZN(G150));
  NAND2_X1  g394(.A1(G80), .A2(G543), .ZN(new_n820));
  INV_X1    g395(.A(G67), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n512), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g397(.A1(G651), .A2(new_n822), .B1(new_n516), .B2(G55), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n523), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n604), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(KEYINPUT103), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n823), .B(new_n832), .C1(new_n824), .C2(new_n523), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n552), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n825), .A2(KEYINPUT103), .A3(new_n551), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n830), .B(new_n836), .Z(new_n837));
  OAI21_X1  g412(.A(new_n827), .B1(new_n837), .B2(G860), .ZN(G145));
  NAND3_X1  g413(.A1(new_n504), .A2(new_n497), .A3(new_n498), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(new_n751), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n704), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n719), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n480), .A2(G130), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n482), .A2(G142), .ZN(new_n844));
  NOR2_X1   g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(new_n479), .B2(G118), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n782), .B(new_n847), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n628), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n623), .B(G160), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n486), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n849), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n850), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(G37), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(KEYINPUT104), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n842), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n842), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n854), .B(new_n855), .C1(new_n859), .C2(new_n852), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g436(.A(G868), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n825), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(G288), .A2(new_n800), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(G288), .A2(new_n800), .ZN(new_n866));
  AOI21_X1  g441(.A(G303), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n868), .A2(G166), .A3(new_n864), .ZN(new_n869));
  OAI21_X1  g444(.A(G290), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(G166), .B1(new_n868), .B2(new_n864), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n865), .A2(G303), .A3(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(new_n588), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n874), .A2(KEYINPUT106), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(KEYINPUT42), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT106), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n593), .A2(new_n594), .B1(G651), .B2(new_n601), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n608), .A3(new_n596), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n608), .B1(new_n881), .B2(new_n596), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n603), .A2(G299), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n886), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n883), .A2(new_n884), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n613), .B(new_n836), .ZN(new_n890));
  MUX2_X1   g465(.A(new_n888), .B(new_n889), .S(new_n890), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n879), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n863), .B1(new_n892), .B2(new_n862), .ZN(G295));
  OAI21_X1  g468(.A(new_n863), .B1(new_n892), .B2(new_n862), .ZN(G331));
  NAND2_X1  g469(.A1(G286), .A2(KEYINPUT107), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n532), .A2(new_n533), .A3(new_n896), .A4(new_n534), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n539), .B(new_n897), .C1(new_n542), .C2(new_n543), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n834), .A2(new_n898), .A3(new_n835), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n834), .B2(new_n835), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n895), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n898), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n836), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n895), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n899), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n906), .A3(new_n889), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT109), .ZN(new_n908));
  INV_X1    g483(.A(new_n874), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n885), .A2(new_n887), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n906), .B2(new_n902), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n902), .A2(new_n906), .A3(new_n889), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n908), .B(new_n909), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n902), .A2(new_n906), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n888), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n915), .B(new_n907), .C1(new_n874), .C2(KEYINPUT109), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n855), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(KEYINPUT110), .A3(KEYINPUT43), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n874), .B1(new_n915), .B2(new_n907), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT108), .B1(new_n923), .B2(G37), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n855), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n915), .A2(new_n874), .A3(new_n907), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n924), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT44), .B1(new_n929), .B2(KEYINPUT43), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  AND4_X1   g506(.A1(new_n931), .A2(new_n913), .A3(new_n855), .A4(new_n916), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(new_n929), .B2(KEYINPUT43), .ZN(new_n933));
  OAI22_X1  g508(.A1(new_n922), .A2(new_n930), .B1(new_n933), .B2(KEYINPUT44), .ZN(G397));
  AND2_X1   g509(.A1(new_n497), .A2(new_n498), .ZN(new_n935));
  AOI21_X1  g510(.A(G1384), .B1(new_n935), .B2(new_n504), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT111), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n494), .B2(new_n499), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G160), .A2(G40), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(G1996), .A3(new_n719), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(KEYINPUT112), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n751), .B(G2067), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n719), .A2(G1996), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(KEYINPUT112), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n947), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n782), .A2(new_n785), .ZN(new_n953));
  OAI22_X1  g528(.A1(new_n952), .A2(new_n953), .B1(G2067), .B2(new_n751), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n945), .ZN(new_n955));
  OR2_X1    g530(.A1(new_n943), .A2(new_n944), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n782), .A2(new_n785), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n956), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n588), .A2(new_n776), .A3(new_n945), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT127), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n956), .B2(G1996), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n945), .B1(new_n719), .B2(new_n948), .ZN(new_n968));
  INV_X1    g543(.A(G1996), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n945), .A2(KEYINPUT46), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  OR2_X1    g546(.A1(new_n971), .A2(KEYINPUT125), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(KEYINPUT125), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(KEYINPUT47), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n964), .A2(new_n965), .A3(new_n974), .A4(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n977), .A2(new_n955), .A3(new_n963), .A4(new_n974), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  AOI211_X1 g557(.A(new_n982), .B(new_n470), .C1(new_n476), .C2(G2105), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n942), .B2(new_n939), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n500), .A2(new_n505), .A3(new_n938), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n986), .A2(KEYINPUT113), .A3(new_n942), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT113), .B1(new_n986), .B2(new_n942), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n797), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT114), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n993), .B(new_n938), .C1(new_n494), .C2(new_n499), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n983), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n996), .A2(G2090), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n998), .A3(new_n797), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n991), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  XOR2_X1   g576(.A(new_n1001), .B(KEYINPUT55), .Z(new_n1002));
  AND3_X1   g577(.A1(new_n1000), .A2(G8), .A3(new_n1002), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT118), .B(G1981), .Z(new_n1004));
  NAND3_X1  g579(.A1(new_n581), .A2(new_n582), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1981), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n581), .B2(new_n582), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT49), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1005), .B(new_n1010), .C1(new_n800), .C2(new_n1007), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n983), .A2(new_n936), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT115), .B(G8), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1014), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1012), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n575), .A2(new_n568), .A3(G1976), .A4(new_n569), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1021), .B(new_n1024), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1022), .B(KEYINPUT117), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1018), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(new_n1016), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1019), .B(new_n1025), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT119), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1024), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT52), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(new_n1019), .A4(new_n1025), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1003), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n790), .A2(new_n1020), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT120), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1005), .B1(new_n1038), .B2(new_n1012), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1002), .B1(new_n1000), .B2(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1015), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n500), .A2(new_n505), .A3(KEYINPUT45), .A4(new_n938), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n939), .A2(new_n942), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n983), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n725), .ZN(new_n1047));
  INV_X1    g622(.A(G2084), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n992), .A2(new_n995), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1043), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G168), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1041), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT63), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1036), .B(new_n1040), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n992), .A2(new_n1048), .A3(new_n995), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT45), .B1(new_n839), .B2(new_n938), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1056), .A2(new_n944), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1966), .B1(new_n1057), .B2(new_n1044), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1015), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n1059), .B2(KEYINPUT123), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G286), .A2(new_n1015), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1062), .B1(new_n1050), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n983), .A2(new_n994), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1065), .B1(KEYINPUT50), .B2(new_n986), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1066), .A2(new_n1048), .B1(new_n1046), .B2(new_n725), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1061), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1060), .A2(new_n1064), .B1(KEYINPUT51), .B2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1067), .A2(new_n1061), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT62), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT124), .B(G1961), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G2078), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(new_n985), .C1(new_n987), .C2(new_n988), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(G2078), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1057), .A2(new_n1080), .A3(new_n1044), .ZN(new_n1081));
  AOI21_X1  g656(.A(G301), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1068), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1083));
  OAI21_X1  g658(.A(KEYINPUT51), .B1(new_n1083), .B2(new_n1062), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1061), .B1(new_n1059), .B2(KEYINPUT123), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1050), .B2(new_n1063), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1084), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1071), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1072), .A2(new_n1082), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1050), .A2(new_n1053), .A3(G168), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n939), .A2(KEYINPUT50), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n500), .A2(new_n505), .A3(new_n993), .A4(new_n938), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n983), .B(new_n1094), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1956), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT56), .B(G2072), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n985), .B(new_n1101), .C1(new_n987), .C2(new_n988), .ZN(new_n1102));
  XOR2_X1   g677(.A(G299), .B(KEYINPUT57), .Z(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1066), .A2(G1348), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1013), .A2(G2067), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n604), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1104), .B(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1348), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n996), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1106), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n604), .A4(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n969), .B(new_n985), .C1(new_n987), .C2(new_n988), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1013), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n551), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1122), .B2(KEYINPUT59), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1115), .A2(new_n603), .A3(new_n1117), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1116), .B1(new_n1107), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1126), .B(new_n551), .C1(new_n1119), .C2(new_n1121), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1111), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n985), .A2(new_n943), .A3(new_n1080), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1079), .A2(G301), .A3(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1130), .B1(new_n1132), .B2(new_n1082), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1079), .A2(G301), .A3(new_n1081), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1131), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1075), .B(new_n1136), .C1(new_n1078), .C2(new_n1077), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1135), .B(KEYINPUT54), .C1(new_n1137), .C2(G301), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1133), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1092), .B(new_n1093), .C1(new_n1129), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n1141));
  AOI21_X1  g716(.A(G2090), .B1(new_n1098), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1141), .B2(new_n1098), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n990), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1002), .B1(new_n1144), .B2(new_n1015), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1145), .A2(new_n1003), .A3(new_n1030), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1054), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n588), .B(G1986), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n959), .B1(new_n956), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n981), .B1(new_n1147), .B2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g725(.A1(new_n860), .A2(new_n648), .A3(new_n667), .ZN(new_n1152));
  NOR2_X1   g726(.A1(G229), .A2(new_n462), .ZN(new_n1153));
  INV_X1    g727(.A(new_n1153), .ZN(new_n1154));
  NOR3_X1   g728(.A1(new_n933), .A2(new_n1152), .A3(new_n1154), .ZN(G308));
  NAND2_X1  g729(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n1156));
  INV_X1    g730(.A(new_n932), .ZN(new_n1157));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g732(.A1(G401), .A2(G227), .ZN(new_n1159));
  NAND4_X1  g733(.A1(new_n1158), .A2(new_n860), .A3(new_n1153), .A4(new_n1159), .ZN(G225));
endmodule


