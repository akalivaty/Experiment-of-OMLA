//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(new_n193), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n189), .B(new_n194), .C1(new_n197), .C2(new_n191), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G110), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(new_n189), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT24), .B(G110), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G125), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n203), .A2(new_n205), .A3(KEYINPUT80), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n204), .A2(KEYINPUT80), .A3(G140), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n203), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n208), .B2(new_n211), .ZN(new_n214));
  OAI221_X1 g028(.A(new_n199), .B1(new_n200), .B2(new_n201), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n214), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n203), .A2(new_n205), .A3(new_n209), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n198), .A2(G110), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n200), .A2(new_n201), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n216), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G137), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n223), .B(new_n225), .Z(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n215), .A2(new_n221), .A3(new_n226), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n187), .B1(new_n230), .B2(G902), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n228), .A2(KEYINPUT25), .A3(new_n232), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(G234), .B2(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(G902), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n229), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT74), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n209), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(KEYINPUT70), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n243), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT65), .B1(new_n209), .B2(G143), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n248), .A2(G128), .B1(new_n253), .B2(new_n243), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(G146), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n243), .A2(new_n255), .A3(G128), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n246), .A2(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n242), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n243), .A2(new_n255), .A3(G128), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT70), .B(KEYINPUT1), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n190), .B1(new_n259), .B2(new_n243), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n251), .A2(G146), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n249), .B2(new_n252), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n264), .B(KEYINPUT74), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G137), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n272));
  INV_X1    g086(.A(G137), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G134), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n276));
  OAI21_X1  g090(.A(G131), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g092(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT66), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n280), .A2(new_n281), .B1(new_n273), .B2(G134), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g097(.A1(KEYINPUT11), .A2(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G137), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n273), .A2(KEYINPUT67), .A3(KEYINPUT11), .A4(G134), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n279), .A2(new_n282), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(G131), .B1(new_n270), .B2(G137), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n278), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n286), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n280), .A2(new_n281), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(new_n274), .A3(new_n279), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n290), .A2(new_n278), .A3(new_n292), .A4(new_n288), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n277), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n290), .A2(new_n292), .A3(new_n288), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n290), .A2(new_n292), .A3(new_n271), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n297), .A2(new_n293), .B1(G131), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT0), .B(G128), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT0), .A2(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n243), .A2(new_n255), .ZN(new_n302));
  OAI22_X1  g116(.A1(new_n267), .A2(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI22_X1  g117(.A1(new_n269), .A2(new_n295), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G116), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT71), .B1(new_n305), .B2(G119), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n188), .A3(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(G119), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT2), .B(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n313));
  XOR2_X1   g127(.A(KEYINPUT2), .B(G113), .Z(new_n314));
  AOI21_X1  g128(.A(KEYINPUT72), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n310), .A2(new_n316), .A3(new_n311), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n312), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT73), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n305), .A2(KEYINPUT71), .A3(G119), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n188), .A2(G116), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n322), .A2(KEYINPUT72), .A3(new_n314), .A4(new_n306), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n316), .B1(new_n310), .B2(new_n311), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n312), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT75), .B1(new_n304), .B2(new_n328), .ZN(new_n329));
  AOI221_X4 g143(.A(KEYINPUT73), .B1(new_n311), .B2(new_n310), .C1(new_n323), .C2(new_n324), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n326), .B1(new_n325), .B2(new_n312), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n298), .A2(G131), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n289), .B2(new_n294), .ZN(new_n335));
  INV_X1    g149(.A(new_n303), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n297), .A2(new_n293), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n338), .A2(new_n261), .A3(new_n277), .A4(new_n268), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n332), .A2(new_n333), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n304), .A2(new_n328), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n329), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT28), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n344));
  NOR2_X1   g158(.A1(G237), .A2(G953), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G210), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT27), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT26), .B(G101), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n332), .A2(new_n337), .A3(new_n339), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n344), .B(new_n350), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n343), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n264), .B1(new_n265), .B2(new_n267), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n277), .B(new_n356), .C1(new_n289), .C2(new_n294), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n303), .B1(new_n338), .B2(new_n334), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n337), .A2(new_n339), .A3(KEYINPUT30), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n328), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n329), .A3(new_n340), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n350), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n344), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n351), .A2(new_n352), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n349), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n328), .B1(new_n359), .B2(new_n358), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n329), .A2(new_n368), .A3(new_n340), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n367), .B1(KEYINPUT28), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n354), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT77), .B1(new_n371), .B2(G472), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT77), .ZN(new_n373));
  INV_X1    g187(.A(G472), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(KEYINPUT28), .ZN(new_n375));
  INV_X1    g189(.A(new_n367), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n363), .B2(new_n350), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI211_X1 g193(.A(new_n373), .B(new_n374), .C1(new_n379), .C2(new_n354), .ZN(new_n380));
  NOR2_X1   g194(.A1(G472), .A2(G902), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n362), .A2(new_n329), .A3(new_n340), .A4(new_n349), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n383), .A2(KEYINPUT76), .A3(KEYINPUT31), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT76), .B1(new_n383), .B2(KEYINPUT31), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n375), .A2(new_n366), .ZN(new_n388));
  INV_X1    g202(.A(new_n383), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT31), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n388), .A2(new_n350), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n382), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  OAI22_X1  g206(.A1(new_n372), .A2(new_n380), .B1(new_n392), .B2(KEYINPUT32), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT32), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n382), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n383), .A2(KEYINPUT31), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n384), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n351), .A2(new_n352), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(new_n369), .B2(KEYINPUT28), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n401), .A2(new_n349), .B1(KEYINPUT31), .B2(new_n383), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n395), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT78), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(new_n395), .C1(new_n399), .C2(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n241), .B1(new_n393), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(G469), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G128), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n262), .A2(new_n263), .B1(new_n414), .B2(new_n302), .ZN(new_n415));
  INV_X1    g229(.A(G104), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT3), .B1(new_n416), .B2(G107), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT3), .ZN(new_n418));
  INV_X1    g232(.A(G107), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n418), .A2(new_n419), .A3(G104), .ZN(new_n420));
  INV_X1    g234(.A(G101), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(G107), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n416), .A2(G107), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n419), .A2(G104), .ZN(new_n425));
  OAI21_X1  g239(.A(G101), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT81), .B1(new_n415), .B2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n423), .A2(new_n426), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n243), .A2(new_n255), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n190), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n431), .A2(new_n432), .B1(new_n256), .B2(new_n259), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n267), .ZN(new_n435));
  OAI21_X1  g249(.A(G128), .B1(new_n263), .B2(new_n266), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n260), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n428), .A2(new_n434), .B1(new_n437), .B2(new_n427), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n411), .B(new_n412), .C1(new_n438), .C2(new_n299), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n427), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n415), .A2(new_n427), .A3(KEYINPUT81), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n430), .B1(new_n429), .B2(new_n433), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n443), .A2(KEYINPUT83), .A3(new_n410), .A4(new_n335), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n439), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n439), .B2(new_n444), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G140), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n224), .A2(G227), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT10), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n441), .B2(new_n442), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n417), .A2(new_n420), .A3(new_n422), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT4), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(new_n455), .A3(G101), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(G101), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT4), .A3(new_n423), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n336), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n261), .A2(KEYINPUT10), .A3(new_n268), .A4(new_n429), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n335), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n299), .A2(KEYINPUT82), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n451), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n446), .A2(new_n447), .A3(new_n466), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n453), .A2(new_n459), .A3(new_n460), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n463), .A2(new_n464), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n461), .A2(new_n335), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n451), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n409), .B(new_n232), .C1(new_n467), .C2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n409), .A2(new_n232), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n450), .B1(new_n468), .B2(new_n469), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n439), .B(new_n444), .C1(new_n461), .C2(new_n465), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n471), .A2(new_n475), .B1(new_n476), .B2(new_n450), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n474), .B1(new_n477), .B2(G469), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G221), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT9), .B(G234), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n480), .B1(new_n482), .B2(new_n232), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT90), .ZN(new_n485));
  INV_X1    g299(.A(G237), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n224), .A3(G214), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n251), .ZN(new_n488));
  AOI21_X1  g302(.A(G143), .B1(new_n345), .B2(G214), .ZN(new_n489));
  OAI211_X1 g303(.A(KEYINPUT18), .B(G131), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n251), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n345), .A2(G143), .A3(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT18), .A2(G131), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n204), .A2(KEYINPUT80), .A3(G140), .ZN(new_n496));
  XNOR2_X1  g310(.A(G125), .B(G140), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(KEYINPUT80), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n217), .B1(new_n498), .B2(G146), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n485), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n206), .A2(new_n207), .A3(G146), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n218), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n502), .A2(new_n490), .A3(KEYINPUT90), .A4(new_n494), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n416), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n508));
  INV_X1    g322(.A(G131), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n491), .A2(new_n509), .A3(new_n492), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n491), .B2(new_n492), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT19), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n497), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n206), .A2(new_n207), .B1(new_n497), .B2(KEYINPUT92), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n209), .B(new_n516), .C1(new_n517), .C2(new_n515), .ZN(new_n518));
  OAI21_X1  g332(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(KEYINPUT91), .A3(new_n510), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n216), .A2(new_n513), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n504), .A2(new_n507), .A3(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(G475), .A2(G902), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT93), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n525), .A3(new_n510), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n512), .A2(KEYINPUT17), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n213), .A2(new_n214), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n528), .A2(new_n529), .B1(new_n500), .B2(new_n503), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n522), .B(new_n524), .C1(new_n530), .C2(new_n507), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT20), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n216), .A2(new_n526), .A3(new_n212), .A4(new_n527), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n504), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n506), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT20), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n522), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n535), .A2(new_n537), .A3(new_n522), .A4(new_n524), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n532), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n535), .A2(new_n522), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n541), .A2(new_n536), .A3(new_n537), .A4(new_n524), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n507), .A2(KEYINPUT95), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n504), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n232), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n504), .B2(new_n533), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT96), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n543), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT96), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n549), .A2(new_n550), .A3(new_n232), .A4(new_n545), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(G475), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n540), .A2(new_n542), .A3(new_n552), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n481), .A2(new_n235), .A3(G953), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n305), .A2(G122), .ZN(new_n556));
  INV_X1    g370(.A(G122), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G116), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(G107), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n558), .A3(new_n419), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n251), .A2(G128), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n190), .A2(G143), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(new_n270), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n560), .A2(new_n561), .B1(KEYINPUT98), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n564), .A2(KEYINPUT98), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n563), .B1(new_n562), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n190), .A2(G143), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT97), .B1(new_n570), .B2(KEYINPUT13), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n562), .A2(new_n572), .A3(new_n568), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(new_n270), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n564), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n270), .B1(new_n562), .B2(new_n563), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n561), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT99), .B1(new_n556), .B2(KEYINPUT14), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT14), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n305), .A4(G122), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n556), .A2(KEYINPUT14), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n580), .A2(new_n583), .A3(new_n558), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n579), .B1(G107), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n555), .B1(new_n576), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n565), .B(new_n566), .C1(new_n270), .C2(new_n574), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n585), .A2(G107), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n589), .B(new_n554), .C1(new_n590), .C2(new_n579), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT100), .B(new_n555), .C1(new_n576), .C2(new_n586), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n594), .A2(KEYINPUT101), .A3(new_n232), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT102), .B(G952), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(G953), .ZN(new_n600));
  NAND2_X1  g414(.A1(G234), .A2(G237), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(G902), .A3(G953), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT103), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT21), .B(G898), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n592), .A2(KEYINPUT101), .A3(new_n232), .A4(new_n593), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n596), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n598), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n553), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n479), .A2(new_n484), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(G110), .B(G122), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n458), .A2(new_n456), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n319), .B2(new_n327), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n313), .A2(KEYINPUT5), .ZN(new_n619));
  INV_X1    g433(.A(G113), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n305), .A2(G119), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT5), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n323), .A2(new_n324), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n429), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n616), .B1(new_n618), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n617), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n330), .B2(new_n331), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n625), .A3(new_n615), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n627), .A2(KEYINPUT6), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n303), .A2(G125), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT85), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n437), .A2(new_n204), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT85), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n303), .A2(new_n635), .A3(G125), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n633), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G224), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(G953), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT86), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n637), .B(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT6), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(new_n616), .C1(new_n618), .C2(new_n626), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n631), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT87), .B(KEYINPUT8), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n615), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n623), .B1(new_n310), .B2(new_n622), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n325), .A2(KEYINPUT88), .A3(new_n429), .A4(new_n647), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n648), .B1(new_n429), .B2(new_n624), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT88), .B1(new_n624), .B2(new_n429), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT7), .B1(new_n638), .B2(G953), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n633), .A2(new_n634), .A3(new_n636), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n632), .B1(G125), .B2(new_n356), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n652), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n630), .A2(new_n651), .A3(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n232), .ZN(new_n659));
  OAI21_X1  g473(.A(G210), .B1(G237), .B2(G902), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n644), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT89), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n644), .A2(new_n659), .A3(new_n660), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n644), .B2(new_n659), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n666), .B2(new_n662), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n668));
  OAI21_X1  g482(.A(G214), .B1(G237), .B2(G902), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n614), .A2(new_n667), .A3(new_n668), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n644), .A2(new_n659), .ZN(new_n671));
  INV_X1    g485(.A(new_n660), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n662), .A3(new_n661), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n664), .A2(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n674), .A2(new_n669), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n483), .B1(new_n473), .B2(new_n478), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n613), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT104), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n670), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n408), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n421), .ZN(G3));
  NAND2_X1  g496(.A1(new_n388), .A2(new_n350), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n389), .A2(new_n390), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n398), .A4(new_n384), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n374), .B1(new_n685), .B2(new_n232), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n392), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n479), .A2(new_n484), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n240), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n669), .B(new_n609), .C1(new_n664), .C2(new_n665), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n594), .A2(new_n232), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n595), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT33), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n594), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n587), .A2(KEYINPUT33), .A3(new_n591), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n232), .A2(G478), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n553), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n691), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n690), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n416), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT105), .B(KEYINPUT34), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G6));
  AND2_X1   g519(.A1(new_n598), .A2(new_n611), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n691), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n532), .A2(new_n539), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n552), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n690), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT35), .B(G107), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G9));
  NOR2_X1   g527(.A1(new_n227), .A2(KEYINPUT36), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n222), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n238), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n237), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n686), .A2(new_n392), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n670), .A3(new_n679), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT37), .B(G110), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT106), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G12));
  NAND2_X1  g537(.A1(new_n371), .A2(G472), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n373), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n371), .A2(KEYINPUT77), .A3(G472), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n685), .A2(new_n381), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n394), .ZN(new_n728));
  INV_X1    g542(.A(new_n406), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n405), .B1(new_n685), .B2(new_n395), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n718), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n669), .B1(new_n664), .B2(new_n665), .ZN(new_n733));
  INV_X1    g547(.A(G900), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n603), .B1(new_n734), .B2(new_n606), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n709), .A2(new_n736), .ZN(new_n737));
  NOR4_X1   g551(.A1(new_n688), .A2(new_n733), .A3(new_n706), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G128), .ZN(G30));
  NAND2_X1  g554(.A1(new_n674), .A2(new_n675), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n553), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n706), .ZN(new_n745));
  INV_X1    g559(.A(new_n669), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n717), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n735), .B(KEYINPUT39), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n688), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT40), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n745), .B(new_n747), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n743), .B(new_n751), .C1(new_n750), .C2(new_n749), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n363), .A2(new_n349), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n754), .B(new_n232), .C1(new_n349), .C2(new_n342), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n727), .A2(new_n394), .B1(G472), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n731), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(G472), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n392), .B2(KEYINPUT32), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT108), .B1(new_n407), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n752), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n752), .A2(new_n764), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n251), .ZN(G45));
  AND2_X1   g581(.A1(new_n699), .A2(new_n553), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n736), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n769), .A2(new_n688), .A3(new_n733), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n770), .B(new_n717), .C1(new_n393), .C2(new_n407), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT110), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n725), .A2(new_n726), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n727), .A2(new_n394), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n404), .A3(new_n406), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n717), .A4(new_n770), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G146), .ZN(G48));
  NAND2_X1  g593(.A1(new_n470), .A2(new_n471), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n450), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n439), .A2(new_n444), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n475), .B1(new_n782), .B2(new_n445), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n781), .B1(new_n783), .B2(new_n446), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n232), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(G469), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n484), .A3(new_n473), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n241), .B(new_n788), .C1(new_n393), .C2(new_n407), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n701), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT41), .B(G113), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G15));
  OAI21_X1  g606(.A(KEYINPUT111), .B1(new_n789), .B2(new_n710), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n240), .B1(new_n728), .B2(new_n731), .ZN(new_n794));
  INV_X1    g608(.A(new_n710), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n796), .A4(new_n788), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G116), .ZN(G18));
  NOR4_X1   g613(.A1(new_n787), .A2(new_n553), .A3(new_n612), .A4(new_n733), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n800), .B(new_n717), .C1(new_n407), .C2(new_n393), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G119), .ZN(G21));
  OAI21_X1  g616(.A(new_n232), .B1(new_n399), .B2(new_n402), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(G472), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n343), .A2(KEYINPUT112), .A3(new_n366), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n350), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT112), .B1(new_n343), .B2(new_n366), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n684), .B(new_n396), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n381), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n804), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n787), .A2(new_n744), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n241), .A3(new_n707), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G122), .ZN(G24));
  NOR2_X1   g627(.A1(new_n700), .A2(new_n735), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n804), .A2(new_n809), .A3(new_n717), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n816));
  INV_X1    g630(.A(new_n733), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n788), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n804), .A2(new_n809), .A3(new_n717), .A4(new_n814), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n788), .A2(new_n817), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT113), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G125), .ZN(G27));
  NOR3_X1   g637(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT89), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n669), .B(new_n484), .C1(new_n824), .C2(new_n663), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n479), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n473), .A2(new_n478), .A3(KEYINPUT114), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n775), .A2(new_n241), .A3(new_n814), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT115), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT42), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n831), .B2(KEYINPUT115), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n240), .B1(new_n728), .B2(new_n403), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n830), .A2(KEYINPUT42), .A3(new_n814), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n833), .A2(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(G131), .ZN(G33));
  NOR2_X1   g654(.A1(new_n737), .A2(new_n706), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n775), .A2(new_n241), .A3(new_n841), .A4(new_n830), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G134), .ZN(G36));
  NAND2_X1  g657(.A1(new_n741), .A2(new_n669), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n744), .A2(new_n699), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT43), .Z(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n717), .C1(new_n392), .C2(new_n686), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT44), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(G469), .B1(new_n477), .B2(KEYINPUT45), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n477), .A2(KEYINPUT45), .ZN(new_n851));
  OAI22_X1  g665(.A1(new_n850), .A2(new_n851), .B1(new_n409), .B2(new_n232), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT46), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n473), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n484), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n748), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n849), .B(new_n858), .C1(new_n848), .C2(new_n847), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(G137), .ZN(G39));
  XNOR2_X1  g674(.A(new_n857), .B(KEYINPUT47), .ZN(new_n861));
  INV_X1    g675(.A(new_n844), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n240), .A3(new_n814), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n861), .A2(new_n775), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n202), .ZN(G42));
  NOR2_X1   g679(.A1(new_n761), .A2(new_n240), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n786), .A2(new_n473), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n867), .A2(KEYINPUT49), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(KEYINPUT49), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n744), .A2(new_n699), .A3(new_n669), .A4(new_n484), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n866), .A2(new_n743), .A3(new_n871), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n818), .A2(new_n821), .B1(new_n732), .B2(new_n738), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n733), .A2(new_n744), .A3(new_n706), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n717), .A2(new_n483), .A3(new_n735), .ZN(new_n875));
  AND4_X1   g689(.A1(new_n827), .A2(new_n874), .A3(new_n828), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n761), .A2(new_n876), .ZN(new_n877));
  AND4_X1   g691(.A1(KEYINPUT52), .A2(new_n873), .A3(new_n778), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n772), .A2(new_n777), .B1(new_n761), .B2(new_n876), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(new_n879), .B2(new_n873), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n737), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(new_n706), .A3(new_n717), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n844), .A2(new_n688), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n775), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n815), .A2(new_n830), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n842), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n676), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n553), .A2(new_n706), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n608), .B1(new_n889), .B2(new_n700), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n687), .A2(new_n888), .A3(new_n689), .A4(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n720), .B(new_n891), .C1(new_n408), .C2(new_n680), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n801), .B(new_n812), .C1(new_n789), .C2(new_n701), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n797), .B2(new_n793), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n839), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n881), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT53), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT53), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n881), .B2(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n837), .A2(new_n838), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n775), .A2(new_n241), .A3(new_n814), .A4(new_n830), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT42), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n906), .B2(new_n832), .ZN(new_n907));
  INV_X1    g721(.A(new_n790), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n798), .A2(new_n908), .A3(new_n801), .A4(new_n812), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT117), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n892), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n885), .A2(new_n886), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n842), .A4(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT116), .B1(new_n887), .B2(new_n892), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n914), .A2(KEYINPUT53), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n873), .A2(new_n778), .A3(new_n877), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT52), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n873), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT117), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n839), .A2(new_n922), .A3(new_n895), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n910), .A2(new_n916), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n900), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n902), .B1(KEYINPUT54), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n825), .A2(new_n602), .A3(new_n867), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n846), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT119), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n929), .A2(new_n717), .A3(new_n810), .ZN(new_n930));
  AND4_X1   g744(.A1(new_n241), .A2(new_n846), .A3(new_n810), .A4(new_n603), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(new_n746), .A3(new_n743), .A4(new_n788), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT50), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n866), .A2(new_n927), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n699), .A2(new_n553), .ZN(new_n935));
  AOI211_X1 g749(.A(new_n930), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n786), .A2(new_n483), .A3(new_n473), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT118), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n861), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n931), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(new_n844), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT51), .B1(new_n936), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n861), .A2(new_n937), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n941), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n936), .A2(KEYINPUT51), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n600), .B1(new_n940), .B2(new_n820), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n934), .B2(new_n768), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n929), .A2(new_n836), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT120), .Z(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT48), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(KEYINPUT48), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n946), .A2(new_n948), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n926), .A2(new_n943), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(G952), .A2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n872), .B1(new_n954), .B2(new_n955), .ZN(G75));
  NOR2_X1   g770(.A1(new_n224), .A2(G952), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n232), .B1(new_n924), .B2(new_n900), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT56), .B1(new_n959), .B2(G210), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n631), .A2(new_n643), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n641), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT55), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n958), .B1(new_n960), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n960), .B2(new_n963), .ZN(G51));
  XNOR2_X1  g779(.A(new_n925), .B(KEYINPUT54), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n474), .B(KEYINPUT57), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n784), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n851), .A2(new_n850), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n959), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n957), .B1(new_n969), .B2(new_n971), .ZN(G54));
  AND3_X1   g786(.A1(new_n959), .A2(KEYINPUT58), .A3(G475), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n958), .B1(new_n973), .B2(new_n541), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n541), .B2(new_n973), .ZN(G60));
  INV_X1    g789(.A(new_n697), .ZN(new_n976));
  NAND2_X1  g790(.A1(G478), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT59), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n976), .B1(new_n926), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n966), .A2(new_n976), .A3(new_n978), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n979), .A2(new_n980), .A3(new_n957), .ZN(G63));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(G217), .A2(G902), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT60), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT121), .B1(new_n925), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT121), .ZN(new_n987));
  AOI211_X1 g801(.A(new_n987), .B(new_n984), .C1(new_n924), .C2(new_n900), .ZN(new_n988));
  OAI211_X1 g802(.A(KEYINPUT122), .B(new_n715), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n925), .A2(new_n985), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n987), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n925), .A2(KEYINPUT121), .A3(new_n985), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n230), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n989), .A2(new_n993), .A3(new_n958), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n991), .A2(new_n992), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT122), .B1(new_n995), .B2(new_n715), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n982), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n993), .A2(KEYINPUT123), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n715), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT123), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n991), .A2(new_n1000), .A3(new_n230), .A4(new_n992), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n957), .A2(new_n982), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n997), .A2(new_n1003), .ZN(G66));
  OAI21_X1  g818(.A(G953), .B1(new_n607), .B2(new_n638), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n909), .A2(new_n892), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1005), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n961), .B1(G898), .B2(new_n224), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G69));
  NAND3_X1  g823(.A1(new_n859), .A2(new_n778), .A3(new_n873), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT126), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n858), .A2(new_n836), .A3(new_n874), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n842), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n907), .A2(new_n864), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(G953), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n224), .A2(G900), .ZN(new_n1017));
  OR3_X1    g831(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n360), .A2(new_n361), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n516), .B1(new_n517), .B2(new_n515), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1016), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n889), .A2(new_n700), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n862), .A2(new_n749), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n859), .B1(new_n408), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1026), .A2(new_n864), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n763), .A2(new_n765), .A3(new_n778), .A4(new_n873), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT62), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT124), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n1028), .A2(new_n1031), .A3(KEYINPUT62), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1031), .B1(new_n1028), .B2(KEYINPUT62), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1021), .B1(new_n1034), .B2(new_n224), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1035), .A2(KEYINPUT125), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n224), .B1(G227), .B2(G900), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1023), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1037), .B1(new_n1023), .B2(new_n1036), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  OAI211_X1 g854(.A(new_n1030), .B(new_n1006), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1041));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  AOI21_X1  g857(.A(new_n754), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n363), .A2(new_n349), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  AND4_X1   g860(.A1(new_n754), .A2(new_n901), .A3(new_n1043), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n1011), .A2(new_n1006), .A3(new_n1014), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1046), .B1(new_n1048), .B2(new_n1043), .ZN(new_n1049));
  NOR4_X1   g863(.A1(new_n1044), .A2(new_n1047), .A3(new_n957), .A4(new_n1049), .ZN(G57));
endmodule


