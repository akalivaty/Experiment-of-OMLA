//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G469), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT12), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n192), .A2(KEYINPUT80), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(KEYINPUT80), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .A4(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(KEYINPUT1), .A3(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(new_n201), .C1(G128), .C2(new_n202), .ZN(new_n203));
  OR2_X1    g017(.A1(KEYINPUT79), .A2(G104), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT79), .A2(G104), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n204), .B(new_n205), .C1(KEYINPUT3), .C2(G107), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT3), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT3), .A2(G107), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(G104), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G107), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(new_n212), .A3(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n213), .B(G101), .C1(new_n214), .C2(new_n212), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n203), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n200), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  AOI21_X1  g032(.A(G128), .B1(new_n196), .B2(new_n198), .ZN(new_n219));
  INV_X1    g033(.A(new_n201), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(KEYINPUT67), .B(new_n201), .C1(new_n202), .C2(G128), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n211), .A2(new_n215), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n216), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT65), .B(G131), .Z(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n227));
  INV_X1    g041(.A(G134), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(G137), .ZN(new_n229));
  NOR2_X1   g043(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G137), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n233), .B2(G134), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(new_n228), .A3(G137), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(G134), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n230), .ZN(new_n239));
  AND4_X1   g053(.A1(new_n226), .A2(new_n232), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G131), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n234), .A2(new_n236), .B1(new_n238), .B2(new_n230), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(new_n232), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n193), .B(new_n194), .C1(new_n225), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n224), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n203), .A2(new_n211), .A3(new_n215), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n244), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(KEYINPUT80), .A3(new_n192), .A4(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT10), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n224), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n221), .A2(new_n222), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n200), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n210), .B1(new_n206), .B2(new_n209), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n202), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n260), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n264), .B2(new_n202), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n211), .A2(KEYINPUT4), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n259), .B(new_n265), .C1(new_n266), .C2(new_n257), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n247), .A2(new_n252), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n256), .A2(new_n244), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(G110), .B(G140), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n270), .B(KEYINPUT78), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n272), .A2(G227), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n271), .B(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT81), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n269), .A2(KEYINPUT81), .A3(new_n274), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n251), .A2(KEYINPUT82), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n256), .A2(new_n267), .A3(new_n268), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n249), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n269), .ZN(new_n282));
  INV_X1    g096(.A(new_n274), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n245), .A2(new_n250), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT81), .B1(new_n269), .B2(new_n274), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT82), .B1(new_n288), .B2(new_n278), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n191), .B(new_n189), .C1(new_n285), .C2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n191), .A2(new_n189), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n251), .A2(new_n269), .ZN(new_n292));
  INV_X1    g106(.A(new_n275), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n292), .A2(new_n283), .B1(new_n293), .B2(new_n281), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n294), .B2(G469), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n190), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G113), .B(G122), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(new_n214), .ZN(new_n298));
  XNOR2_X1  g112(.A(G125), .B(G140), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n299), .A2(KEYINPUT19), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(KEYINPUT19), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n195), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(KEYINPUT16), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n305), .A2(KEYINPUT16), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(G146), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n272), .A3(G214), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(new_n197), .ZN(new_n311));
  NOR2_X1   g125(.A1(G237), .A2(G953), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n312), .B(G214), .C1(KEYINPUT88), .C2(G143), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n226), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n226), .A3(new_n313), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n302), .B(new_n307), .C1(new_n314), .C2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n299), .B2(new_n195), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  AND4_X1   g135(.A1(new_n318), .A2(new_n305), .A3(new_n321), .A4(new_n195), .ZN(new_n322));
  OAI22_X1  g136(.A1(new_n319), .A2(new_n322), .B1(new_n195), .B2(new_n299), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT18), .A2(G131), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n311), .A2(new_n324), .A3(new_n313), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n311), .A2(new_n313), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT18), .A3(G131), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n298), .B1(new_n317), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n303), .A2(new_n306), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n195), .ZN(new_n331));
  INV_X1    g145(.A(new_n226), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n326), .A2(KEYINPUT17), .A3(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(new_n333), .A3(new_n307), .ZN(new_n334));
  INV_X1    g148(.A(new_n314), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT17), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n315), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n327), .A2(new_n325), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n334), .A2(new_n337), .B1(new_n338), .B2(new_n323), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n329), .B1(new_n339), .B2(new_n298), .ZN(new_n340));
  NOR2_X1   g154(.A1(G475), .A2(G902), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n334), .A2(new_n337), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n298), .A3(new_n328), .ZN(new_n345));
  INV_X1    g159(.A(new_n329), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n341), .ZN(new_n349));
  INV_X1    g163(.A(new_n345), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n298), .B1(new_n344), .B2(new_n328), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n189), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n343), .A2(new_n349), .B1(new_n352), .B2(G475), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n197), .A2(G128), .ZN(new_n355));
  INV_X1    g169(.A(G128), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G143), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(new_n228), .ZN(new_n359));
  INV_X1    g173(.A(G122), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G116), .ZN(new_n361));
  INV_X1    g175(.A(G116), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G122), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G116), .B(G122), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT89), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n212), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n362), .A2(KEYINPUT14), .A3(G122), .ZN(new_n370));
  OAI211_X1 g184(.A(G107), .B(new_n370), .C1(new_n364), .C2(KEYINPUT14), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n359), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n365), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(KEYINPUT89), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(G107), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n358), .A2(new_n228), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT13), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n357), .B1(new_n355), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n355), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT90), .B1(new_n380), .B2(KEYINPUT13), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n355), .A2(new_n382), .A3(new_n378), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n379), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n377), .B1(new_n384), .B2(new_n228), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n372), .B1(new_n376), .B2(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT71), .B(G217), .Z(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n188), .A3(new_n272), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n388), .B(KEYINPUT91), .Z(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT92), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n389), .B(new_n372), .C1(new_n376), .C2(new_n385), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n386), .A2(new_n390), .A3(KEYINPUT92), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n189), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n394), .A2(new_n189), .A3(new_n395), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G952), .ZN(new_n403));
  AOI211_X1 g217(.A(G953), .B(new_n403), .C1(G234), .C2(G237), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n189), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT21), .B(G898), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n354), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT86), .Z(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(KEYINPUT87), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n265), .A2(G125), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n223), .B2(G125), .ZN(new_n413));
  INV_X1    g227(.A(G224), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G953), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n413), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT2), .B(G113), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G116), .B(G119), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n419), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n259), .B(new_n423), .C1(new_n266), .C2(new_n257), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(KEYINPUT5), .ZN(new_n425));
  NOR3_X1   g239(.A1(new_n362), .A2(KEYINPUT5), .A3(G119), .ZN(new_n426));
  INV_X1    g240(.A(G113), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n211), .A2(new_n215), .A3(new_n429), .A4(new_n420), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G122), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n424), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT6), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n430), .ZN(new_n434));
  XOR2_X1   g248(.A(new_n431), .B(KEYINPUT83), .Z(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(KEYINPUT6), .A3(new_n435), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n416), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT7), .B1(new_n414), .B2(G953), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n412), .B(new_n440), .C1(new_n223), .C2(G125), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT85), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n429), .A2(new_n420), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n224), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n430), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n431), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n440), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n413), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n432), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n189), .B1(new_n442), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n411), .B1(new_n439), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n416), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n432), .A2(KEYINPUT6), .B1(new_n434), .B2(new_n435), .ZN(new_n455));
  INV_X1    g269(.A(new_n438), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n432), .A2(new_n448), .A3(new_n450), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n441), .B(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(G902), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n410), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n296), .A2(new_n408), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT30), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n232), .A2(new_n226), .A3(new_n237), .A4(new_n239), .ZN(new_n471));
  INV_X1    g285(.A(new_n238), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n233), .A2(G134), .ZN(new_n473));
  OAI21_X1  g287(.A(G131), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n255), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n265), .B1(new_n240), .B2(new_n243), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n223), .A2(new_n475), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n196), .A2(new_n198), .A3(new_n260), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n196), .A2(new_n198), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n263), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n232), .A2(new_n237), .A3(new_n239), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(G131), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n483), .B1(new_n485), .B2(new_n471), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n480), .A2(new_n486), .A3(KEYINPUT30), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n423), .B1(new_n479), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT31), .ZN(new_n489));
  INV_X1    g303(.A(new_n423), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n478), .B(new_n490), .C1(new_n223), .C2(new_n475), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n312), .A2(G210), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT27), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G101), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n488), .A2(new_n489), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n495), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n423), .B1(new_n480), .B2(new_n486), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n491), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n491), .A2(new_n500), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT30), .B1(new_n480), .B2(new_n486), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n478), .B(new_n470), .C1(new_n223), .C2(new_n475), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n490), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT31), .B1(new_n507), .B2(new_n496), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n498), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT68), .ZN(new_n510));
  NOR2_X1   g324(.A1(G472), .A2(G902), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n498), .A2(new_n504), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT32), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n510), .A2(new_n516), .A3(new_n511), .A4(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n501), .A2(new_n491), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(KEYINPUT28), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n491), .A2(new_n500), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n495), .A3(new_n521), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n480), .A2(new_n486), .A3(new_n423), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n499), .B1(new_n507), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT29), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT69), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n522), .A2(new_n524), .A3(new_n528), .A4(new_n525), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n502), .A2(new_n503), .A3(new_n499), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n530), .B2(KEYINPUT29), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G472), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n518), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT70), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n518), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n307), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n319), .A2(new_n322), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G119), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n542), .A2(KEYINPUT72), .A3(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n356), .A2(G119), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT72), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT73), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n542), .B2(G128), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n356), .A2(KEYINPUT73), .A3(G119), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n543), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT23), .B1(new_n356), .B2(G119), .ZN(new_n553));
  AND2_X1   g367(.A1(KEYINPUT23), .A2(G119), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n553), .A2(new_n544), .B1(new_n356), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n541), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT76), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n541), .B(new_n562), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n331), .A2(new_n307), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n549), .A2(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  INV_X1    g384(.A(G234), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n187), .A2(new_n571), .A3(G953), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n570), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n564), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n189), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n564), .B2(new_n568), .ZN(new_n580));
  AOI211_X1 g394(.A(new_n567), .B(new_n573), .C1(new_n561), .C2(new_n563), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(KEYINPUT25), .A3(new_n189), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n387), .B1(new_n571), .B2(G902), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G902), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n584), .A2(new_n586), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT77), .B1(new_n538), .B2(new_n588), .ZN(new_n589));
  AOI221_X4 g403(.A(KEYINPUT70), .B1(new_n532), .B2(G472), .C1(new_n515), .C2(new_n517), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n536), .B1(new_n518), .B2(new_n533), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT77), .B(new_n588), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n469), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  NAND3_X1  g409(.A1(new_n510), .A2(new_n189), .A3(new_n513), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n296), .A2(new_n514), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n407), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n410), .B1(new_n439), .B2(new_n452), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n467), .B1(new_n601), .B2(new_n463), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n588), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT33), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n394), .A2(new_n604), .A3(new_n395), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT93), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n391), .A2(KEYINPUT94), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n393), .ZN(new_n608));
  INV_X1    g422(.A(new_n393), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT94), .A3(new_n391), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n608), .A2(new_n610), .A3(KEYINPUT33), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n394), .A2(new_n612), .A3(new_n604), .A4(new_n395), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n397), .A2(G902), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n606), .A2(new_n611), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n396), .A2(new_n397), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n353), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n603), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n599), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  NAND2_X1  g436(.A1(new_n402), .A2(new_n353), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n588), .A2(new_n600), .A3(new_n602), .A4(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n598), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT95), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NAND2_X1  g443(.A1(new_n296), .A2(new_n468), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT25), .B1(new_n582), .B2(new_n189), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n580), .A2(new_n581), .A3(new_n578), .A4(G902), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n586), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n564), .B2(new_n568), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n564), .A2(new_n634), .A3(new_n568), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n636), .B2(new_n638), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n587), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n633), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n642), .A2(new_n514), .A3(new_n597), .A4(new_n408), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n630), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT97), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT37), .B(G110), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n404), .B1(new_n405), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n623), .A2(new_n649), .ZN(new_n650));
  AND4_X1   g464(.A1(new_n296), .A2(new_n602), .A3(new_n642), .A4(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n590), .B2(new_n591), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XOR2_X1   g467(.A(new_n649), .B(KEYINPUT39), .Z(new_n654));
  NAND2_X1  g468(.A1(new_n296), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  INV_X1    g470(.A(new_n642), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n464), .B(KEYINPUT38), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n343), .A2(new_n349), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n352), .A2(G475), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n399), .A2(new_n401), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND4_X1   g475(.A1(new_n466), .A2(new_n657), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n507), .A2(new_n523), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n499), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n189), .B1(new_n519), .B2(new_n495), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n518), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n656), .A2(new_n662), .A3(new_n663), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  AND3_X1   g484(.A1(new_n296), .A2(new_n602), .A3(new_n642), .ZN(new_n671));
  INV_X1    g485(.A(new_n649), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n617), .A2(new_n672), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n671), .B(new_n673), .C1(new_n590), .C2(new_n591), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  OAI21_X1  g489(.A(new_n189), .B1(new_n285), .B2(new_n289), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n191), .A2(KEYINPUT98), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n251), .A2(new_n278), .A3(new_n277), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT82), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n284), .A3(new_n279), .ZN(new_n682));
  INV_X1    g496(.A(new_n677), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n189), .A3(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n190), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n678), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n619), .B(new_n687), .C1(new_n590), .C2(new_n591), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT99), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT99), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT41), .B(G113), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G15));
  NOR2_X1   g507(.A1(new_n625), .A2(new_n686), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n538), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NAND4_X1  g510(.A1(new_n678), .A2(new_n684), .A3(new_n685), .A4(new_n602), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n642), .A2(new_n408), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n538), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G119), .ZN(G21));
  AND3_X1   g515(.A1(new_n602), .A2(new_n661), .A3(new_n600), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(new_n685), .A3(new_n678), .A4(new_n684), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT100), .B(G472), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n596), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n509), .A2(new_n511), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n588), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n360), .ZN(G24));
  NAND4_X1  g523(.A1(new_n673), .A2(new_n642), .A3(new_n706), .A4(new_n705), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n697), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n320), .ZN(G27));
  NAND2_X1  g526(.A1(new_n518), .A2(KEYINPUT102), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n515), .A2(new_n714), .A3(new_n517), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n713), .A2(new_n533), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n615), .A2(new_n616), .ZN(new_n717));
  AND4_X1   g531(.A1(KEYINPUT42), .A2(new_n717), .A3(new_n354), .A4(new_n672), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n292), .A2(new_n283), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT101), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n293), .A2(new_n281), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n292), .A2(KEYINPUT101), .A3(new_n283), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n721), .A2(G469), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(new_n291), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n290), .A3(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n464), .A2(new_n467), .A3(new_n190), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n718), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n716), .A2(new_n588), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT103), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n716), .A2(new_n728), .A3(KEYINPUT103), .A4(new_n588), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n726), .A2(new_n727), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n588), .B(new_n735), .C1(new_n590), .C2(new_n591), .ZN(new_n736));
  INV_X1    g550(.A(new_n673), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  INV_X1    g554(.A(new_n650), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n228), .ZN(G36));
  NAND2_X1  g557(.A1(new_n465), .A2(new_n466), .ZN(new_n744));
  XOR2_X1   g558(.A(new_n744), .B(KEYINPUT106), .Z(new_n745));
  AOI21_X1  g559(.A(new_n657), .B1(new_n514), .B2(new_n597), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n354), .B1(new_n615), .B2(new_n616), .ZN(new_n748));
  NOR2_X1   g562(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n749));
  AND2_X1   g563(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n748), .B2(new_n750), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n746), .A2(new_n747), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n747), .B1(new_n746), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n745), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(KEYINPUT107), .B(new_n745), .C1(new_n753), .C2(new_n754), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n294), .A2(KEYINPUT45), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n191), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n721), .A2(KEYINPUT45), .A3(new_n722), .A4(new_n723), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n291), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT46), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n290), .B1(new_n763), .B2(KEYINPUT46), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n685), .B(new_n654), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n759), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G137), .ZN(G39));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n685), .B(new_n774), .C1(new_n765), .C2(new_n766), .ZN(new_n775));
  INV_X1    g589(.A(new_n290), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n761), .A2(new_n762), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n725), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT46), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n190), .B1(new_n780), .B2(new_n764), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n775), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n737), .A2(new_n588), .A3(new_n744), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n535), .A2(new_n537), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n304), .ZN(G42));
  AND2_X1   g601(.A1(new_n678), .A2(new_n684), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT49), .ZN(new_n789));
  INV_X1    g603(.A(new_n668), .ZN(new_n790));
  INV_X1    g604(.A(new_n658), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n190), .A2(new_n467), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n588), .A2(new_n791), .A3(new_n792), .A4(new_n748), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n752), .A2(new_n404), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n752), .A2(KEYINPUT111), .A3(new_n404), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n707), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n602), .A3(new_n687), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n686), .A2(new_n744), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n790), .A2(new_n801), .A3(new_n588), .A4(new_n404), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n618), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n403), .A3(G953), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n686), .B(new_n744), .C1(new_n797), .C2(new_n798), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT48), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n716), .A2(new_n588), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n805), .B2(new_n807), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n800), .B(new_n804), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n687), .A2(new_n467), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(KEYINPUT113), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n658), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT114), .B1(new_n814), .B2(new_n799), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT50), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n642), .A2(new_n706), .A3(new_n705), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n805), .A2(new_n817), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n802), .A2(new_n354), .A3(new_n717), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n816), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n815), .A2(KEYINPUT50), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n799), .A2(new_n745), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n788), .A2(new_n190), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n783), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n810), .B1(new_n822), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT115), .B1(new_n820), .B2(new_n821), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n783), .A2(KEYINPUT112), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n190), .B2(new_n788), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n783), .A2(KEYINPUT112), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n825), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n694), .A2(new_n699), .B1(new_n590), .B2(new_n591), .ZN(new_n838));
  OAI22_X1  g652(.A1(new_n630), .A2(new_n643), .B1(new_n703), .B2(new_n707), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n588), .A2(new_n468), .A3(new_n600), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n599), .B(new_n841), .C1(new_n617), .C2(new_n624), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n689), .B2(new_n690), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n594), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n735), .A2(new_n817), .A3(new_n673), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n353), .A2(new_n672), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(new_n402), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n850), .B2(new_n744), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n849), .A2(new_n402), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT109), .A3(new_n466), .A4(new_n465), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n296), .A2(new_n642), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n854), .B(new_n855), .C1(new_n590), .C2(new_n591), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n847), .B(new_n856), .C1(new_n736), .C2(new_n741), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n733), .B2(new_n738), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n710), .A2(new_n697), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n642), .A2(new_n190), .A3(new_n649), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n602), .A2(new_n661), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n668), .A2(new_n860), .A3(new_n862), .A4(new_n726), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n674), .A2(new_n652), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n711), .B1(new_n538), .B2(new_n651), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(KEYINPUT52), .A3(new_n674), .A4(new_n863), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n858), .A4(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n866), .A2(new_n868), .A3(KEYINPUT110), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n864), .A2(KEYINPUT110), .A3(new_n865), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n858), .A2(new_n844), .A3(new_n594), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT54), .ZN(new_n878));
  AND4_X1   g692(.A1(KEYINPUT53), .A2(new_n858), .A3(new_n594), .A4(new_n844), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n872), .A2(new_n873), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n869), .A2(new_n858), .A3(new_n594), .A4(new_n844), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n871), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n878), .B1(new_n884), .B2(KEYINPUT54), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n837), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n794), .B1(new_n886), .B2(new_n887), .ZN(G75));
  NOR2_X1   g702(.A1(new_n272), .A2(G952), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n189), .B1(new_n881), .B2(new_n883), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n891), .B2(new_n410), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n439), .ZN(new_n894));
  XOR2_X1   g708(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n895));
  XNOR2_X1  g709(.A(new_n894), .B(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n890), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n879), .A2(new_n880), .B1(new_n882), .B2(new_n871), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT117), .B1(new_n900), .B2(new_n189), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n882), .A2(new_n871), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n858), .A2(new_n844), .A3(KEYINPUT53), .A4(new_n594), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(new_n874), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n902), .B(G902), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n411), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n899), .B1(new_n907), .B2(KEYINPUT118), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n901), .A2(new_n906), .A3(new_n909), .A4(new_n411), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n897), .B1(new_n908), .B2(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n291), .B(KEYINPUT57), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT54), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n900), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n682), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n901), .A2(new_n762), .A3(new_n906), .A4(new_n761), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n889), .B1(new_n917), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n901), .A2(new_n906), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n340), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n901), .A2(new_n906), .A3(new_n347), .A4(new_n920), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n890), .A3(new_n923), .ZN(G60));
  AND3_X1   g738(.A1(new_n606), .A2(new_n613), .A3(new_n611), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT59), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n927), .C1(new_n913), .C2(new_n915), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n890), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n925), .B1(new_n885), .B2(new_n927), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT119), .Z(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n639), .A2(new_n640), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT120), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n934), .B(new_n936), .C1(new_n903), .C2(new_n905), .ZN(new_n937));
  INV_X1    g751(.A(new_n934), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n900), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n890), .B(new_n937), .C1(new_n939), .C2(new_n582), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G66));
  OAI21_X1  g756(.A(G953), .B1(new_n406), .B2(new_n414), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n846), .B2(G953), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n437), .B(new_n438), .C1(G898), .C2(new_n272), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT121), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n944), .B(new_n946), .ZN(G69));
  AOI21_X1  g761(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n479), .A2(new_n487), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT122), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n300), .A2(new_n301), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(new_n952));
  AOI211_X1 g766(.A(new_n744), .B(new_n655), .C1(new_n618), .C2(new_n623), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n589), .B2(new_n593), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n786), .B1(new_n759), .B2(new_n769), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n674), .A2(new_n652), .A3(new_n859), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n669), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT123), .B1(new_n960), .B2(KEYINPUT62), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT62), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n959), .A2(new_n964), .A3(new_n965), .A4(new_n669), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT125), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  AOI22_X1  g783(.A1(new_n955), .A2(new_n956), .B1(KEYINPUT62), .B2(new_n960), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n970), .A2(new_n967), .A3(new_n971), .A4(new_n958), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n952), .B1(new_n973), .B2(new_n272), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n769), .A2(new_n862), .A3(new_n807), .ZN(new_n975));
  INV_X1    g789(.A(new_n959), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n976), .A2(new_n742), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n739), .A2(new_n958), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n272), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n952), .B1(new_n648), .B2(new_n272), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n948), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n948), .ZN(new_n983));
  AOI21_X1  g797(.A(G953), .B1(new_n969), .B2(new_n972), .ZN(new_n984));
  OAI221_X1 g798(.A(new_n983), .B1(new_n979), .B2(new_n980), .C1(new_n984), .C2(new_n952), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n985), .ZN(G72));
  XNOR2_X1  g800(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n524), .B1(new_n507), .B2(new_n496), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n877), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n989), .B(KEYINPUT127), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n978), .B2(new_n846), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n664), .A2(new_n499), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n991), .B(new_n890), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n992), .B1(new_n973), .B2(new_n845), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n665), .B2(new_n997), .ZN(G57));
endmodule


