

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  XOR2_X1 U321 ( .A(n383), .B(n382), .Z(n558) );
  XNOR2_X1 U322 ( .A(KEYINPUT48), .B(KEYINPUT109), .ZN(n380) );
  XNOR2_X1 U323 ( .A(n545), .B(n372), .ZN(n578) );
  XNOR2_X1 U324 ( .A(n343), .B(n342), .ZN(n346) );
  AND2_X1 U325 ( .A1(G232GAT), .A2(G233GAT), .ZN(n289) );
  XNOR2_X1 U326 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n373) );
  XNOR2_X1 U327 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U328 ( .A(KEYINPUT116), .B(KEYINPUT54), .ZN(n382) );
  XNOR2_X1 U329 ( .A(n341), .B(KEYINPUT31), .ZN(n342) );
  XNOR2_X1 U330 ( .A(n296), .B(n289), .ZN(n297) );
  XNOR2_X1 U331 ( .A(n371), .B(KEYINPUT94), .ZN(n372) );
  XNOR2_X1 U332 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U333 ( .A(n445), .B(KEYINPUT118), .Z(n556) );
  XNOR2_X1 U334 ( .A(n446), .B(G190GAT), .ZN(n447) );
  XOR2_X1 U335 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n291) );
  XNOR2_X1 U336 ( .A(KEYINPUT72), .B(KEYINPUT11), .ZN(n290) );
  XNOR2_X1 U337 ( .A(n291), .B(n290), .ZN(n300) );
  XOR2_X1 U338 ( .A(G99GAT), .B(G85GAT), .Z(n340) );
  XOR2_X1 U339 ( .A(n340), .B(G92GAT), .Z(n293) );
  XOR2_X1 U340 ( .A(G162GAT), .B(G106GAT), .Z(n419) );
  XNOR2_X1 U341 ( .A(G218GAT), .B(n419), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n298) );
  XOR2_X1 U343 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n295) );
  XNOR2_X1 U344 ( .A(G134GAT), .B(G190GAT), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n306) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n301), .B(G29GAT), .ZN(n302) );
  XOR2_X1 U349 ( .A(n302), .B(KEYINPUT8), .Z(n304) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G50GAT), .ZN(n303) );
  XOR2_X1 U351 ( .A(n304), .B(n303), .Z(n361) );
  INV_X1 U352 ( .A(n361), .ZN(n305) );
  XOR2_X1 U353 ( .A(n306), .B(n305), .Z(n545) );
  INV_X1 U354 ( .A(n545), .ZN(n530) );
  XOR2_X1 U355 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n308) );
  XNOR2_X1 U356 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U358 ( .A(G190GAT), .B(KEYINPUT17), .Z(n309) );
  XOR2_X1 U359 ( .A(n310), .B(n309), .Z(n441) );
  XOR2_X1 U360 ( .A(G169GAT), .B(G8GAT), .Z(n351) );
  XOR2_X1 U361 ( .A(n351), .B(KEYINPUT91), .Z(n312) );
  NAND2_X1 U362 ( .A1(G226GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U364 ( .A(G92GAT), .B(G64GAT), .Z(n314) );
  XNOR2_X1 U365 ( .A(G176GAT), .B(KEYINPUT71), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U367 ( .A(G204GAT), .B(n315), .Z(n348) );
  XOR2_X1 U368 ( .A(n316), .B(n348), .Z(n322) );
  XNOR2_X1 U369 ( .A(G211GAT), .B(KEYINPUT80), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n317), .B(KEYINPUT21), .ZN(n318) );
  XOR2_X1 U371 ( .A(n318), .B(KEYINPUT79), .Z(n320) );
  XNOR2_X1 U372 ( .A(G197GAT), .B(G218GAT), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n320), .B(n319), .ZN(n423) );
  XNOR2_X1 U374 ( .A(G36GAT), .B(n423), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(n441), .B(n323), .Z(n494) );
  INV_X1 U377 ( .A(n494), .ZN(n509) );
  XNOR2_X1 U378 ( .A(G15GAT), .B(G22GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n324), .B(G1GAT), .ZN(n350) );
  XOR2_X1 U380 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n326) );
  XNOR2_X1 U381 ( .A(G8GAT), .B(G64GAT), .ZN(n325) );
  XNOR2_X1 U382 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U383 ( .A(n350), .B(n327), .ZN(n336) );
  XOR2_X1 U384 ( .A(KEYINPUT13), .B(G57GAT), .Z(n329) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(G78GAT), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n344) );
  XOR2_X1 U387 ( .A(n344), .B(KEYINPUT15), .Z(n331) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(G127GAT), .B(G155GAT), .Z(n387) );
  XOR2_X1 U391 ( .A(n332), .B(n387), .Z(n334) );
  XNOR2_X1 U392 ( .A(G183GAT), .B(G211GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U394 ( .A(n336), .B(n335), .ZN(n473) );
  INV_X1 U395 ( .A(n473), .ZN(n571) );
  XOR2_X1 U396 ( .A(KEYINPUT104), .B(n571), .Z(n555) );
  XNOR2_X1 U397 ( .A(KEYINPUT105), .B(KEYINPUT46), .ZN(n365) );
  INV_X1 U398 ( .A(KEYINPUT41), .ZN(n349) );
  XOR2_X1 U399 ( .A(KEYINPUT33), .B(G106GAT), .Z(n338) );
  XNOR2_X1 U400 ( .A(G120GAT), .B(G148GAT), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U402 ( .A(n340), .B(n339), .Z(n343) );
  NAND2_X1 U403 ( .A1(G230GAT), .A2(G233GAT), .ZN(n341) );
  XOR2_X1 U404 ( .A(n344), .B(KEYINPUT32), .Z(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X2 U406 ( .A(n348), .B(n347), .Z(n566) );
  XNOR2_X1 U407 ( .A(n349), .B(n566), .ZN(n488) );
  XOR2_X1 U408 ( .A(n351), .B(n350), .Z(n353) );
  NAND2_X1 U409 ( .A1(G229GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U411 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n355) );
  XNOR2_X1 U412 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U414 ( .A(n357), .B(n356), .Z(n363) );
  XOR2_X1 U415 ( .A(KEYINPUT68), .B(G197GAT), .Z(n359) );
  XNOR2_X1 U416 ( .A(G113GAT), .B(G141GAT), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U418 ( .A(n361), .B(n360), .Z(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n562) );
  NOR2_X1 U420 ( .A1(n488), .A2(n562), .ZN(n364) );
  XOR2_X1 U421 ( .A(n365), .B(n364), .Z(n366) );
  NOR2_X1 U422 ( .A1(n555), .A2(n366), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n367), .B(KEYINPUT106), .ZN(n368) );
  NAND2_X1 U424 ( .A1(n368), .A2(n545), .ZN(n369) );
  XNOR2_X1 U425 ( .A(n369), .B(KEYINPUT47), .ZN(n370) );
  XOR2_X1 U426 ( .A(KEYINPUT107), .B(n370), .Z(n379) );
  XOR2_X1 U427 ( .A(n562), .B(KEYINPUT70), .Z(n547) );
  INV_X1 U428 ( .A(KEYINPUT36), .ZN(n371) );
  NAND2_X1 U429 ( .A1(n578), .A2(n473), .ZN(n374) );
  NAND2_X1 U430 ( .A1(n375), .A2(n566), .ZN(n376) );
  NOR2_X1 U431 ( .A1(n547), .A2(n376), .ZN(n377) );
  XNOR2_X1 U432 ( .A(KEYINPUT108), .B(n377), .ZN(n378) );
  NOR2_X1 U433 ( .A1(n379), .A2(n378), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n381), .B(n380), .ZN(n516) );
  NAND2_X1 U435 ( .A1(n509), .A2(n516), .ZN(n383) );
  XOR2_X1 U436 ( .A(KEYINPUT90), .B(G85GAT), .Z(n385) );
  XNOR2_X1 U437 ( .A(G29GAT), .B(G162GAT), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U439 ( .A(n387), .B(n386), .Z(n389) );
  NAND2_X1 U440 ( .A1(G225GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n405) );
  XOR2_X1 U442 ( .A(KEYINPUT86), .B(G57GAT), .Z(n391) );
  XNOR2_X1 U443 ( .A(G1GAT), .B(KEYINPUT87), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U445 ( .A(KEYINPUT84), .B(KEYINPUT1), .Z(n393) );
  XNOR2_X1 U446 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U448 ( .A(n395), .B(n394), .Z(n403) );
  XOR2_X1 U449 ( .A(KEYINPUT0), .B(G134GAT), .Z(n397) );
  XNOR2_X1 U450 ( .A(KEYINPUT74), .B(G120GAT), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U452 ( .A(G113GAT), .B(n398), .Z(n443) );
  XOR2_X1 U453 ( .A(KEYINPUT4), .B(KEYINPUT85), .Z(n400) );
  XNOR2_X1 U454 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n443), .B(n401), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U459 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n407) );
  XNOR2_X1 U460 ( .A(KEYINPUT81), .B(G148GAT), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U462 ( .A(G141GAT), .B(n408), .ZN(n427) );
  XOR2_X1 U463 ( .A(n409), .B(n427), .Z(n559) );
  XOR2_X1 U464 ( .A(G204GAT), .B(KEYINPUT83), .Z(n411) );
  XNOR2_X1 U465 ( .A(G22GAT), .B(KEYINPUT77), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U467 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n413) );
  XNOR2_X1 U468 ( .A(G155GAT), .B(G78GAT), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U470 ( .A(n415), .B(n414), .Z(n425) );
  XOR2_X1 U471 ( .A(KEYINPUT78), .B(KEYINPUT22), .Z(n417) );
  XNOR2_X1 U472 ( .A(G50GAT), .B(KEYINPUT82), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U474 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U479 ( .A(n427), .B(n426), .Z(n455) );
  AND2_X1 U480 ( .A1(n559), .A2(n455), .ZN(n428) );
  NAND2_X1 U481 ( .A1(n558), .A2(n428), .ZN(n430) );
  XOR2_X1 U482 ( .A(KEYINPUT117), .B(KEYINPUT55), .Z(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n444) );
  XOR2_X1 U484 ( .A(G176GAT), .B(KEYINPUT20), .Z(n432) );
  XNOR2_X1 U485 ( .A(G169GAT), .B(KEYINPUT75), .ZN(n431) );
  XNOR2_X1 U486 ( .A(n432), .B(n431), .ZN(n439) );
  XOR2_X1 U487 ( .A(G71GAT), .B(G99GAT), .Z(n434) );
  XNOR2_X1 U488 ( .A(G43GAT), .B(G15GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(G127GAT), .B(n435), .Z(n437) );
  NAND2_X1 U491 ( .A1(G227GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U493 ( .A(n439), .B(n438), .Z(n440) );
  XOR2_X1 U494 ( .A(n441), .B(n440), .Z(n442) );
  XOR2_X1 U495 ( .A(n443), .B(n442), .Z(n496) );
  INV_X1 U496 ( .A(n496), .ZN(n517) );
  NAND2_X1 U497 ( .A1(n444), .A2(n517), .ZN(n445) );
  NAND2_X1 U498 ( .A1(n530), .A2(n556), .ZN(n448) );
  XOR2_X1 U499 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n446) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(G1351GAT) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n464) );
  NAND2_X1 U502 ( .A1(n547), .A2(n566), .ZN(n476) );
  NOR2_X1 U503 ( .A1(n530), .A2(n571), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n449), .B(KEYINPUT16), .ZN(n462) );
  XOR2_X1 U505 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n450) );
  XOR2_X1 U506 ( .A(n455), .B(n450), .Z(n499) );
  XOR2_X1 U507 ( .A(KEYINPUT27), .B(n494), .Z(n457) );
  AND2_X1 U508 ( .A1(n499), .A2(n457), .ZN(n451) );
  INV_X1 U509 ( .A(n559), .ZN(n507) );
  NAND2_X1 U510 ( .A1(n451), .A2(n507), .ZN(n518) );
  XOR2_X1 U511 ( .A(KEYINPUT92), .B(n518), .Z(n452) );
  NAND2_X1 U512 ( .A1(n496), .A2(n452), .ZN(n461) );
  NAND2_X1 U513 ( .A1(n517), .A2(n509), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n455), .A2(n453), .ZN(n454) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n454), .Z(n458) );
  NOR2_X1 U516 ( .A1(n455), .A2(n517), .ZN(n456) );
  XNOR2_X1 U517 ( .A(n456), .B(KEYINPUT26), .ZN(n561) );
  NAND2_X1 U518 ( .A1(n457), .A2(n561), .ZN(n534) );
  NAND2_X1 U519 ( .A1(n458), .A2(n534), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n559), .A2(n459), .ZN(n460) );
  NAND2_X1 U521 ( .A1(n461), .A2(n460), .ZN(n471) );
  NAND2_X1 U522 ( .A1(n462), .A2(n471), .ZN(n489) );
  NOR2_X1 U523 ( .A1(n476), .A2(n489), .ZN(n469) );
  NAND2_X1 U524 ( .A1(n469), .A2(n507), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n464), .B(n463), .ZN(G1324GAT) );
  XOR2_X1 U526 ( .A(G8GAT), .B(KEYINPUT93), .Z(n466) );
  NAND2_X1 U527 ( .A1(n469), .A2(n509), .ZN(n465) );
  XNOR2_X1 U528 ( .A(n466), .B(n465), .ZN(G1325GAT) );
  XOR2_X1 U529 ( .A(G15GAT), .B(KEYINPUT35), .Z(n468) );
  NAND2_X1 U530 ( .A1(n469), .A2(n517), .ZN(n467) );
  XNOR2_X1 U531 ( .A(n468), .B(n467), .ZN(G1326GAT) );
  INV_X1 U532 ( .A(n499), .ZN(n512) );
  NAND2_X1 U533 ( .A1(n469), .A2(n512), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n470), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U535 ( .A1(n578), .A2(n471), .ZN(n472) );
  NOR2_X1 U536 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U537 ( .A(KEYINPUT37), .B(n474), .Z(n475) );
  XNOR2_X1 U538 ( .A(KEYINPUT95), .B(n475), .ZN(n506) );
  NOR2_X1 U539 ( .A1(n506), .A2(n476), .ZN(n477) );
  XOR2_X1 U540 ( .A(KEYINPUT38), .B(n477), .Z(n486) );
  NOR2_X1 U541 ( .A1(n486), .A2(n559), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n478), .B(KEYINPUT39), .ZN(n479) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(n479), .ZN(G1328GAT) );
  NOR2_X1 U544 ( .A1(n494), .A2(n486), .ZN(n480) );
  XOR2_X1 U545 ( .A(G36GAT), .B(n480), .Z(n481) );
  XNOR2_X1 U546 ( .A(KEYINPUT96), .B(n481), .ZN(G1329GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n483) );
  XNOR2_X1 U548 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n482) );
  XNOR2_X1 U549 ( .A(n483), .B(n482), .ZN(n485) );
  NOR2_X1 U550 ( .A1(n496), .A2(n486), .ZN(n484) );
  XOR2_X1 U551 ( .A(n485), .B(n484), .Z(G1330GAT) );
  NOR2_X1 U552 ( .A1(n486), .A2(n499), .ZN(n487) );
  XOR2_X1 U553 ( .A(G50GAT), .B(n487), .Z(G1331GAT) );
  BUF_X1 U554 ( .A(n488), .Z(n539) );
  INV_X1 U555 ( .A(n539), .ZN(n552) );
  NAND2_X1 U556 ( .A1(n562), .A2(n552), .ZN(n505) );
  NOR2_X1 U557 ( .A1(n489), .A2(n505), .ZN(n490) );
  XNOR2_X1 U558 ( .A(n490), .B(KEYINPUT99), .ZN(n500) );
  NOR2_X1 U559 ( .A1(n559), .A2(n500), .ZN(n492) );
  XNOR2_X1 U560 ( .A(KEYINPUT100), .B(KEYINPUT42), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U562 ( .A(G57GAT), .B(n493), .Z(G1332GAT) );
  NOR2_X1 U563 ( .A1(n494), .A2(n500), .ZN(n495) );
  XOR2_X1 U564 ( .A(G64GAT), .B(n495), .Z(G1333GAT) );
  NOR2_X1 U565 ( .A1(n496), .A2(n500), .ZN(n498) );
  XNOR2_X1 U566 ( .A(G71GAT), .B(KEYINPUT101), .ZN(n497) );
  XNOR2_X1 U567 ( .A(n498), .B(n497), .ZN(G1334GAT) );
  NOR2_X1 U568 ( .A1(n500), .A2(n499), .ZN(n504) );
  XOR2_X1 U569 ( .A(KEYINPUT102), .B(KEYINPUT43), .Z(n502) );
  XNOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT103), .ZN(n501) );
  XNOR2_X1 U571 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NOR2_X1 U573 ( .A1(n506), .A2(n505), .ZN(n513) );
  NAND2_X1 U574 ( .A1(n513), .A2(n507), .ZN(n508) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n509), .A2(n513), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n517), .A2(n513), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT44), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n515), .ZN(G1339GAT) );
  XOR2_X1 U583 ( .A(G113GAT), .B(KEYINPUT111), .Z(n522) );
  BUF_X1 U584 ( .A(n516), .Z(n536) );
  NAND2_X1 U585 ( .A1(n536), .A2(n517), .ZN(n519) );
  NOR2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(KEYINPUT110), .ZN(n529) );
  NAND2_X1 U588 ( .A1(n547), .A2(n529), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n524) );
  NAND2_X1 U591 ( .A1(n529), .A2(n552), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(n526) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT112), .Z(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1341GAT) );
  NAND2_X1 U595 ( .A1(n529), .A2(n555), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n527), .B(KEYINPUT50), .ZN(n528) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n532) );
  NAND2_X1 U599 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n533), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n559), .A2(n534), .ZN(n535) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n544) );
  NOR2_X1 U604 ( .A1(n562), .A2(n544), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1344GAT) );
  NOR2_X1 U607 ( .A1(n539), .A2(n544), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n542), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n571), .A2(n544), .ZN(n543) );
  XOR2_X1 U612 ( .A(G155GAT), .B(n543), .Z(G1346GAT) );
  NOR2_X1 U613 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U614 ( .A(G162GAT), .B(n546), .Z(G1347GAT) );
  NAND2_X1 U615 ( .A1(n556), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n550) );
  XNOR2_X1 U618 ( .A(G176GAT), .B(KEYINPUT119), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(n551), .Z(n554) );
  NAND2_X1 U621 ( .A1(n556), .A2(n552), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n576) );
  XNOR2_X1 U627 ( .A(n576), .B(KEYINPUT122), .ZN(n572) );
  NOR2_X1 U628 ( .A1(n572), .A2(n562), .ZN(n565) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1352GAT) );
  NOR2_X1 U632 ( .A1(n572), .A2(n566), .ZN(n570) );
  XOR2_X1 U633 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U634 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n580) );
  XOR2_X1 U642 ( .A(n576), .B(KEYINPUT122), .Z(n577) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

