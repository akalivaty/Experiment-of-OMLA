//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NAND2_X1  g003(.A1(G125), .A2(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  OR3_X1    g006(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n194), .B(G146), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT66), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G128), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT69), .B(G119), .ZN(new_n201));
  AOI22_X1  g015(.A1(G119), .A2(new_n200), .B1(new_n201), .B2(G128), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT24), .B(G110), .Z(new_n203));
  AOI21_X1  g017(.A(new_n195), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G110), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n206));
  OR3_X1    g020(.A1(new_n201), .A2(KEYINPUT23), .A3(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n204), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n191), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(G110), .B1(new_n206), .B2(new_n207), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n202), .A2(new_n203), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n192), .A2(G146), .A3(new_n193), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT75), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n215), .B(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT22), .ZN(new_n221));
  INV_X1    g035(.A(G137), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n223), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT25), .B1(new_n226), .B2(G902), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(G234), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n224), .A2(new_n231), .A3(new_n229), .A4(new_n225), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT77), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(G902), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(KEYINPUT76), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n224), .A2(new_n236), .A3(new_n225), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n233), .B2(new_n237), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n210), .A2(G143), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(G143), .B2(new_n210), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n200), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G143), .B(G146), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n245), .A3(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(G134), .A2(G137), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT64), .B(G137), .ZN(new_n252));
  OAI211_X1 g066(.A(G131), .B(new_n251), .C1(new_n252), .C2(G134), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT11), .A2(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT11), .A2(G134), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(G137), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n256), .B(new_n257), .C1(new_n252), .C2(new_n255), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n250), .A2(new_n253), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT70), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT2), .A2(G113), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(KEYINPUT2), .A2(G113), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n201), .A2(G116), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G119), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n263), .A2(new_n264), .B1(new_n266), .B2(new_n268), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n250), .A2(new_n273), .A3(new_n253), .A4(new_n258), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT0), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(new_n196), .ZN(new_n276));
  NOR2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n244), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n248), .B1(new_n275), .B2(new_n196), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT64), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G137), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n255), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n257), .B1(new_n286), .B2(new_n256), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n255), .B1(new_n281), .B2(new_n283), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n255), .A2(G137), .ZN(new_n289));
  OR2_X1    g103(.A1(KEYINPUT11), .A2(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n288), .A2(new_n291), .A3(G131), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n280), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n260), .A2(new_n272), .A3(new_n274), .A4(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n288), .B2(new_n291), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n258), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n259), .A2(KEYINPUT70), .B1(new_n298), .B2(new_n280), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(KEYINPUT72), .A3(new_n272), .A4(new_n274), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(G101), .ZN(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n310));
  INV_X1    g124(.A(new_n259), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n293), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n298), .A2(KEYINPUT65), .A3(new_n280), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n310), .B1(new_n315), .B2(KEYINPUT30), .ZN(new_n316));
  OR2_X1    g130(.A1(new_n270), .A2(new_n271), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n299), .A2(KEYINPUT30), .A3(new_n274), .ZN(new_n318));
  AOI221_X4 g132(.A(new_n312), .B1(new_n278), .B2(new_n279), .C1(new_n258), .C2(new_n297), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT65), .B1(new_n298), .B2(new_n280), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n259), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(KEYINPUT67), .A3(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n316), .A2(new_n317), .A3(new_n318), .A4(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n324), .A2(new_n325), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n309), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT31), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n315), .A2(new_n272), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n302), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n272), .A2(new_n259), .A3(new_n293), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n308), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n337), .B(new_n309), .C1(new_n326), .C2(new_n327), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n329), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(G472), .A2(G902), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(KEYINPUT32), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n339), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G472), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n339), .A2(new_n346), .A3(new_n229), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT32), .ZN(new_n348));
  INV_X1    g162(.A(new_n334), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n299), .A2(new_n274), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n317), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n301), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n349), .B1(new_n352), .B2(KEYINPUT28), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT29), .A4(new_n307), .ZN(new_n355));
  AOI22_X1  g169(.A1(new_n296), .A2(new_n300), .B1(new_n350), .B2(new_n317), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT29), .B(new_n334), .C1(new_n356), .C2(new_n333), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT73), .B1(new_n357), .B2(new_n308), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n308), .B1(new_n331), .B2(new_n334), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n316), .A2(new_n323), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(KEYINPUT71), .A3(new_n317), .A4(new_n318), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n324), .A2(new_n325), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n302), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n360), .B1(new_n364), .B2(new_n308), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n229), .B(new_n359), .C1(new_n365), .C2(KEYINPUT29), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n347), .A2(new_n348), .B1(new_n366), .B2(G472), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n240), .B1(new_n345), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT9), .B(G234), .Z(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G221), .B1(new_n371), .B2(G902), .ZN(new_n372));
  INV_X1    g186(.A(G469), .ZN(new_n373));
  INV_X1    g187(.A(G107), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G104), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT78), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT78), .A2(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n375), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  OAI211_X1 g195(.A(G104), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G107), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n380), .A2(new_n381), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n375), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT79), .B1(new_n383), .B2(G107), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g203(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n244), .B1(new_n246), .B2(new_n196), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n249), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n380), .A2(new_n382), .A3(new_n384), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G101), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n396), .A2(new_n399), .A3(G101), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n280), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(KEYINPUT10), .A3(new_n250), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(new_n298), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n385), .A2(new_n389), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n247), .A3(new_n249), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n393), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI211_X1 g224(.A(KEYINPUT80), .B(KEYINPUT12), .C1(new_n393), .C2(new_n407), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n298), .B(new_n410), .C1(new_n411), .C2(new_n409), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT80), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n408), .A2(new_n413), .A3(new_n298), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT12), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n405), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G140), .ZN(new_n417));
  INV_X1    g231(.A(G227), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G953), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n417), .B(new_n419), .Z(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n404), .A2(new_n421), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n403), .A2(new_n298), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT82), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n425), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n373), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n423), .A2(new_n415), .A3(new_n412), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n420), .B1(new_n405), .B2(new_n424), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n373), .B(new_n229), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(G469), .A2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n372), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n317), .A2(new_n398), .A3(new_n400), .ZN(new_n439));
  INV_X1    g253(.A(new_n270), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n266), .A2(KEYINPUT5), .A3(new_n268), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n441), .B(G113), .C1(KEYINPUT5), .C2(new_n266), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n390), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(G110), .B(G122), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n439), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(KEYINPUT6), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n278), .A2(new_n279), .A3(G125), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n250), .B2(G125), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(KEYINPUT83), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G224), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(G953), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n455), .B(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n444), .A2(new_n459), .A3(new_n445), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n449), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n440), .A2(new_n442), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n406), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n443), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n445), .B(KEYINPUT8), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n451), .B1(new_n468), .B2(new_n457), .ZN(new_n469));
  INV_X1    g283(.A(new_n457), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n453), .A2(KEYINPUT7), .A3(new_n470), .A4(new_n454), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n467), .A2(new_n469), .A3(new_n448), .A4(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n461), .A2(new_n229), .A3(new_n462), .A4(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT87), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n461), .A2(new_n229), .A3(new_n472), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n461), .A2(KEYINPUT84), .A3(new_n229), .A4(new_n472), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n462), .B(KEYINPUT85), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n475), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AOI211_X1 g297(.A(KEYINPUT86), .B(new_n481), .C1(new_n478), .C2(new_n479), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n474), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(G234), .A2(G237), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(G952), .A3(new_n219), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT21), .B(G898), .Z(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(G902), .A3(G953), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(G214), .B1(G237), .B2(G902), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(G475), .A2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n305), .A2(G214), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n242), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n305), .A2(G143), .A3(G214), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT18), .A2(G131), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n189), .A2(KEYINPUT89), .A3(new_n190), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT89), .B1(new_n189), .B2(new_n190), .ZN(new_n506));
  OAI21_X1  g320(.A(G146), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n211), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n500), .A2(new_n257), .A3(new_n501), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n257), .B1(new_n500), .B2(new_n501), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT90), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n502), .A2(G131), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n500), .A2(new_n257), .A3(new_n501), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT19), .B1(new_n505), .B2(new_n506), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT19), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n191), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n512), .B(new_n516), .C1(G146), .C2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n509), .B1(new_n521), .B2(new_n217), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n523));
  XOR2_X1   g337(.A(G113), .B(G122), .Z(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT92), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(new_n383), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n509), .B(new_n527), .C1(new_n521), .C2(new_n217), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n526), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n511), .A2(KEYINPUT17), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n513), .A2(new_n515), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n195), .B(new_n531), .C1(new_n532), .C2(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n533), .A3(new_n509), .ZN(new_n534));
  AOI211_X1 g348(.A(KEYINPUT20), .B(new_n498), .C1(new_n529), .C2(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n529), .A2(new_n534), .A3(KEYINPUT93), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT93), .B1(new_n529), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n497), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XOR2_X1   g352(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n539));
  AOI21_X1  g353(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(G475), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n509), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n526), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n534), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n541), .B1(new_n544), .B2(new_n229), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n267), .A2(G122), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n267), .A2(G122), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(G107), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n552));
  INV_X1    g366(.A(new_n549), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n374), .B1(new_n553), .B2(KEYINPUT14), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n242), .A2(G128), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT66), .B(G128), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n242), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT95), .ZN(new_n559));
  INV_X1    g373(.A(G134), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n555), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n557), .A2(new_n242), .B1(new_n564), .B2(new_n556), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT13), .B1(new_n242), .B2(G128), .ZN(new_n566));
  OAI21_X1  g380(.A(G134), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT94), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n559), .A2(new_n560), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n550), .B(G107), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n371), .A2(new_n228), .A3(G953), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT96), .ZN(new_n575));
  INV_X1    g389(.A(new_n573), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n563), .A2(new_n571), .A3(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n575), .A3(new_n229), .A4(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n547), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n438), .A2(new_n485), .A3(new_n496), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n369), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n381), .ZN(G3));
  NAND2_X1  g401(.A1(new_n339), .A2(new_n229), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n346), .A2(KEYINPUT97), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n240), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n438), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n493), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n574), .A2(new_n595), .A3(new_n577), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n579), .A2(G902), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT100), .B1(new_n572), .B2(KEYINPUT99), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT100), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n599), .B1(new_n576), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n598), .A2(new_n576), .B1(new_n572), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n596), .B(new_n597), .C1(new_n602), .C2(new_n595), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n574), .A2(new_n577), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n229), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n579), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n547), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n462), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n476), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(KEYINPUT98), .A3(new_n473), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n473), .A2(KEYINPUT98), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n494), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n593), .A2(new_n594), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT101), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  XNOR2_X1  g432(.A(new_n538), .B(new_n539), .ZN(new_n619));
  INV_X1    g433(.A(new_n545), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n583), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n613), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n593), .A2(new_n594), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT102), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G107), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  INV_X1    g440(.A(new_n590), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n223), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n218), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n236), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n233), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n585), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT37), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G110), .ZN(G12));
  NAND2_X1  g449(.A1(new_n345), .A2(new_n367), .ZN(new_n636));
  INV_X1    g450(.A(new_n613), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n631), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n492), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n487), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n619), .A2(new_n620), .A3(new_n583), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n437), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n636), .A2(new_n639), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  OR2_X1    g460(.A1(new_n485), .A2(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n485), .A2(KEYINPUT103), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(KEYINPUT38), .A3(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT38), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n650), .A2(new_n495), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n642), .B(KEYINPUT39), .Z(new_n653));
  NOR2_X1   g467(.A1(new_n437), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n347), .A2(new_n348), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n364), .A2(new_n308), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n229), .B1(new_n352), .B2(new_n307), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n345), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n656), .A2(new_n662), .A3(new_n631), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n547), .A2(new_n583), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n655), .A2(KEYINPUT40), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n652), .A2(new_n663), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  OAI211_X1 g482(.A(new_n607), .B(new_n642), .C1(new_n540), .C2(new_n545), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n437), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n636), .A2(new_n639), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  NOR2_X1   g486(.A1(new_n432), .A2(new_n433), .ZN(new_n673));
  OAI21_X1  g487(.A(G469), .B1(new_n673), .B2(G902), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n674), .A2(new_n372), .A3(new_n434), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n594), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n368), .A2(new_n614), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G113), .ZN(G15));
  NAND3_X1  g494(.A1(new_n368), .A2(new_n622), .A3(new_n677), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  AOI21_X1  g496(.A(new_n638), .B1(new_n345), .B2(new_n367), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n584), .A3(new_n677), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  NOR3_X1   g499(.A1(new_n664), .A2(new_n676), .A3(new_n613), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n353), .A2(new_n307), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n329), .A2(new_n338), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n340), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n688), .A2(KEYINPUT104), .A3(new_n340), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n233), .A2(new_n237), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT105), .B(G472), .Z(new_n696));
  NAND2_X1  g510(.A1(new_n588), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n686), .A2(new_n693), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  AND4_X1   g513(.A1(new_n631), .A2(new_n691), .A3(new_n697), .A4(new_n692), .ZN(new_n700));
  INV_X1    g514(.A(new_n675), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n613), .A3(new_n669), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT106), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n187), .ZN(G27));
  INV_X1    g519(.A(new_n669), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n428), .A2(new_n373), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n372), .B1(new_n436), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n474), .B(new_n494), .C1(new_n483), .C2(new_n484), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n368), .A2(new_n706), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n366), .A2(G472), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n657), .A2(new_n714), .A3(new_n341), .ZN(new_n715));
  AND4_X1   g529(.A1(KEYINPUT42), .A2(new_n715), .A3(new_n711), .A4(new_n695), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n669), .A2(new_n708), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n712), .A2(new_n713), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n257), .ZN(G33));
  INV_X1    g533(.A(new_n643), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n368), .A2(new_n720), .A3(new_n709), .A4(new_n711), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  INV_X1    g536(.A(new_n607), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(KEYINPUT43), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n546), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n546), .B(KEYINPUT107), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n723), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n627), .A3(new_n631), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n426), .A2(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n427), .A2(new_n430), .ZN(new_n735));
  OAI211_X1 g549(.A(G469), .B(new_n734), .C1(new_n735), .C2(KEYINPUT45), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n435), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT46), .B1(new_n736), .B2(new_n435), .ZN(new_n739));
  INV_X1    g553(.A(new_n434), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n372), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n741), .A2(new_n742), .A3(new_n653), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n731), .A2(new_n732), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n733), .A2(new_n711), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT108), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G137), .ZN(G39));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n741), .B2(new_n742), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n739), .A2(new_n740), .ZN(new_n750));
  OAI211_X1 g564(.A(KEYINPUT47), .B(new_n372), .C1(new_n750), .C2(new_n738), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n636), .A2(new_n669), .A3(new_n710), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n240), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  AOI21_X1  g569(.A(new_n694), .B1(new_n367), .B2(new_n341), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n710), .A2(new_n487), .A3(new_n701), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n730), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n693), .A2(new_n697), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n695), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n729), .A3(new_n487), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n674), .A2(new_n434), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(new_n742), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n711), .B(new_n764), .C1(new_n752), .C2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n730), .A2(new_n700), .A3(new_n757), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n770));
  INV_X1    g584(.A(new_n763), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n730), .A3(new_n488), .A4(new_n675), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n495), .B1(new_n650), .B2(new_n651), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n773), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n775), .A2(new_n764), .A3(KEYINPUT50), .A4(new_n675), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n769), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n662), .A2(new_n591), .A3(new_n757), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT116), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n546), .A3(new_n723), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT51), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n774), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n781), .A3(new_n768), .A4(new_n767), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT117), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n547), .A3(new_n607), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n758), .B(new_n759), .ZN(new_n789));
  OAI211_X1 g603(.A(G952), .B(new_n219), .C1(new_n789), .C2(new_n760), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n784), .B2(new_n785), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n761), .A2(new_n787), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n678), .A2(new_n681), .A3(new_n684), .A4(new_n698), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n718), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n645), .A2(new_n671), .A3(new_n703), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n664), .A2(new_n613), .A3(new_n708), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n661), .A2(new_n632), .A3(new_n642), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n683), .A2(new_n644), .B1(new_n700), .B2(new_n702), .ZN(new_n799));
  AND4_X1   g613(.A1(KEYINPUT52), .A2(new_n799), .A3(new_n671), .A4(new_n797), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n794), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT109), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n583), .B(new_n802), .ZN(new_n803));
  MUX2_X1   g617(.A(new_n723), .B(new_n803), .S(new_n546), .Z(new_n804));
  NAND2_X1  g618(.A1(new_n485), .A2(new_n496), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n592), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n586), .A2(new_n806), .A3(new_n633), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n691), .A2(new_n717), .A3(new_n692), .A4(new_n697), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n803), .A2(new_n620), .A3(new_n619), .A4(new_n642), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n345), .B2(new_n367), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n810), .B2(new_n438), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n710), .A2(new_n632), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n721), .B(KEYINPUT110), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n437), .B(new_n809), .C1(new_n345), .C2(new_n367), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n812), .B1(new_n816), .B2(new_n808), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT110), .B1(new_n817), .B2(new_n721), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n807), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n801), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT112), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n795), .A2(KEYINPUT52), .A3(new_n797), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n798), .B2(KEYINPUT111), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n795), .A2(new_n826), .A3(KEYINPUT52), .A4(new_n797), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n586), .A2(new_n806), .A3(new_n633), .ZN(new_n829));
  INV_X1    g643(.A(new_n818), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n814), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n794), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n820), .A2(KEYINPUT112), .A3(KEYINPUT53), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n823), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n833), .B1(new_n801), .B2(new_n819), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n833), .B1(new_n794), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT114), .B1(new_n718), .B2(new_n793), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n828), .A2(new_n840), .A3(new_n841), .A4(new_n831), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT113), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n844), .B(new_n833), .C1(new_n801), .C2(new_n819), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n838), .A2(new_n842), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n836), .A2(KEYINPUT54), .B1(new_n846), .B2(KEYINPUT115), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(KEYINPUT115), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n764), .A2(new_n637), .A3(new_n675), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n792), .A2(new_n847), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OR2_X1    g664(.A1(G952), .A2(G953), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n651), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n495), .B1(new_n853), .B2(new_n649), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n765), .B(KEYINPUT49), .Z(new_n855));
  NOR3_X1   g669(.A1(new_n855), .A2(new_n694), .A3(new_n742), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n662), .A3(new_n727), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(G75));
  NAND3_X1  g672(.A1(new_n838), .A2(new_n842), .A3(new_n845), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n859), .A2(G902), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n482), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n449), .A2(new_n460), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT119), .Z(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT55), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(new_n458), .Z(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n861), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT56), .B1(new_n860), .B2(G210), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n865), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n219), .A2(G952), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(G51));
  INV_X1    g685(.A(new_n673), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n846), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n435), .B(KEYINPUT57), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT121), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT121), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n878), .B(new_n875), .C1(new_n873), .C2(new_n846), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n872), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n736), .B(KEYINPUT122), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n860), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n870), .B1(new_n880), .B2(new_n882), .ZN(G54));
  NAND3_X1  g697(.A1(new_n860), .A2(KEYINPUT58), .A3(G475), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n536), .A2(new_n537), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n870), .ZN(G60));
  NOR2_X1   g702(.A1(new_n602), .A2(new_n595), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n595), .B2(new_n604), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n847), .A2(new_n848), .ZN(new_n891));
  NAND2_X1  g705(.A1(G478), .A2(G902), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT59), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n874), .A2(new_n890), .A3(new_n893), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n870), .A3(new_n895), .ZN(G63));
  INV_X1    g710(.A(new_n870), .ZN(new_n897));
  NAND2_X1  g711(.A1(G217), .A2(G902), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT60), .Z(new_n899));
  NAND3_X1  g713(.A1(new_n859), .A2(new_n629), .A3(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n859), .A2(new_n899), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n226), .B(KEYINPUT123), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n897), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g718(.A(G953), .B1(new_n490), .B2(new_n456), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n829), .A2(new_n793), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(G953), .ZN(new_n907));
  INV_X1    g721(.A(new_n863), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(G898), .B2(new_n219), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n907), .B(new_n909), .ZN(G69));
  NAND2_X1  g724(.A1(new_n361), .A2(new_n318), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n520), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n743), .A2(new_n637), .A3(new_n665), .A4(new_n756), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n745), .A2(new_n754), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n799), .A2(new_n671), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n718), .A2(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n917), .A2(new_n721), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n219), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n219), .A2(G900), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(G953), .B1(new_n915), .B2(new_n918), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT126), .B1(new_n925), .B2(new_n922), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n913), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n418), .B2(new_n640), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT125), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n667), .A2(new_n795), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT62), .Z(new_n931));
  NOR4_X1   g745(.A1(new_n369), .A2(new_n804), .A3(new_n655), .A4(new_n710), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT124), .Z(new_n933));
  NAND4_X1  g747(.A1(new_n931), .A2(new_n745), .A3(new_n754), .A4(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n912), .B1(new_n934), .B2(new_n219), .ZN(new_n935));
  OR3_X1    g749(.A1(new_n927), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n927), .B2(new_n935), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(G72));
  NAND2_X1  g752(.A1(G472), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT63), .Z(new_n940));
  INV_X1    g754(.A(new_n906), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n919), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n364), .A2(new_n308), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n870), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT127), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n940), .B1(new_n934), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n658), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n943), .A2(new_n658), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n836), .A2(new_n940), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n945), .A2(new_n950), .ZN(G57));
endmodule


