

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U549 ( .A1(n680), .A2(n755), .ZN(n719) );
  INV_X1 U550 ( .A(n719), .ZN(n704) );
  INV_X1 U551 ( .A(n754), .ZN(n680) );
  NOR2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XOR2_X2 U553 ( .A(KEYINPUT17), .B(n514), .Z(n882) );
  NOR2_X1 U554 ( .A1(G1384), .A2(G164), .ZN(n679) );
  XNOR2_X1 U555 ( .A(n693), .B(n692), .ZN(n735) );
  INV_X1 U556 ( .A(KEYINPUT31), .ZN(n691) );
  XNOR2_X1 U557 ( .A(n691), .B(KEYINPUT98), .ZN(n692) );
  INV_X1 U558 ( .A(KEYINPUT96), .ZN(n681) );
  NOR2_X1 U559 ( .A1(G651), .A2(n620), .ZN(n640) );
  INV_X1 U560 ( .A(G2104), .ZN(n517) );
  NOR2_X1 U561 ( .A1(G2105), .A2(n517), .ZN(n879) );
  NAND2_X1 U562 ( .A1(G102), .A2(n879), .ZN(n516) );
  NAND2_X1 U563 ( .A1(G138), .A2(n882), .ZN(n515) );
  NAND2_X1 U564 ( .A1(n516), .A2(n515), .ZN(n522) );
  AND2_X1 U565 ( .A1(n517), .A2(G2105), .ZN(n874) );
  NAND2_X1 U566 ( .A1(G126), .A2(n874), .ZN(n520) );
  NAND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XOR2_X1 U568 ( .A(KEYINPUT66), .B(n518), .Z(n875) );
  NAND2_X1 U569 ( .A1(G114), .A2(n875), .ZN(n519) );
  NAND2_X1 U570 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U571 ( .A1(n522), .A2(n521), .ZN(G164) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n631) );
  NAND2_X1 U573 ( .A1(G85), .A2(n631), .ZN(n524) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n620) );
  INV_X1 U575 ( .A(G651), .ZN(n525) );
  NOR2_X1 U576 ( .A1(n620), .A2(n525), .ZN(n635) );
  NAND2_X1 U577 ( .A1(G72), .A2(n635), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n524), .A2(n523), .ZN(n530) );
  NOR2_X1 U579 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n526), .Z(n632) );
  NAND2_X1 U581 ( .A1(G60), .A2(n632), .ZN(n528) );
  NAND2_X1 U582 ( .A1(G47), .A2(n640), .ZN(n527) );
  NAND2_X1 U583 ( .A1(n528), .A2(n527), .ZN(n529) );
  OR2_X1 U584 ( .A1(n530), .A2(n529), .ZN(G290) );
  NAND2_X1 U585 ( .A1(G64), .A2(n632), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G52), .A2(n640), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U588 ( .A(KEYINPUT67), .B(n533), .Z(n538) );
  NAND2_X1 U589 ( .A1(G90), .A2(n631), .ZN(n535) );
  NAND2_X1 U590 ( .A1(G77), .A2(n635), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U592 ( .A(KEYINPUT9), .B(n536), .Z(n537) );
  NOR2_X1 U593 ( .A1(n538), .A2(n537), .ZN(G171) );
  AND2_X1 U594 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U595 ( .A(G132), .ZN(G219) );
  INV_X1 U596 ( .A(G82), .ZN(G220) );
  INV_X1 U597 ( .A(G108), .ZN(G238) );
  NAND2_X1 U598 ( .A1(G63), .A2(n632), .ZN(n540) );
  NAND2_X1 U599 ( .A1(G51), .A2(n640), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n542) );
  XOR2_X1 U601 ( .A(KEYINPUT79), .B(KEYINPUT6), .Z(n541) );
  XNOR2_X1 U602 ( .A(n542), .B(n541), .ZN(n551) );
  XNOR2_X1 U603 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G89), .A2(n631), .ZN(n543) );
  XNOR2_X1 U605 ( .A(n543), .B(KEYINPUT76), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n544), .B(KEYINPUT4), .ZN(n546) );
  NAND2_X1 U607 ( .A1(G76), .A2(n635), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n547), .B(KEYINPUT5), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n549), .B(n548), .ZN(n550) );
  NOR2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U612 ( .A(KEYINPUT7), .B(n552), .Z(G168) );
  XOR2_X1 U613 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U614 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n554) );
  NAND2_X1 U615 ( .A1(G7), .A2(G661), .ZN(n553) );
  XNOR2_X1 U616 ( .A(n554), .B(n553), .ZN(G223) );
  INV_X1 U617 ( .A(G223), .ZN(n820) );
  NAND2_X1 U618 ( .A1(n820), .A2(G567), .ZN(n555) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(n555), .Z(G234) );
  XNOR2_X1 U620 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G81), .A2(n631), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(KEYINPUT12), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT70), .ZN(n559) );
  NAND2_X1 U624 ( .A1(G68), .A2(n635), .ZN(n558) );
  NAND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n561), .B(n560), .ZN(n564) );
  NAND2_X1 U627 ( .A1(n632), .A2(G56), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n562), .Z(n563) );
  NOR2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n640), .A2(G43), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n962) );
  INV_X1 U632 ( .A(G860), .ZN(n589) );
  NOR2_X1 U633 ( .A1(n962), .A2(n589), .ZN(n567) );
  XOR2_X1 U634 ( .A(KEYINPUT72), .B(n567), .Z(G153) );
  XNOR2_X1 U635 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G66), .A2(n632), .ZN(n568) );
  XNOR2_X1 U638 ( .A(n568), .B(KEYINPUT74), .ZN(n575) );
  NAND2_X1 U639 ( .A1(G92), .A2(n631), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G54), .A2(n640), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G79), .A2(n635), .ZN(n571) );
  XNOR2_X1 U643 ( .A(KEYINPUT75), .B(n571), .ZN(n572) );
  NOR2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n576), .Z(n971) );
  INV_X1 U647 ( .A(G868), .ZN(n654) );
  NAND2_X1 U648 ( .A1(n971), .A2(n654), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n578), .A2(n577), .ZN(G284) );
  NAND2_X1 U650 ( .A1(G65), .A2(n632), .ZN(n580) );
  NAND2_X1 U651 ( .A1(G53), .A2(n640), .ZN(n579) );
  NAND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U653 ( .A(KEYINPUT68), .B(n581), .Z(n585) );
  NAND2_X1 U654 ( .A1(G91), .A2(n631), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G78), .A2(n635), .ZN(n582) );
  AND2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G299) );
  NOR2_X1 U658 ( .A1(G286), .A2(n654), .ZN(n587) );
  NOR2_X1 U659 ( .A1(G868), .A2(G299), .ZN(n586) );
  NOR2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U661 ( .A(KEYINPUT80), .B(n588), .ZN(G297) );
  NAND2_X1 U662 ( .A1(n589), .A2(G559), .ZN(n590) );
  INV_X1 U663 ( .A(n971), .ZN(n606) );
  NAND2_X1 U664 ( .A1(n590), .A2(n606), .ZN(n591) );
  XNOR2_X1 U665 ( .A(n591), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n962), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT81), .B(n592), .Z(n595) );
  NAND2_X1 U668 ( .A1(G868), .A2(n606), .ZN(n593) );
  NOR2_X1 U669 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U670 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U671 ( .A1(G123), .A2(n874), .ZN(n596) );
  XNOR2_X1 U672 ( .A(n596), .B(KEYINPUT18), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT82), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G99), .A2(n879), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G135), .A2(n882), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G111), .A2(n875), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(n917) );
  XNOR2_X1 U680 ( .A(G2096), .B(n917), .ZN(n605) );
  INV_X1 U681 ( .A(G2100), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G156) );
  NAND2_X1 U683 ( .A1(n606), .A2(G559), .ZN(n651) );
  XNOR2_X1 U684 ( .A(n962), .B(n651), .ZN(n607) );
  NOR2_X1 U685 ( .A1(n607), .A2(G860), .ZN(n616) );
  NAND2_X1 U686 ( .A1(G93), .A2(n631), .ZN(n609) );
  NAND2_X1 U687 ( .A1(G80), .A2(n635), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U689 ( .A(n610), .B(KEYINPUT83), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G55), .A2(n640), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n632), .A2(G67), .ZN(n613) );
  XOR2_X1 U693 ( .A(KEYINPUT84), .B(n613), .Z(n614) );
  OR2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n653) );
  XOR2_X1 U695 ( .A(n616), .B(n653), .Z(G145) );
  NAND2_X1 U696 ( .A1(G49), .A2(n640), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U699 ( .A1(n632), .A2(n619), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n620), .A2(G87), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(G288) );
  NAND2_X1 U702 ( .A1(G62), .A2(n632), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G50), .A2(n640), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G88), .A2(n631), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G75), .A2(n635), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT87), .B(n627), .Z(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U710 ( .A(KEYINPUT88), .B(n630), .Z(G303) );
  NAND2_X1 U711 ( .A1(G86), .A2(n631), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G61), .A2(n632), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n635), .A2(G73), .ZN(n636) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(n636), .Z(n637) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U717 ( .A(KEYINPUT85), .B(n639), .Z(n642) );
  NAND2_X1 U718 ( .A1(n640), .A2(G48), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U720 ( .A(KEYINPUT86), .B(n643), .ZN(G305) );
  XNOR2_X1 U721 ( .A(KEYINPUT19), .B(KEYINPUT89), .ZN(n645) );
  XOR2_X1 U722 ( .A(G288), .B(n653), .Z(n644) );
  XNOR2_X1 U723 ( .A(n645), .B(n644), .ZN(n649) );
  XNOR2_X1 U724 ( .A(G303), .B(G305), .ZN(n647) );
  INV_X1 U725 ( .A(G299), .ZN(n969) );
  XNOR2_X1 U726 ( .A(n962), .B(n969), .ZN(n646) );
  XNOR2_X1 U727 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n650), .B(G290), .ZN(n893) );
  XNOR2_X1 U730 ( .A(n651), .B(n893), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n652), .A2(G868), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U734 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U735 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U736 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U737 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U738 ( .A1(n660), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U740 ( .A1(G69), .A2(G120), .ZN(n661) );
  XNOR2_X1 U741 ( .A(KEYINPUT90), .B(n661), .ZN(n662) );
  NOR2_X1 U742 ( .A1(G238), .A2(n662), .ZN(n663) );
  NAND2_X1 U743 ( .A1(G57), .A2(n663), .ZN(n826) );
  NAND2_X1 U744 ( .A1(n826), .A2(G567), .ZN(n668) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT22), .B(n664), .Z(n665) );
  NOR2_X1 U747 ( .A1(G218), .A2(n665), .ZN(n666) );
  NAND2_X1 U748 ( .A1(G96), .A2(n666), .ZN(n825) );
  NAND2_X1 U749 ( .A1(n825), .A2(G2106), .ZN(n667) );
  NAND2_X1 U750 ( .A1(n668), .A2(n667), .ZN(n828) );
  NAND2_X1 U751 ( .A1(G483), .A2(G661), .ZN(n669) );
  NOR2_X1 U752 ( .A1(n828), .A2(n669), .ZN(n824) );
  NAND2_X1 U753 ( .A1(n824), .A2(G36), .ZN(n670) );
  XOR2_X1 U754 ( .A(KEYINPUT91), .B(n670), .Z(G176) );
  NAND2_X1 U755 ( .A1(G101), .A2(n879), .ZN(n671) );
  XOR2_X1 U756 ( .A(KEYINPUT23), .B(n671), .Z(n674) );
  NAND2_X1 U757 ( .A1(G125), .A2(n874), .ZN(n672) );
  XOR2_X1 U758 ( .A(KEYINPUT65), .B(n672), .Z(n673) );
  NAND2_X1 U759 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U760 ( .A1(G137), .A2(n882), .ZN(n676) );
  NAND2_X1 U761 ( .A1(G113), .A2(n875), .ZN(n675) );
  NAND2_X1 U762 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U763 ( .A1(n678), .A2(n677), .ZN(G160) );
  XNOR2_X1 U764 ( .A(n679), .B(KEYINPUT64), .ZN(n754) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n755) );
  NOR2_X1 U766 ( .A1(G2084), .A2(n719), .ZN(n734) );
  NAND2_X1 U767 ( .A1(G8), .A2(n719), .ZN(n795) );
  NOR2_X1 U768 ( .A1(G1966), .A2(n795), .ZN(n682) );
  XNOR2_X1 U769 ( .A(n682), .B(n681), .ZN(n738) );
  NAND2_X1 U770 ( .A1(n738), .A2(G8), .ZN(n683) );
  NOR2_X1 U771 ( .A1(n734), .A2(n683), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT30), .B(n684), .Z(n685) );
  NOR2_X1 U773 ( .A1(G168), .A2(n685), .ZN(n690) );
  INV_X1 U774 ( .A(G1961), .ZN(n1003) );
  NAND2_X1 U775 ( .A1(n719), .A2(n1003), .ZN(n687) );
  XNOR2_X1 U776 ( .A(G2078), .B(KEYINPUT25), .ZN(n944) );
  NAND2_X1 U777 ( .A1(n704), .A2(n944), .ZN(n686) );
  NAND2_X1 U778 ( .A1(n687), .A2(n686), .ZN(n694) );
  NOR2_X1 U779 ( .A1(G171), .A2(n694), .ZN(n688) );
  XOR2_X1 U780 ( .A(KEYINPUT97), .B(n688), .Z(n689) );
  NOR2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n694), .A2(G171), .ZN(n718) );
  NAND2_X1 U783 ( .A1(n704), .A2(G2072), .ZN(n695) );
  XNOR2_X1 U784 ( .A(n695), .B(KEYINPUT27), .ZN(n697) );
  INV_X1 U785 ( .A(G1956), .ZN(n994) );
  NOR2_X1 U786 ( .A1(n994), .A2(n704), .ZN(n696) );
  NOR2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n699) );
  NOR2_X1 U788 ( .A1(n969), .A2(n699), .ZN(n698) );
  XOR2_X1 U789 ( .A(n698), .B(KEYINPUT28), .Z(n715) );
  NAND2_X1 U790 ( .A1(n969), .A2(n699), .ZN(n713) );
  INV_X1 U791 ( .A(G1996), .ZN(n945) );
  NOR2_X1 U792 ( .A1(n719), .A2(n945), .ZN(n700) );
  XOR2_X1 U793 ( .A(n700), .B(KEYINPUT26), .Z(n702) );
  NAND2_X1 U794 ( .A1(n719), .A2(G1341), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U796 ( .A1(n962), .A2(n703), .ZN(n708) );
  NAND2_X1 U797 ( .A1(G1348), .A2(n719), .ZN(n706) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n704), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U800 ( .A1(n971), .A2(n709), .ZN(n707) );
  OR2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n971), .A2(n709), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U806 ( .A(KEYINPUT29), .B(n716), .Z(n717) );
  NAND2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n736) );
  INV_X1 U808 ( .A(G8), .ZN(n726) );
  NOR2_X1 U809 ( .A1(G1971), .A2(n795), .ZN(n721) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n719), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U812 ( .A(KEYINPUT99), .B(n722), .Z(n723) );
  NAND2_X1 U813 ( .A1(G303), .A2(n723), .ZN(n724) );
  XNOR2_X1 U814 ( .A(n724), .B(KEYINPUT100), .ZN(n725) );
  OR2_X1 U815 ( .A1(n726), .A2(n725), .ZN(n728) );
  AND2_X1 U816 ( .A1(n736), .A2(n728), .ZN(n727) );
  NAND2_X1 U817 ( .A1(n735), .A2(n727), .ZN(n732) );
  INV_X1 U818 ( .A(n728), .ZN(n730) );
  AND2_X1 U819 ( .A1(G286), .A2(G8), .ZN(n729) );
  OR2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U822 ( .A(n733), .B(KEYINPUT32), .ZN(n742) );
  NAND2_X1 U823 ( .A1(G8), .A2(n734), .ZN(n740) );
  NAND2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n737) );
  AND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n791) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U829 ( .A1(G303), .A2(G1971), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n749), .A2(n743), .ZN(n982) );
  NAND2_X1 U831 ( .A1(n791), .A2(n982), .ZN(n746) );
  INV_X1 U832 ( .A(KEYINPUT33), .ZN(n744) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n967) );
  AND2_X1 U834 ( .A1(n744), .A2(n967), .ZN(n745) );
  AND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  INV_X1 U836 ( .A(n795), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n747), .A2(n748), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U841 ( .A(KEYINPUT101), .B(n753), .Z(n788) );
  XOR2_X1 U842 ( .A(G305), .B(G1981), .Z(n976) );
  NOR2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n814) );
  XNOR2_X1 U844 ( .A(G2067), .B(KEYINPUT37), .ZN(n807) );
  XNOR2_X1 U845 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n759) );
  NAND2_X1 U846 ( .A1(G104), .A2(n879), .ZN(n757) );
  NAND2_X1 U847 ( .A1(G140), .A2(n882), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U849 ( .A(n759), .B(n758), .ZN(n764) );
  NAND2_X1 U850 ( .A1(G128), .A2(n874), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G116), .A2(n875), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U853 ( .A(KEYINPUT35), .B(n762), .Z(n763) );
  NOR2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U855 ( .A(KEYINPUT36), .B(n765), .ZN(n890) );
  NOR2_X1 U856 ( .A1(n807), .A2(n890), .ZN(n923) );
  NAND2_X1 U857 ( .A1(n814), .A2(n923), .ZN(n766) );
  XOR2_X1 U858 ( .A(KEYINPUT93), .B(n766), .Z(n805) );
  NAND2_X1 U859 ( .A1(G119), .A2(n874), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G95), .A2(n879), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n875), .A2(G107), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n769), .B(KEYINPUT94), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n882), .A2(G131), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n772) );
  OR2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n887) );
  AND2_X1 U867 ( .A1(n887), .A2(G1991), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G117), .A2(n875), .ZN(n780) );
  NAND2_X1 U869 ( .A1(G129), .A2(n874), .ZN(n775) );
  NAND2_X1 U870 ( .A1(G141), .A2(n882), .ZN(n774) );
  NAND2_X1 U871 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n879), .A2(G105), .ZN(n776) );
  XOR2_X1 U873 ( .A(KEYINPUT38), .B(n776), .Z(n777) );
  NOR2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U876 ( .A(KEYINPUT95), .B(n781), .ZN(n871) );
  NOR2_X1 U877 ( .A1(n871), .A2(n945), .ZN(n782) );
  NOR2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n921) );
  INV_X1 U879 ( .A(n814), .ZN(n784) );
  NOR2_X1 U880 ( .A1(n921), .A2(n784), .ZN(n802) );
  INV_X1 U881 ( .A(n802), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n805), .A2(n785), .ZN(n799) );
  INV_X1 U883 ( .A(n799), .ZN(n786) );
  AND2_X1 U884 ( .A1(n976), .A2(n786), .ZN(n787) );
  NAND2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n812) );
  NOR2_X1 U886 ( .A1(G2090), .A2(G303), .ZN(n789) );
  NAND2_X1 U887 ( .A1(G8), .A2(n789), .ZN(n790) );
  NAND2_X1 U888 ( .A1(n791), .A2(n790), .ZN(n792) );
  AND2_X1 U889 ( .A1(n792), .A2(n795), .ZN(n797) );
  NOR2_X1 U890 ( .A1(G305), .A2(G1981), .ZN(n793) );
  XOR2_X1 U891 ( .A(n793), .B(KEYINPUT24), .Z(n794) );
  NOR2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n810) );
  AND2_X1 U895 ( .A1(n945), .A2(n871), .ZN(n930) );
  NOR2_X1 U896 ( .A1(G1991), .A2(n887), .ZN(n918) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U898 ( .A1(n918), .A2(n800), .ZN(n801) );
  NOR2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n930), .A2(n803), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n804), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n807), .A2(n890), .ZN(n927) );
  NAND2_X1 U904 ( .A1(n808), .A2(n927), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n809), .A2(n814), .ZN(n813) );
  AND2_X1 U906 ( .A1(n810), .A2(n813), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n818) );
  INV_X1 U908 ( .A(n813), .ZN(n816) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n966) );
  NAND2_X1 U910 ( .A1(n966), .A2(n814), .ZN(n815) );
  OR2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  AND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U913 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  INV_X1 U914 ( .A(G303), .ZN(G166) );
  NAND2_X1 U915 ( .A1(n820), .A2(G2106), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n821), .Z(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U918 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U921 ( .A(G120), .B(KEYINPUT104), .Z(G236) );
  XNOR2_X1 U922 ( .A(G96), .B(KEYINPUT105), .ZN(G221) );
  NOR2_X1 U924 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n827), .B(KEYINPUT106), .ZN(G325) );
  XNOR2_X1 U926 ( .A(KEYINPUT107), .B(G325), .ZN(G261) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  INV_X1 U928 ( .A(n828), .ZN(G319) );
  XOR2_X1 U929 ( .A(KEYINPUT112), .B(G1976), .Z(n830) );
  XNOR2_X1 U930 ( .A(G1986), .B(G1956), .ZN(n829) );
  XNOR2_X1 U931 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U932 ( .A(n831), .B(KEYINPUT41), .Z(n833) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1991), .ZN(n832) );
  XNOR2_X1 U934 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U935 ( .A(G1981), .B(G1971), .Z(n835) );
  XNOR2_X1 U936 ( .A(G1966), .B(G1961), .ZN(n834) );
  XNOR2_X1 U937 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U938 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U939 ( .A(KEYINPUT111), .B(G2474), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(G229) );
  XOR2_X1 U941 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n841) );
  XNOR2_X1 U942 ( .A(KEYINPUT109), .B(G2096), .ZN(n840) );
  XNOR2_X1 U943 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U944 ( .A(n842), .B(KEYINPUT42), .Z(n844) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2084), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U947 ( .A(G2100), .B(G2090), .Z(n846) );
  XNOR2_X1 U948 ( .A(G2078), .B(G2072), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U950 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U951 ( .A(G2678), .B(KEYINPUT108), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(G227) );
  NAND2_X1 U953 ( .A1(G124), .A2(n874), .ZN(n851) );
  XNOR2_X1 U954 ( .A(n851), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n875), .A2(G112), .ZN(n852) );
  XOR2_X1 U956 ( .A(KEYINPUT113), .B(n852), .Z(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G100), .A2(n879), .ZN(n856) );
  NAND2_X1 U959 ( .A1(G136), .A2(n882), .ZN(n855) );
  NAND2_X1 U960 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U961 ( .A1(n858), .A2(n857), .ZN(G162) );
  XOR2_X1 U962 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n860) );
  XNOR2_X1 U963 ( .A(G164), .B(n917), .ZN(n859) );
  XNOR2_X1 U964 ( .A(n860), .B(n859), .ZN(n870) );
  NAND2_X1 U965 ( .A1(G130), .A2(n874), .ZN(n862) );
  NAND2_X1 U966 ( .A1(G118), .A2(n875), .ZN(n861) );
  NAND2_X1 U967 ( .A1(n862), .A2(n861), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G106), .A2(n879), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G142), .A2(n882), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U971 ( .A(KEYINPUT114), .B(n865), .Z(n866) );
  XNOR2_X1 U972 ( .A(KEYINPUT45), .B(n866), .ZN(n867) );
  NOR2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U974 ( .A(n870), .B(n869), .Z(n873) );
  XNOR2_X1 U975 ( .A(G160), .B(n871), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n873), .B(n872), .ZN(n886) );
  NAND2_X1 U977 ( .A1(G127), .A2(n874), .ZN(n877) );
  NAND2_X1 U978 ( .A1(G115), .A2(n875), .ZN(n876) );
  NAND2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U980 ( .A(n878), .B(KEYINPUT47), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G103), .A2(n879), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G139), .A2(n882), .ZN(n883) );
  XNOR2_X1 U984 ( .A(KEYINPUT115), .B(n883), .ZN(n884) );
  NOR2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n913) );
  XOR2_X1 U986 ( .A(n886), .B(n913), .Z(n889) );
  XOR2_X1 U987 ( .A(n887), .B(G162), .Z(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U989 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U990 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G286), .B(n971), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U993 ( .A(n895), .B(G171), .ZN(n896) );
  NOR2_X1 U994 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U995 ( .A(G2438), .B(KEYINPUT102), .Z(n898) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2430), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U998 ( .A(n899), .B(G2435), .Z(n901) );
  XNOR2_X1 U999 ( .A(G1341), .B(G1348), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U1001 ( .A(G2451), .B(G2427), .Z(n903) );
  XNOR2_X1 U1002 ( .A(G2454), .B(G2446), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(n905), .B(n904), .Z(n906) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n906), .ZN(n912) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n912), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n907) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n911) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G57), .ZN(G237) );
  INV_X1 U1014 ( .A(n912), .ZN(G401) );
  XOR2_X1 U1015 ( .A(G2072), .B(n913), .Z(n915) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1018 ( .A(KEYINPUT50), .B(n916), .Z(n936) );
  XNOR2_X1 U1019 ( .A(G160), .B(G2084), .ZN(n925) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(n919), .B(KEYINPUT116), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n926), .B(KEYINPUT117), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n933) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n931), .B(KEYINPUT51), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1031 ( .A(KEYINPUT118), .B(n934), .Z(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(n937), .B(KEYINPUT52), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n959) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n959), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(KEYINPUT120), .B(n939), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(G1991), .B(G25), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n952) );
  XOR2_X1 U1041 ( .A(G2072), .B(G33), .Z(n943) );
  NAND2_X1 U1042 ( .A1(n943), .A2(G28), .ZN(n950) );
  XOR2_X1 U1043 ( .A(n944), .B(G27), .Z(n947) );
  XOR2_X1 U1044 ( .A(n945), .B(G32), .Z(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT121), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1049 ( .A(n953), .B(KEYINPUT53), .ZN(n956) );
  XOR2_X1 U1050 ( .A(G2084), .B(G34), .Z(n954) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(n954), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G35), .B(G2090), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(n959), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(G29), .A2(n961), .ZN(n1019) );
  XOR2_X1 U1057 ( .A(G16), .B(KEYINPUT56), .Z(n986) );
  NAND2_X1 U1058 ( .A1(G303), .A2(G1971), .ZN(n964) );
  XOR2_X1 U1059 ( .A(G1341), .B(n962), .Z(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n984) );
  XNOR2_X1 U1063 ( .A(n969), .B(G1956), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(n970), .B(KEYINPUT122), .ZN(n975) );
  XOR2_X1 U1065 ( .A(G171), .B(G1961), .Z(n973) );
  XNOR2_X1 U1066 ( .A(n971), .B(G1348), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1071 ( .A(KEYINPUT57), .B(n978), .Z(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NOR2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n1015) );
  XOR2_X1 U1076 ( .A(G16), .B(KEYINPUT123), .Z(n1013) );
  XNOR2_X1 U1077 ( .A(G1986), .B(G24), .ZN(n991) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G22), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(G1976), .B(G23), .ZN(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(KEYINPUT125), .B(n989), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT126), .B(n992), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(n993), .B(KEYINPUT58), .ZN(n1010) );
  XNOR2_X1 U1085 ( .A(G20), .B(n994), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G6), .B(G1981), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT59), .B(G1348), .Z(n999) );
  XNOR2_X1 U1091 ( .A(G4), .B(n999), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1002), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1003), .B(G5), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(KEYINPUT124), .B(G1966), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(G21), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(n1011), .B(KEYINPUT61), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1016), .Z(n1017) );
  NAND2_X1 U1104 ( .A1(G11), .A2(n1017), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

