//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n204));
  NAND2_X1  g0004(.A1(G87), .A2(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT64), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(new_n208), .A2(new_n209), .B1(G77), .B2(G244), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G116), .A2(G270), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G68), .A2(G238), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  AND2_X1   g0014(.A1(G50), .A2(G226), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n203), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n203), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT0), .Z(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR3_X1   g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n217), .A2(new_n220), .A3(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G270), .ZN(new_n232));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n230), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  INV_X1    g0036(.A(G107), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NOR2_X1   g0044(.A1(G20), .A2(G33), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n245), .A2(G50), .B1(G20), .B2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT69), .B1(new_n248), .B2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT69), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(new_n222), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n247), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n223), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n257), .B(KEYINPUT11), .Z(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n256), .B1(new_n259), .B2(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n246), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n263), .A2(new_n222), .A3(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n246), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT12), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n258), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G33), .ZN(new_n271));
  AND2_X1   g0071(.A1(G232), .A2(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G97), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n269), .A2(new_n271), .A3(G226), .A4(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n269), .A2(new_n271), .A3(new_n272), .A4(KEYINPUT72), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n275), .A2(new_n276), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(G1), .B(G13), .C1(new_n248), .C2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n285));
  INV_X1    g0085(.A(G274), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT66), .B(G41), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI211_X1 g0088(.A(G1), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT67), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT67), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n282), .A2(new_n293), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n289), .B1(new_n295), .B2(G238), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT73), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n280), .A2(new_n297), .A3(new_n283), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n285), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT74), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT13), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n285), .A2(new_n302), .A3(new_n296), .A4(new_n298), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n299), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(G169), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT14), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n304), .A2(KEYINPUT14), .A3(G169), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n300), .A2(G179), .A3(new_n303), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT76), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(KEYINPUT76), .A3(new_n311), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n268), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n304), .A2(G200), .A3(new_n305), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n300), .A2(G190), .A3(new_n303), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n268), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT75), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n289), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n295), .A2(G226), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n269), .A2(new_n271), .ZN(new_n325));
  MUX2_X1   g0125(.A(G222), .B(G223), .S(G1698), .Z(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n253), .B2(new_n325), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT68), .Z(new_n329));
  OAI211_X1 g0129(.A(new_n323), .B(new_n324), .C1(new_n329), .C2(new_n282), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  NOR2_X1   g0131(.A1(G58), .A2(G68), .ZN(new_n332));
  INV_X1    g0132(.A(G50), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n222), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(G150), .B2(new_n245), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n252), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(new_n256), .B1(new_n333), .B2(new_n264), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n333), .B2(new_n261), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT9), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n331), .B(new_n340), .C1(new_n341), .C2(new_n330), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT10), .ZN(new_n343));
  INV_X1    g0143(.A(G169), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n330), .A2(new_n344), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n339), .C1(G179), .C2(new_n330), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n269), .A2(new_n271), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT7), .B1(new_n348), .B2(new_n222), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT78), .B1(new_n270), .B2(G33), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT78), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(new_n248), .A3(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n350), .A2(new_n352), .A3(new_n271), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT79), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT79), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n358), .A3(new_n355), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n349), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT80), .B1(new_n360), .B2(new_n246), .ZN(new_n361));
  INV_X1    g0161(.A(G58), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n246), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n332), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n245), .A2(G159), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n354), .B1(new_n325), .B2(G20), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n353), .A2(new_n358), .A3(new_n355), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n358), .B1(new_n353), .B2(new_n355), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT80), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n372), .A3(G68), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n361), .A2(new_n367), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n366), .B(KEYINPUT77), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n348), .A2(new_n355), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n378), .B2(new_n349), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n256), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n291), .A2(new_n227), .ZN(new_n384));
  XOR2_X1   g0184(.A(new_n384), .B(KEYINPUT81), .Z(new_n385));
  OAI21_X1  g0185(.A(new_n325), .B1(G226), .B2(new_n277), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  INV_X1    g0187(.A(G87), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n386), .A2(new_n387), .B1(new_n248), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n289), .B1(new_n389), .B2(new_n283), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G200), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n385), .A2(new_n390), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G190), .ZN(new_n394));
  INV_X1    g0194(.A(new_n336), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(new_n264), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n396), .B1(new_n261), .B2(new_n395), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n383), .A2(new_n392), .A3(new_n394), .A4(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n381), .B1(new_n374), .B2(new_n375), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n397), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n403), .A2(KEYINPUT17), .A3(new_n392), .A4(new_n394), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n393), .A2(new_n344), .ZN(new_n406));
  INV_X1    g0206(.A(G179), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n391), .A2(new_n407), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n402), .A2(new_n397), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT18), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G20), .A2(G77), .ZN(new_n411));
  INV_X1    g0211(.A(new_n245), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT15), .B(G87), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n411), .B1(new_n336), .B2(new_n412), .C1(new_n252), .C2(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(new_n256), .B1(new_n253), .B2(new_n264), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n253), .B2(new_n261), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n289), .B1(new_n295), .B2(G244), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G238), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n325), .B(new_n418), .C1(new_n227), .C2(G1698), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT70), .B(G107), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n325), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n417), .B1(new_n282), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n416), .B1(G200), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT71), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n341), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n347), .A2(new_n405), .A3(new_n410), .A4(new_n428), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n422), .A2(G179), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n422), .A2(new_n344), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n416), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n322), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G283), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n222), .C1(G33), .C2(new_n206), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n256), .B1(new_n222), .B2(G116), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT84), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(new_n437), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT20), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT85), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n440), .A2(new_n441), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT85), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n445), .A3(new_n441), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n443), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n256), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(G1), .B2(new_n248), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n264), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G116), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n264), .A2(new_n239), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n288), .A2(G1), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(new_n287), .C2(KEYINPUT5), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n456), .A2(new_n282), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G270), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n456), .A2(new_n286), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G264), .A2(G1698), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n325), .B(new_n461), .C1(new_n207), .C2(G1698), .ZN(new_n462));
  XOR2_X1   g0262(.A(KEYINPUT83), .B(G303), .Z(new_n463));
  OAI211_X1 g0263(.A(new_n462), .B(new_n283), .C1(new_n325), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n458), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G200), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n465), .A2(new_n341), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n453), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n466), .A2(new_n344), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n453), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT21), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT86), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n465), .A2(new_n407), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n453), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(KEYINPUT86), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n453), .A2(new_n477), .A3(new_n471), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n325), .B1(G257), .B2(new_n277), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G250), .A2(G1698), .ZN(new_n480));
  INV_X1    g0280(.A(G294), .ZN(new_n481));
  OAI22_X1  g0281(.A1(new_n479), .A2(new_n480), .B1(new_n248), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n283), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n457), .A2(G264), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n460), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G179), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n344), .B2(new_n485), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT22), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n489));
  OAI21_X1  g0289(.A(G87), .B1(new_n488), .B2(KEYINPUT87), .ZN(new_n490));
  OR4_X1    g0290(.A1(G20), .A2(new_n348), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n325), .A2(new_n222), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n492), .B2(new_n490), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  XOR2_X1   g0294(.A(KEYINPUT89), .B(KEYINPUT23), .Z(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n222), .B2(new_n420), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n222), .A2(G33), .A3(G116), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT88), .ZN(new_n498));
  OR3_X1    g0298(.A1(new_n222), .A2(KEYINPUT23), .A3(G107), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT24), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n494), .A2(KEYINPUT24), .A3(new_n500), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n256), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n450), .A2(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n264), .A2(new_n237), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT25), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n505), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n487), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n474), .A2(new_n476), .A3(new_n478), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n504), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT24), .B1(new_n494), .B2(new_n500), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n508), .B1(new_n515), .B2(new_n256), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n485), .A2(G200), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n483), .A2(new_n484), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(G190), .A3(new_n460), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n516), .A2(new_n506), .A3(new_n517), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n450), .A2(G97), .ZN(new_n521));
  INV_X1    g0321(.A(new_n264), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT6), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n523), .A2(new_n206), .A3(G107), .ZN(new_n524));
  XNOR2_X1  g0324(.A(G97), .B(G107), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n526), .A2(new_n222), .B1(new_n253), .B2(new_n412), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n527), .B1(new_n371), .B2(new_n420), .ZN(new_n528));
  OAI221_X1 g0328(.A(new_n521), .B1(G97), .B2(new_n522), .C1(new_n528), .C2(new_n448), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n325), .A2(KEYINPUT4), .A3(G244), .A4(new_n277), .ZN(new_n531));
  INV_X1    g0331(.A(G244), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n348), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n531), .B(new_n434), .C1(KEYINPUT4), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n325), .A2(G250), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n277), .B1(new_n535), .B2(KEYINPUT4), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n283), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n459), .B1(new_n457), .B2(G257), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n539), .A2(new_n467), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(G190), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n530), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n539), .A2(new_n407), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n529), .B(new_n543), .C1(G169), .C2(new_n539), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n532), .A2(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n325), .B(new_n545), .C1(G238), .C2(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n282), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n282), .B1(G250), .B2(new_n455), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n286), .B2(new_n455), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n551), .A2(new_n467), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(G190), .B2(new_n551), .ZN(new_n553));
  NOR3_X1   g0353(.A1(new_n449), .A2(new_n388), .A3(new_n264), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n554), .B(KEYINPUT82), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(new_n252), .B2(new_n206), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n222), .B1(new_n276), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n388), .A2(new_n206), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n558), .B1(new_n420), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n557), .B(new_n560), .C1(new_n246), .C2(new_n492), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n256), .B1(new_n264), .B2(new_n413), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n551), .ZN(new_n564));
  INV_X1    g0364(.A(new_n413), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n450), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n564), .A2(new_n344), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n551), .A2(new_n407), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n553), .A2(new_n563), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n520), .A2(new_n542), .A3(new_n544), .A4(new_n569), .ZN(new_n570));
  NOR4_X1   g0370(.A1(new_n433), .A2(new_n470), .A3(new_n512), .A4(new_n570), .ZN(G372));
  INV_X1    g0371(.A(new_n433), .ZN(new_n572));
  INV_X1    g0372(.A(new_n569), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n573), .A2(new_n544), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n574), .B(KEYINPUT26), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n567), .A2(new_n568), .ZN(new_n576));
  INV_X1    g0376(.A(new_n570), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n512), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n572), .A2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n268), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT76), .B1(new_n310), .B2(new_n311), .ZN(new_n582));
  INV_X1    g0382(.A(new_n311), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n313), .B(new_n583), .C1(new_n308), .C2(new_n309), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n432), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n320), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n405), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n410), .A2(KEYINPUT90), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n410), .A2(KEYINPUT90), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n343), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT91), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n592), .A2(new_n593), .A3(new_n346), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n592), .B2(new_n346), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n580), .B1(new_n594), .B2(new_n595), .ZN(G369));
  NOR2_X1   g0396(.A1(new_n263), .A2(G20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n259), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT92), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT27), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(G213), .ZN(new_n603));
  INV_X1    g0403(.A(G343), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n453), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g0406(.A(new_n606), .B(KEYINPUT93), .Z(new_n607));
  NAND3_X1  g0407(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n608));
  OR3_X1    g0408(.A1(new_n607), .A2(new_n608), .A3(new_n470), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n610), .A2(KEYINPUT94), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(KEYINPUT94), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(G330), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT95), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n511), .A2(new_n605), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n510), .A2(new_n605), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n520), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n487), .A2(new_n510), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n616), .B(new_n618), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n520), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT95), .B1(new_n623), .B2(new_n617), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n605), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n608), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT96), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n608), .A2(KEYINPUT96), .A3(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n617), .B1(new_n632), .B2(new_n625), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n626), .A2(new_n633), .ZN(G399));
  INV_X1    g0434(.A(new_n287), .ZN(new_n635));
  INV_X1    g0435(.A(new_n218), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n420), .A2(G116), .A3(new_n559), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G1), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n221), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT28), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n579), .A2(new_n627), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT29), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR4_X1   g0445(.A1(new_n512), .A2(new_n570), .A3(new_n470), .A4(new_n605), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n539), .A2(new_n518), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(KEYINPUT30), .A3(new_n475), .A4(new_n551), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n539), .A2(new_n466), .A3(G179), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n485), .A3(new_n564), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n539), .A2(new_n475), .A3(new_n518), .A4(new_n551), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT30), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n605), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT31), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(KEYINPUT31), .A3(new_n605), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n646), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G330), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n579), .A2(new_n627), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT29), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n645), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n642), .B1(new_n667), .B2(G1), .ZN(G364));
  NAND2_X1  g0468(.A1(new_n597), .A2(G45), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n638), .A2(G1), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n615), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(G330), .B2(new_n613), .ZN(new_n673));
  NOR2_X1   g0473(.A1(G13), .A2(G33), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G20), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n613), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n222), .B1(KEYINPUT97), .B2(new_n344), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n344), .A2(KEYINPUT97), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n223), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n407), .A2(new_n467), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n222), .A2(G190), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(G317), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT33), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n686), .A2(KEYINPUT33), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(G179), .A2(G200), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G329), .ZN(new_n693));
  INV_X1    g0493(.A(G283), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n467), .A2(G179), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n683), .A2(new_n695), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n689), .B(new_n693), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n222), .A2(new_n341), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n682), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n697), .B1(G326), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n695), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G303), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n407), .A2(G200), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n325), .B1(new_n707), .B2(G322), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n222), .B1(new_n690), .B2(G190), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G294), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n701), .A2(new_n704), .A3(new_n708), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n683), .A2(new_n705), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(G311), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n699), .A2(new_n333), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n709), .A2(new_n206), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n348), .B(new_n717), .C1(G58), .C2(new_n707), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n703), .A2(G87), .ZN(new_n719));
  INV_X1    g0519(.A(G159), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n691), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT32), .ZN(new_n722));
  INV_X1    g0522(.A(new_n696), .ZN(new_n723));
  AOI22_X1  g0523(.A1(G77), .A2(new_n714), .B1(new_n723), .B2(G107), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n718), .A2(new_n719), .A3(new_n722), .A4(new_n724), .ZN(new_n725));
  AOI211_X1 g0525(.A(new_n716), .B(new_n725), .C1(G68), .C2(new_n685), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n681), .B1(new_n715), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n243), .A2(G45), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n325), .A2(new_n636), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n728), .B(new_n729), .C1(G45), .C2(new_n221), .ZN(new_n730));
  INV_X1    g0530(.A(G355), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n325), .A2(new_n218), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n730), .B1(G116), .B2(new_n218), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n681), .A2(new_n676), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n678), .A2(new_n727), .A3(new_n735), .A4(new_n671), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n673), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(G396));
  NOR2_X1   g0538(.A1(new_n432), .A2(new_n605), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n605), .A2(new_n416), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n427), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n739), .B1(new_n741), .B2(new_n432), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n643), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n742), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n664), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(new_n662), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n670), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n674), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n681), .A2(new_n674), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n253), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n717), .B1(G303), .B2(new_n700), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n237), .B2(new_n702), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n696), .A2(new_n388), .ZN(new_n755));
  INV_X1    g0555(.A(G311), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n691), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n348), .B1(new_n713), .B2(new_n239), .ZN(new_n758));
  NOR4_X1   g0558(.A1(new_n754), .A2(new_n755), .A3(new_n757), .A4(new_n758), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n759), .B1(new_n694), .B2(new_n684), .C1(new_n481), .C2(new_n706), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n696), .A2(new_n246), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n348), .B(new_n761), .C1(G50), .C2(new_n703), .ZN(new_n762));
  INV_X1    g0562(.A(G132), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n762), .B1(new_n362), .B2(new_n709), .C1(new_n763), .C2(new_n691), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT99), .ZN(new_n765));
  AOI22_X1  g0565(.A1(G143), .A2(new_n707), .B1(new_n714), .B2(G159), .ZN(new_n766));
  INV_X1    g0566(.A(G137), .ZN(new_n767));
  INV_X1    g0567(.A(G150), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n766), .B1(new_n767), .B2(new_n699), .C1(new_n768), .C2(new_n684), .ZN(new_n769));
  XOR2_X1   g0569(.A(new_n769), .B(KEYINPUT34), .Z(new_n770));
  OAI21_X1  g0570(.A(new_n760), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n681), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n749), .A2(new_n671), .A3(new_n752), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n748), .A2(new_n773), .ZN(G384));
  INV_X1    g0574(.A(KEYINPUT35), .ZN(new_n775));
  AOI211_X1 g0575(.A(new_n222), .B(new_n223), .C1(new_n526), .C2(new_n775), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n776), .B(G116), .C1(new_n775), .C2(new_n526), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT36), .ZN(new_n778));
  OAI21_X1  g0578(.A(G77), .B1(new_n362), .B2(new_n246), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n779), .A2(new_n221), .B1(G50), .B2(new_n246), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G1), .A3(new_n263), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT100), .Z(new_n783));
  INV_X1    g0583(.A(new_n405), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n589), .B2(new_n590), .ZN(new_n785));
  INV_X1    g0585(.A(new_n603), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n402), .B2(new_n397), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n399), .A2(new_n409), .A3(new_n787), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT37), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT37), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n399), .A2(new_n792), .A3(new_n409), .A4(new_n787), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(KEYINPUT38), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n377), .A2(new_n379), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n375), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n397), .B1(new_n382), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n786), .B(new_n799), .C1(new_n410), .C2(new_n405), .ZN(new_n800));
  INV_X1    g0600(.A(new_n399), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n406), .A2(new_n408), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n798), .B1(new_n802), .B2(new_n603), .ZN(new_n803));
  OAI21_X1  g0603(.A(KEYINPUT37), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n793), .ZN(new_n805));
  AND3_X1   g0605(.A1(new_n800), .A2(KEYINPUT38), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n795), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT40), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n512), .A2(new_n570), .A3(new_n470), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n627), .ZN(new_n810));
  INV_X1    g0610(.A(new_n659), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n744), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n581), .A2(new_n605), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n585), .A2(new_n320), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(new_n585), .B2(new_n320), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n807), .A2(new_n808), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT102), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n818), .B(new_n812), .C1(new_n814), .C2(new_n815), .ZN(new_n819));
  AOI21_X1  g0619(.A(KEYINPUT38), .B1(new_n800), .B2(new_n805), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n806), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n314), .A2(new_n315), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n581), .B(new_n605), .C1(new_n823), .C2(new_n321), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n585), .A2(new_n320), .A3(new_n813), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n818), .B1(new_n826), .B2(new_n812), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n808), .B1(new_n822), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT103), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT103), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n830), .B(new_n808), .C1(new_n822), .C2(new_n827), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n817), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n433), .A2(new_n660), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n832), .B(new_n833), .Z(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(G330), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT39), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n795), .B2(new_n806), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n316), .A2(new_n627), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT101), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n806), .A2(new_n820), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n837), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n664), .A2(new_n744), .B1(new_n432), .B2(new_n605), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n821), .A2(new_n844), .A3(new_n826), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n591), .A2(new_n603), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n645), .A2(new_n665), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n572), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n594), .B2(new_n595), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n847), .B(new_n850), .Z(new_n851));
  XOR2_X1   g0651(.A(new_n835), .B(new_n851), .Z(new_n852));
  NOR2_X1   g0652(.A1(new_n597), .A2(new_n259), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n783), .B1(new_n852), .B2(new_n853), .ZN(G367));
  NOR2_X1   g0654(.A1(new_n699), .A2(new_n756), .ZN(new_n855));
  INV_X1    g0655(.A(new_n463), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n856), .A2(new_n706), .B1(new_n481), .B2(new_n684), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n855), .B(new_n857), .C1(G317), .C2(new_n692), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n723), .A2(G97), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G283), .A2(new_n714), .B1(new_n710), .B2(new_n420), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT109), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(KEYINPUT109), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n325), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n858), .A2(new_n859), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT46), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT110), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n865), .A2(KEYINPUT110), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n703), .A2(G116), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n703), .A2(G116), .A3(new_n866), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n696), .A2(new_n253), .ZN(new_n871));
  INV_X1    g0671(.A(G143), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n699), .A2(new_n872), .B1(new_n713), .B2(new_n333), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n702), .A2(new_n362), .B1(new_n691), .B2(new_n767), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n709), .A2(new_n246), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n348), .B1(new_n685), .B2(G159), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n876), .B(new_n877), .C1(new_n768), .C2(new_n706), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT47), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n681), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n627), .A2(new_n563), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(new_n576), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n569), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n676), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n729), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n734), .B1(new_n218), .B2(new_n413), .C1(new_n234), .C2(new_n886), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n881), .A2(new_n671), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT106), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n544), .A2(new_n627), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n529), .A2(new_n605), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n542), .A2(new_n544), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n632), .A2(new_n625), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT42), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n621), .A2(new_n544), .A3(new_n542), .A4(new_n891), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n896), .A2(KEYINPUT105), .A3(new_n544), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT105), .B1(new_n896), .B2(new_n544), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n897), .A2(new_n898), .A3(new_n605), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n889), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  AOI211_X1 g0701(.A(KEYINPUT106), .B(new_n899), .C1(new_n894), .C2(KEYINPUT42), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n883), .A2(new_n884), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT104), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n630), .A2(new_n631), .B1(new_n622), .B2(new_n624), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT42), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n893), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n903), .A2(KEYINPUT107), .A3(new_n906), .A4(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n908), .B1(new_n907), .B2(new_n893), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT106), .B1(new_n911), .B2(new_n899), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n895), .A2(new_n889), .A3(new_n900), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(new_n906), .A4(new_n909), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT107), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n903), .A2(new_n909), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n906), .B1(KEYINPUT43), .B2(new_n904), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n893), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n626), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(KEYINPUT108), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT108), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n910), .A2(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n923), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n927), .A2(new_n923), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n637), .B(KEYINPUT41), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n625), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n614), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n633), .A2(KEYINPUT45), .A3(new_n893), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT45), .B1(new_n633), .B2(new_n893), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n633), .A2(KEYINPUT44), .A3(new_n893), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT44), .B1(new_n633), .B2(new_n893), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n934), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n937), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n935), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n944), .A2(new_n626), .A3(new_n940), .A4(new_n939), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n933), .A2(new_n630), .A3(new_n631), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n632), .A2(new_n625), .ZN(new_n947));
  AND4_X1   g0747(.A1(G330), .A2(new_n613), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(G330), .A2(new_n613), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n666), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n932), .B1(new_n951), .B2(new_n667), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n669), .A2(G1), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n930), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n888), .B1(new_n929), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT111), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT111), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n957), .B(new_n888), .C1(new_n929), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n956), .A2(new_n958), .ZN(G387));
  INV_X1    g0759(.A(new_n950), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n666), .B1(new_n948), .B2(new_n949), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n960), .A2(new_n637), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n948), .A2(new_n949), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n933), .A2(new_n676), .ZN(new_n964));
  INV_X1    g0764(.A(new_n681), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G322), .A2(new_n700), .B1(new_n685), .B2(G311), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n966), .B1(new_n686), .B2(new_n706), .C1(new_n856), .C2(new_n713), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT48), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n694), .B2(new_n709), .C1(new_n481), .C2(new_n702), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n325), .B1(new_n692), .B2(G326), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n239), .C2(new_n696), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n700), .A2(G159), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT113), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G77), .A2(new_n703), .B1(new_n685), .B2(new_n395), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n710), .A2(new_n565), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n246), .C2(new_n713), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n859), .B1(new_n768), .B2(new_n691), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n325), .B1(new_n706), .B2(new_n333), .ZN(new_n980));
  NOR4_X1   g0780(.A1(new_n975), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT114), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n965), .B1(new_n973), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n230), .A2(G45), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT112), .Z(new_n985));
  NOR2_X1   g0785(.A1(new_n336), .A2(G50), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT50), .ZN(new_n987));
  AOI21_X1  g0787(.A(G45), .B1(G68), .B2(G77), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n987), .A2(new_n639), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n729), .A3(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(G107), .B2(new_n218), .C1(new_n639), .C2(new_n732), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n670), .B(new_n983), .C1(new_n734), .C2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n963), .A2(new_n953), .B1(new_n964), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n962), .A2(new_n993), .ZN(G393));
  NAND2_X1  g0794(.A1(new_n942), .A2(new_n945), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n960), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n996), .A2(new_n637), .A3(new_n951), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n942), .A2(new_n945), .A3(new_n953), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n893), .A2(new_n677), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n734), .B1(new_n206), .B2(new_n218), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n240), .B2(new_n729), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n699), .A2(new_n768), .B1(new_n706), .B2(new_n720), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT51), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n325), .B1(new_n253), .B2(new_n709), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n702), .A2(new_n246), .B1(new_n713), .B2(new_n336), .ZN(new_n1005));
  NOR4_X1   g0805(.A1(new_n1003), .A2(new_n755), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n333), .B2(new_n684), .C1(new_n872), .C2(new_n691), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n699), .A2(new_n686), .B1(new_n706), .B2(new_n756), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT52), .Z(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n463), .B2(new_n685), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n714), .A2(G294), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n692), .A2(G322), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n702), .A2(new_n694), .B1(new_n696), .B2(new_n237), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n325), .B(new_n1013), .C1(G116), .C2(new_n710), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n965), .B1(new_n1007), .B2(new_n1015), .ZN(new_n1016));
  OR4_X1    g0816(.A1(new_n670), .A2(new_n999), .A3(new_n1001), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n997), .A2(new_n998), .A3(new_n1017), .ZN(G390));
  OAI221_X1 g0818(.A(new_n348), .B1(new_n709), .B2(new_n253), .C1(new_n481), .C2(new_n691), .ZN(new_n1019));
  AOI211_X1 g0819(.A(new_n761), .B(new_n1019), .C1(G87), .C2(new_n703), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G283), .A2(new_n700), .B1(new_n707), .B2(G116), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n420), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1022), .B1(new_n206), .B2(new_n713), .C1(new_n1023), .C2(new_n684), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n325), .B1(new_n684), .B2(new_n767), .C1(new_n763), .C2(new_n706), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n703), .A2(G150), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT53), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1025), .B(new_n1027), .C1(G159), .C2(new_n710), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G50), .A2(new_n723), .B1(new_n692), .B2(G125), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT54), .B(G143), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1028), .B(new_n1029), .C1(new_n713), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(G128), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n699), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n681), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n751), .A2(new_n336), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n671), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT117), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n837), .A2(new_n842), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n675), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g0843(.A1(new_n660), .A2(new_n661), .A3(new_n744), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n826), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n844), .A2(new_n826), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1047), .A2(new_n839), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n807), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n837), .A2(new_n842), .B1(new_n1047), .B2(new_n839), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n1045), .C1(new_n1040), .C2(new_n1048), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT116), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1044), .A2(new_n826), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n844), .B1(new_n1046), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1044), .A2(new_n826), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n844), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1059), .A2(new_n1060), .A3(new_n1045), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n833), .A2(G330), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n849), .B(new_n1063), .C1(new_n594), .C2(new_n595), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1056), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1064), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(KEYINPUT116), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1055), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n638), .B1(new_n1055), .B2(new_n1069), .ZN(new_n1071));
  AOI221_X4 g0871(.A(new_n1043), .B1(new_n953), .B2(new_n1055), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G378));
  XNOR2_X1  g0873(.A(new_n347), .B(KEYINPUT55), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n786), .A2(new_n339), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n1074), .B(new_n1075), .Z(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n674), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n751), .A2(new_n333), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G77), .A2(new_n703), .B1(new_n692), .B2(G283), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n362), .B2(new_n696), .C1(new_n413), .C2(new_n713), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n875), .B(new_n1083), .C1(G107), .C2(new_n707), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n206), .B2(new_n684), .C1(new_n239), .C2(new_n699), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n348), .A2(new_n287), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(new_n1087), .B(KEYINPUT118), .Z(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT58), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1086), .B(new_n333), .C1(G33), .C2(G41), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(KEYINPUT58), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n702), .A2(new_n1030), .B1(new_n709), .B2(new_n768), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n706), .A2(new_n1032), .B1(new_n713), .B2(new_n767), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1092), .B(new_n1093), .C1(G125), .C2(new_n700), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n763), .B2(new_n684), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT59), .Z(new_n1096));
  AOI211_X1 g0896(.A(G33), .B(G41), .C1(new_n692), .C2(G124), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n720), .C2(new_n696), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n681), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1080), .A2(new_n671), .A3(new_n1081), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n817), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n742), .B1(new_n646), .B2(new_n659), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n824), .B2(new_n825), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n841), .B1(new_n1105), .B2(new_n818), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n830), .B1(new_n1108), .B2(new_n808), .ZN(new_n1109));
  AOI211_X1 g0909(.A(KEYINPUT103), .B(KEYINPUT40), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1110));
  OAI211_X1 g0910(.A(G330), .B(new_n1103), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT120), .B1(new_n1111), .B2(new_n1079), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n661), .B(new_n817), .C1(new_n829), .C2(new_n831), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n847), .B1(new_n1113), .B2(new_n1078), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n847), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1111), .A2(new_n1115), .A3(new_n1079), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1111), .B2(new_n1079), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n832), .A2(G330), .A3(new_n847), .A4(new_n1078), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1078), .B1(new_n832), .B2(G330), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1119), .C1(KEYINPUT120), .C2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1102), .B1(new_n1122), .B2(new_n953), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1064), .B1(new_n1055), .B2(new_n1069), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(KEYINPUT57), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n637), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1124), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(KEYINPUT57), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1123), .B1(new_n1127), .B2(new_n1129), .ZN(G375));
  NAND2_X1  g0930(.A1(new_n1067), .A2(new_n953), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n824), .A2(new_n674), .A3(new_n825), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n699), .A2(new_n763), .B1(new_n684), .B2(new_n1030), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G137), .B2(new_n707), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT121), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n362), .A2(new_n696), .B1(new_n713), .B2(new_n768), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n348), .B(new_n1136), .C1(G128), .C2(new_n692), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n333), .C2(new_n709), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G159), .B2(new_n703), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1023), .A2(new_n713), .B1(new_n696), .B2(new_n253), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n977), .B1(new_n481), .B2(new_n699), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1140), .B(new_n1141), .C1(G303), .C2(new_n692), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n325), .B1(new_n703), .B2(G97), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1142), .B(new_n1143), .C1(new_n239), .C2(new_n684), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G283), .B2(new_n707), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n681), .B1(new_n1139), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n751), .A2(new_n246), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1132), .A2(new_n671), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1131), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n931), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1150), .B1(new_n1069), .B2(new_n1152), .ZN(G381));
  NAND2_X1  g0953(.A1(new_n1122), .A2(new_n953), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1101), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1128), .A2(KEYINPUT57), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n638), .B1(new_n1128), .B2(KEYINPUT57), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1072), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n1159), .A2(G384), .A3(G381), .ZN(new_n1160));
  INV_X1    g0960(.A(G390), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n956), .A2(new_n958), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(G393), .A2(G396), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1160), .A2(new_n1163), .A3(new_n1164), .ZN(G407));
  OAI211_X1 g0965(.A(G407), .B(G213), .C1(G343), .C2(new_n1159), .ZN(G409));
  INV_X1    g0966(.A(G213), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(G343), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1122), .A2(new_n931), .A3(new_n1125), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1123), .A2(new_n1072), .A3(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n1158), .C2(new_n1072), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1062), .A2(KEYINPUT60), .A3(new_n1064), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1065), .A2(new_n1068), .A3(KEYINPUT60), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n638), .B(new_n1174), .C1(new_n1175), .C2(new_n1151), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n748), .B(new_n773), .C1(new_n1176), .C2(new_n1149), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1174), .B1(new_n1175), .B2(new_n1151), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n637), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(G384), .A3(new_n1150), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1173), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(KEYINPUT62), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT61), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT122), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1177), .A2(new_n1180), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1185), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1168), .A2(G2897), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1186), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1185), .B(new_n1188), .C1(new_n1177), .C2(new_n1180), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1172), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT62), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1173), .A2(new_n1194), .A3(new_n1181), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1183), .A2(new_n1184), .A3(new_n1193), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n955), .A2(G390), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1161), .B(new_n888), .C1(new_n929), .C2(new_n954), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n737), .B1(new_n962), .B2(new_n993), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1164), .A2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1162), .A2(new_n1197), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1200), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1196), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(KEYINPUT123), .B1(new_n1204), .B2(KEYINPUT61), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT123), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1200), .B1(new_n1162), .B2(new_n1197), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1184), .C1(new_n1208), .C2(new_n1201), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1206), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1193), .A2(KEYINPUT63), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1182), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT124), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1173), .A2(new_n1213), .A3(KEYINPUT63), .A4(new_n1181), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1168), .B1(G375), .B2(G378), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1215), .A2(KEYINPUT63), .A3(new_n1181), .A4(new_n1171), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT124), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT125), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1212), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1212), .B2(new_n1218), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1205), .B1(new_n1220), .B2(new_n1221), .ZN(G405));
  NAND2_X1  g1022(.A1(G375), .A2(G378), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1159), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT126), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1181), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1224), .B(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(new_n1204), .ZN(G402));
endmodule


