//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G952), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n188), .B1(G234), .B2(G237), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI211_X1 g004(.A(new_n190), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT21), .B(G898), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(G475), .A2(G902), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n200), .A3(KEYINPUT88), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(KEYINPUT19), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n201), .A2(KEYINPUT19), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n197), .A3(G125), .ZN(new_n210));
  OAI211_X1 g024(.A(G146), .B(new_n210), .C1(new_n201), .C2(new_n209), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT90), .ZN(new_n212));
  NOR2_X1   g026(.A1(G237), .A2(G953), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(G143), .A3(G214), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(G143), .B1(new_n213), .B2(G214), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n212), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(G131), .B1(new_n215), .B2(new_n216), .ZN(new_n220));
  INV_X1    g034(.A(G237), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n187), .A3(G214), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n224), .A2(new_n212), .A3(new_n218), .A4(new_n214), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n208), .B(new_n211), .C1(new_n219), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n214), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT18), .A2(G131), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n203), .A2(G146), .A3(new_n204), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n198), .A2(new_n200), .A3(new_n206), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(new_n217), .B2(new_n229), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n228), .A2(KEYINPUT89), .A3(new_n230), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n231), .B(new_n234), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n227), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G113), .B(G122), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n210), .B1(new_n201), .B2(new_n209), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n206), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT17), .B(G131), .C1(new_n215), .C2(new_n216), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n246), .A2(new_n211), .A3(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT90), .B1(new_n228), .B2(G131), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT17), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n249), .A2(new_n250), .A3(new_n220), .A4(new_n225), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n242), .A3(new_n238), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n196), .B1(new_n244), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT91), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n252), .A2(new_n242), .A3(new_n238), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n242), .B1(new_n227), .B2(new_n238), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n195), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT20), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(new_n255), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n256), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n242), .B1(new_n252), .B2(new_n238), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n190), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G475), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT93), .B1(new_n269), .B2(G143), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n223), .A3(G128), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n223), .A2(G128), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT95), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n273), .A2(KEYINPUT95), .A3(new_n275), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G134), .ZN(new_n281));
  INV_X1    g095(.A(G122), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G116), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G122), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT92), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT92), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(G107), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G107), .ZN(new_n290));
  INV_X1    g104(.A(new_n288), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(new_n286), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n280), .A2(new_n281), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT13), .B1(new_n270), .B2(new_n272), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT94), .B1(new_n294), .B2(new_n274), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n270), .A2(new_n272), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT13), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n294), .A2(KEYINPUT94), .A3(new_n274), .ZN(new_n299));
  OAI21_X1  g113(.A(G134), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n285), .A2(KEYINPUT14), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n285), .A2(KEYINPUT14), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n283), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G107), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n278), .A2(G134), .A3(new_n279), .ZN(new_n306));
  AOI21_X1  g120(.A(G134), .B1(new_n278), .B2(new_n279), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n292), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT9), .B(G234), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(G217), .A3(new_n187), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n301), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n301), .B2(new_n308), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n190), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT96), .ZN(new_n316));
  INV_X1    g130(.A(G478), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(KEYINPUT15), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT96), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n319), .B(new_n190), .C1(new_n313), .C2(new_n314), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT97), .ZN(new_n322));
  OR2_X1    g136(.A1(new_n315), .A2(new_n318), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n321), .B2(new_n323), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n194), .B(new_n268), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G104), .B(G107), .ZN(new_n328));
  INV_X1    g142(.A(G101), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT80), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n290), .A2(G104), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n241), .A2(G107), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G101), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT81), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT1), .B1(new_n223), .B2(G146), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G128), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n206), .A2(G143), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n223), .A2(G146), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n340), .A2(new_n341), .A3(new_n344), .A4(G128), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n241), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n290), .A3(G104), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n347), .A2(new_n349), .A3(new_n329), .A4(new_n332), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n336), .A2(new_n337), .A3(new_n346), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n330), .A2(new_n335), .A3(new_n350), .ZN(new_n352));
  INV_X1    g166(.A(new_n345), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n338), .A2(G128), .B1(new_n340), .B2(new_n341), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT81), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n342), .A2(KEYINPUT0), .A3(G128), .ZN(new_n359));
  OR2_X1    g173(.A1(KEYINPUT0), .A2(G128), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT0), .A2(G128), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n340), .A2(new_n341), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n347), .A2(new_n349), .A3(new_n332), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G101), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n364), .A2(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n363), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n336), .A2(KEYINPUT10), .A3(new_n346), .A4(new_n350), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT11), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n281), .B2(G137), .ZN(new_n373));
  AOI21_X1  g187(.A(G131), .B1(new_n281), .B2(G137), .ZN(new_n374));
  INV_X1    g188(.A(G137), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT11), .A3(G134), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT65), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n373), .A2(new_n374), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n281), .A2(G137), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n373), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G131), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n371), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n378), .A2(new_n380), .B1(G131), .B2(new_n383), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n358), .A2(new_n387), .A3(new_n369), .A4(new_n370), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G110), .B(G140), .ZN(new_n390));
  INV_X1    g204(.A(G227), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G953), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n390), .B(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n352), .A2(new_n355), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n351), .A2(new_n356), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n385), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT12), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(KEYINPUT12), .A3(new_n385), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n394), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G469), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n190), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n403), .A2(new_n388), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n393), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n386), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(G469), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(G469), .A2(G902), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n414), .B(KEYINPUT87), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G113), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n284), .A2(G119), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G119), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G116), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n284), .A2(G119), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n417), .A2(KEYINPUT2), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G113), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(G116), .B(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n352), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n420), .A2(new_n424), .B1(new_n430), .B2(new_n429), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n434), .A2(new_n350), .A3(new_n335), .A4(new_n330), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(KEYINPUT8), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n359), .A2(G125), .A3(new_n360), .A4(new_n362), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n343), .A2(new_n199), .A3(new_n345), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n187), .A2(G224), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT84), .Z(new_n443));
  OR2_X1    g257(.A1(KEYINPUT85), .A2(KEYINPUT7), .ZN(new_n444));
  NAND2_X1  g258(.A1(KEYINPUT85), .A2(KEYINPUT7), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n436), .A2(new_n438), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT83), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n441), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n439), .A2(KEYINPUT83), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(KEYINPUT7), .A3(new_n443), .A4(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n447), .A2(new_n451), .A3(KEYINPUT86), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT86), .B1(new_n447), .B2(new_n451), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n422), .A2(new_n423), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(new_n426), .A3(new_n428), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n431), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n456), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n435), .A3(new_n437), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n452), .A2(new_n453), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n435), .ZN(new_n461));
  INV_X1    g275(.A(new_n437), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT6), .A3(new_n458), .ZN(new_n464));
  INV_X1    g278(.A(new_n443), .ZN(new_n465));
  INV_X1    g279(.A(new_n450), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT83), .B1(new_n439), .B2(new_n440), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n449), .A2(new_n443), .A3(new_n450), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n461), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n464), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n190), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n416), .B1(new_n460), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G214), .B1(G237), .B2(G902), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT82), .Z(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n447), .A2(new_n451), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n447), .A2(KEYINPUT86), .A3(new_n451), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n458), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n483), .A2(new_n190), .A3(new_n415), .A4(new_n473), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n475), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G221), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n310), .B2(new_n190), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n413), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n327), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT70), .ZN(new_n491));
  NOR2_X1   g305(.A1(G472), .A2(G902), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT31), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n385), .A2(new_n363), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n382), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n375), .A2(G134), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n281), .A2(KEYINPUT66), .A3(G137), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n378), .A2(new_n380), .B1(G131), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT68), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n346), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(G131), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n381), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(KEYINPUT30), .B(new_n495), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n381), .A2(new_n346), .A3(new_n504), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT64), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n362), .A2(new_n360), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n361), .B1(new_n340), .B2(new_n341), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n359), .A2(KEYINPUT64), .A3(new_n360), .A4(new_n362), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n507), .B1(new_n513), .B2(new_n387), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n456), .B(new_n506), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n456), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n520), .B(new_n495), .C1(new_n503), .C2(new_n505), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n213), .A2(G210), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n523), .B(KEYINPUT27), .Z(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G101), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n494), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n526), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n514), .A2(new_n456), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n521), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n529), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n519), .A2(new_n494), .A3(new_n527), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n493), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n491), .B1(new_n539), .B2(KEYINPUT32), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n519), .A2(new_n527), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT31), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n535), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n526), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n492), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT32), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(KEYINPUT70), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n495), .B1(new_n503), .B2(new_n505), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n456), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n534), .B1(new_n550), .B2(new_n521), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n521), .B2(new_n534), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n535), .A2(KEYINPUT71), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n529), .A2(KEYINPUT29), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n190), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n543), .A2(new_n526), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n529), .B1(new_n519), .B2(new_n521), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT29), .ZN(new_n562));
  OAI21_X1  g376(.A(G472), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n539), .A2(KEYINPUT32), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n540), .A2(new_n548), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT22), .B(G137), .ZN(new_n566));
  INV_X1    g380(.A(G234), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n486), .A2(new_n567), .A3(G953), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n566), .B(new_n568), .Z(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n269), .A2(G119), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n421), .A2(G128), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n246), .B2(new_n211), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(G110), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT72), .A4(KEYINPUT23), .ZN(new_n579));
  OR2_X1    g393(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n580));
  NAND2_X1  g394(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n580), .A2(G119), .A3(new_n269), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n578), .B1(new_n583), .B2(KEYINPUT73), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT73), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n579), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n584), .A2(KEYINPUT74), .A3(new_n586), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n577), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(KEYINPUT75), .B(G110), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n573), .A2(new_n574), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(new_n233), .A3(new_n211), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n570), .B1(new_n591), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n590), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT74), .B1(new_n584), .B2(new_n586), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n576), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n596), .A3(new_n569), .ZN(new_n602));
  OAI21_X1  g416(.A(G217), .B1(new_n567), .B2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n190), .ZN(new_n604));
  XOR2_X1   g418(.A(new_n604), .B(KEYINPUT77), .Z(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT78), .Z(new_n608));
  INV_X1    g422(.A(KEYINPUT76), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(KEYINPUT25), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n598), .A2(new_n602), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n610), .B1(new_n611), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n610), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n598), .A2(new_n602), .A3(new_n190), .A4(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n603), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n608), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n565), .A2(KEYINPUT79), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT79), .B1(new_n565), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n490), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT98), .B(G101), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G3));
  INV_X1    g436(.A(G472), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n623), .B1(new_n545), .B2(new_n190), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n624), .A2(new_n539), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n413), .A2(new_n488), .ZN(new_n626));
  INV_X1    g440(.A(new_n616), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n485), .A2(new_n194), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n316), .A2(new_n317), .A3(new_n320), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n317), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  INV_X1    g446(.A(new_n314), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n301), .A2(new_n308), .A3(new_n312), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT33), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n267), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n629), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n628), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n321), .A2(new_n323), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT97), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n324), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT99), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n266), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n265), .A2(KEYINPUT99), .A3(G475), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n263), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n646), .A2(new_n629), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n628), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n624), .A2(new_n539), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT100), .B1(new_n591), .B2(new_n597), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n601), .A2(new_n657), .A3(new_n596), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n570), .A2(KEYINPUT36), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n656), .A2(new_n658), .A3(new_n660), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n662), .A2(new_n606), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n615), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n490), .A2(new_n655), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT37), .B(G110), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT101), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n667), .B(new_n669), .ZN(G12));
  INV_X1    g484(.A(new_n626), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n565), .A2(new_n671), .A3(new_n666), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT102), .B(G900), .Z(new_n673));
  AOI21_X1  g487(.A(new_n189), .B1(new_n191), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  AND4_X1   g489(.A1(new_n263), .A2(new_n648), .A3(new_n649), .A4(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n645), .A2(new_n676), .A3(new_n485), .A4(new_n324), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT103), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n674), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n671), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n519), .A2(new_n521), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n529), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n550), .A2(new_n521), .ZN(new_n686));
  AOI21_X1  g500(.A(G902), .B1(new_n686), .B2(new_n526), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n623), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n539), .B2(KEYINPUT32), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n540), .A2(new_n689), .A3(new_n548), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n540), .A2(new_n689), .A3(new_n692), .A4(new_n548), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n646), .A2(new_n268), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n475), .A2(new_n484), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT38), .Z(new_n698));
  NAND4_X1  g512(.A1(new_n696), .A2(new_n698), .A3(new_n478), .A4(new_n665), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n683), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n223), .ZN(G45));
  NAND3_X1  g515(.A1(new_n638), .A2(new_n267), .A3(new_n675), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n489), .A2(new_n702), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n565), .A2(new_n703), .A3(new_n666), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n206), .ZN(G48));
  AOI22_X1  g519(.A1(new_n393), .A2(new_n389), .B1(new_n396), .B2(new_n403), .ZN(new_n706));
  OAI21_X1  g520(.A(G469), .B1(new_n706), .B2(G902), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n407), .A3(new_n488), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n565), .A2(new_n709), .A3(new_n616), .A4(new_n640), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND4_X1  g526(.A1(new_n651), .A2(new_n565), .A3(new_n709), .A4(new_n616), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NAND2_X1  g528(.A1(new_n709), .A2(new_n485), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n327), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n565), .A3(new_n666), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  AND4_X1   g532(.A1(new_n485), .A2(new_n645), .A3(new_n324), .A4(new_n267), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n529), .B1(new_n554), .B2(new_n556), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT105), .B1(new_n720), .B2(new_n528), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n551), .A2(new_n555), .A3(new_n553), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n722), .B(new_n542), .C1(new_n723), .C2(new_n529), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n721), .A2(new_n538), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n624), .B1(new_n725), .B2(new_n492), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n708), .A2(new_n193), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n719), .A2(new_n726), .A3(new_n616), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NAND3_X1  g543(.A1(new_n475), .A2(new_n484), .A3(new_n478), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n702), .A2(new_n708), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n726), .A2(new_n731), .A3(new_n666), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G125), .ZN(G27));
  AOI21_X1  g547(.A(KEYINPUT106), .B1(new_n697), .B2(new_n478), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  AOI211_X1 g549(.A(new_n735), .B(new_n477), .C1(new_n475), .C2(new_n484), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n626), .A2(new_n734), .A3(new_n702), .A4(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n564), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n546), .A2(new_n547), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n539), .A2(KEYINPUT107), .A3(KEYINPUT32), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n740), .A3(new_n563), .A4(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n737), .A2(KEYINPUT42), .A3(new_n742), .A4(new_n616), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n565), .A2(new_n616), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n626), .A2(new_n734), .A3(new_n736), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n744), .A2(new_n746), .A3(new_n702), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n743), .B1(new_n747), .B2(KEYINPUT42), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  NOR3_X1   g563(.A1(new_n646), .A2(new_n650), .A3(new_n674), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n745), .A3(new_n565), .A4(new_n616), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NOR2_X1   g566(.A1(new_n734), .A2(new_n736), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n630), .A2(new_n637), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n267), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n267), .B2(KEYINPUT109), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n756), .B(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n625), .A3(new_n666), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n754), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n409), .A2(new_n410), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n406), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n765), .B2(new_n764), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT46), .B1(new_n767), .B2(new_n412), .ZN(new_n768));
  INV_X1    g582(.A(new_n407), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(KEYINPUT46), .A3(new_n412), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n487), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n681), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n488), .ZN(new_n776));
  INV_X1    g590(.A(new_n681), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT108), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n763), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  XNOR2_X1  g594(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n772), .A2(new_n781), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n565), .A2(new_n754), .A3(new_n616), .A4(new_n702), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  AND2_X1   g601(.A1(new_n707), .A2(new_n407), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT49), .Z(new_n789));
  NOR3_X1   g603(.A1(new_n627), .A2(new_n477), .A3(new_n487), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n756), .B1(new_n790), .B2(KEYINPUT111), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n791), .B1(KEYINPUT111), .B2(new_n790), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n698), .B(new_n789), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n794), .B(new_n695), .C1(new_n793), .C2(new_n792), .ZN(new_n795));
  INV_X1    g609(.A(new_n644), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n639), .B1(new_n796), .B2(new_n267), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(new_n485), .A3(new_n194), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n628), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n667), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT79), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n744), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n617), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n800), .B1(new_n803), .B2(new_n490), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n710), .A2(new_n717), .A3(new_n713), .A4(new_n728), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n676), .A2(new_n796), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n806), .A2(new_n734), .A3(new_n736), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n565), .A3(new_n671), .A4(new_n666), .ZN(new_n808));
  INV_X1    g622(.A(new_n702), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n745), .A2(new_n666), .A3(new_n726), .A4(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n751), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n804), .A2(new_n748), .A3(new_n805), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n488), .A2(new_n413), .A3(new_n665), .A4(new_n675), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n719), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT70), .B1(new_n546), .B2(new_n547), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n491), .B(KEYINPUT32), .C1(new_n545), .C2(new_n492), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n692), .B1(new_n820), .B2(new_n689), .ZN(new_n821));
  INV_X1    g635(.A(new_n693), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n817), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n704), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT103), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n677), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n565), .A2(new_n671), .A3(new_n666), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n732), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n814), .B1(new_n825), .B2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n563), .A2(new_n564), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n665), .B1(new_n820), .B2(new_n831), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n694), .A2(new_n817), .B1(new_n832), .B2(new_n703), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n726), .A2(new_n731), .A3(new_n666), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n672), .B2(new_n678), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n833), .A2(KEYINPUT52), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n830), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n813), .A2(new_n837), .A3(KEYINPUT53), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n816), .B1(new_n691), .B2(new_n693), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n829), .A2(new_n840), .A3(new_n814), .A4(new_n704), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT52), .B1(new_n833), .B2(new_n835), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n839), .B1(new_n843), .B2(new_n812), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n748), .A2(new_n805), .A3(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n799), .A2(new_n667), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n811), .A2(new_n848), .A3(new_n620), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n804), .A2(KEYINPUT113), .A3(new_n811), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n837), .A2(new_n847), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n844), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n846), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n783), .A2(new_n784), .B1(new_n487), .B2(new_n788), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n759), .A2(new_n189), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n726), .A2(new_n616), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n753), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n695), .A2(new_n616), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n753), .A2(new_n709), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(KEYINPUT115), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(KEYINPUT115), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n189), .A3(new_n865), .ZN(new_n866));
  OR4_X1    g680(.A1(new_n267), .A2(new_n862), .A3(new_n638), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(new_n189), .A3(new_n759), .A4(new_n865), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n726), .A2(new_n666), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n861), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n698), .A2(new_n478), .A3(new_n708), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n858), .A2(new_n859), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT50), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n877), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT51), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n862), .A2(new_n639), .A3(new_n866), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n858), .A2(new_n859), .ZN(new_n882));
  OAI211_X1 g696(.A(G952), .B(new_n187), .C1(new_n882), .C2(new_n715), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n881), .A2(new_n883), .A3(KEYINPUT116), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT116), .B1(new_n881), .B2(new_n883), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n861), .A2(new_n867), .A3(new_n870), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n877), .A2(KEYINPUT51), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n742), .A2(new_n616), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n868), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT48), .B1(new_n891), .B2(KEYINPUT117), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT117), .B1(new_n868), .B2(new_n889), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n892), .B(new_n893), .Z(new_n894));
  NOR4_X1   g708(.A1(new_n856), .A2(new_n880), .A3(new_n888), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(G952), .A2(G953), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n795), .B1(new_n895), .B2(new_n896), .ZN(G75));
  AOI21_X1  g711(.A(new_n190), .B1(new_n844), .B2(new_n853), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n415), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n464), .A2(new_n472), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n470), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n903), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n187), .A2(G952), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(G51));
  XOR2_X1   g721(.A(new_n412), .B(KEYINPUT57), .Z(new_n908));
  AND3_X1   g722(.A1(new_n844), .A2(new_n853), .A3(new_n854), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n854), .B1(new_n844), .B2(new_n853), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(KEYINPUT118), .B(new_n908), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n405), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n898), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(new_n767), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n906), .B1(new_n915), .B2(new_n917), .ZN(G54));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  AOI211_X1 g733(.A(new_n919), .B(new_n916), .C1(new_n253), .C2(new_n244), .ZN(new_n920));
  INV_X1    g734(.A(new_n919), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n257), .B(new_n258), .C1(new_n898), .C2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n920), .A2(new_n906), .A3(new_n922), .ZN(G60));
  OR2_X1    g737(.A1(new_n635), .A2(new_n636), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT119), .ZN(new_n925));
  XNOR2_X1  g739(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n317), .A2(new_n190), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n925), .B(new_n928), .C1(new_n909), .C2(new_n910), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(G952), .B2(new_n187), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n925), .B1(new_n856), .B2(new_n928), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(new_n844), .A2(new_n853), .ZN(new_n933));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT121), .Z(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT60), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n906), .B1(new_n937), .B2(new_n611), .ZN(new_n938));
  INV_X1    g752(.A(new_n936), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n844), .B2(new_n853), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n662), .A2(new_n663), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n941), .B1(new_n940), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n938), .B(KEYINPUT61), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  AND2_X1   g763(.A1(new_n804), .A2(new_n805), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(G224), .A2(G953), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n952), .A2(G953), .B1(new_n192), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n901), .B1(G898), .B2(new_n187), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n954), .B(new_n956), .ZN(G69));
  NAND3_X1  g771(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n506), .B1(new_n517), .B2(new_n518), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT125), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n205), .A2(new_n207), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n803), .A2(new_n681), .A3(new_n745), .A4(new_n797), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n786), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n835), .A2(new_n824), .ZN(new_n965));
  OR3_X1    g779(.A1(new_n700), .A2(new_n965), .A3(KEYINPUT62), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT62), .B1(new_n700), .B2(new_n965), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n964), .A2(new_n966), .A3(new_n779), .A4(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n958), .B(new_n962), .C1(new_n968), .C2(G953), .ZN(new_n969));
  INV_X1    g783(.A(new_n965), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n779), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n786), .A2(new_n748), .A3(new_n751), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n742), .A2(new_n616), .A3(new_n719), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n778), .A2(new_n774), .A3(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n971), .A2(KEYINPUT126), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n779), .A2(new_n970), .A3(new_n975), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n972), .ZN(new_n979));
  AOI21_X1  g793(.A(G953), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n391), .A2(G900), .A3(G953), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n962), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n969), .B1(new_n980), .B2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n952), .B2(new_n968), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n685), .B1(new_n986), .B2(KEYINPUT127), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(KEYINPUT127), .B2(new_n986), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n684), .A2(new_n529), .ZN(new_n989));
  INV_X1    g803(.A(new_n952), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n976), .A2(new_n990), .A3(new_n979), .ZN(new_n991));
  INV_X1    g805(.A(new_n985), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n684), .A2(new_n526), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n992), .B1(new_n994), .B2(new_n541), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n906), .B1(new_n845), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n988), .A2(new_n993), .A3(new_n996), .ZN(G57));
endmodule


