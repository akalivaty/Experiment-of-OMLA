//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n773, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996;
  INV_X1    g000(.A(G120gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G113gat), .ZN(new_n203));
  INV_X1    g002(.A(G113gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G127gat), .ZN(new_n212));
  INV_X1    g011(.A(G127gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G134gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n209), .A2(new_n207), .ZN(new_n216));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n215), .B(new_n216), .C1(new_n217), .C2(KEYINPUT1), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT70), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n210), .A2(new_n218), .A3(KEYINPUT70), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224));
  INV_X1    g023(.A(G169gat), .ZN(new_n225));
  INV_X1    g024(.A(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n224), .B1(new_n227), .B2(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n227), .A2(KEYINPUT26), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT26), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n235), .A2(new_n225), .A3(new_n226), .A4(KEYINPUT68), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n228), .A2(new_n233), .A3(new_n234), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT27), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT27), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G183gat), .ZN(new_n241));
  INV_X1    g040(.A(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n243), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n239), .A2(new_n241), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n242), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n237), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(G183gat), .B2(G190gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  AND4_X1   g054(.A1(new_n250), .A2(new_n251), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(new_n225), .A3(new_n226), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n233), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT25), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n238), .A2(new_n242), .A3(KEYINPUT65), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(G183gat), .B2(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n255), .A2(KEYINPUT64), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n268), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n266), .A2(new_n254), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n259), .A2(new_n258), .B1(new_n231), .B2(new_n232), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n248), .A2(new_n262), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n223), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n251), .A3(new_n250), .A4(new_n255), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  AND3_X1   g076(.A1(new_n260), .A2(new_n233), .A3(new_n271), .ZN(new_n278));
  AOI22_X1  g077(.A1(KEYINPUT25), .A2(new_n277), .B1(new_n278), .B2(new_n270), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n279), .A2(new_n222), .A3(new_n221), .A4(new_n248), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT34), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT34), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n275), .A2(new_n280), .A3(new_n285), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G15gat), .B(G43gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(G71gat), .B(G99gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n281), .A2(new_n283), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT33), .B1(new_n281), .B2(new_n283), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n284), .B(new_n286), .C1(new_n295), .C2(new_n290), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(KEYINPUT32), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n300), .A3(new_n296), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT36), .B1(new_n302), .B2(KEYINPUT71), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n294), .A2(new_n300), .A3(new_n296), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n294), .B2(new_n296), .ZN(new_n305));
  OAI211_X1 g104(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT0), .ZN(new_n310));
  XNOR2_X1  g109(.A(G57gat), .B(G85gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  XOR2_X1   g111(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n313));
  INV_X1    g112(.A(KEYINPUT5), .ZN(new_n314));
  NAND2_X1  g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT2), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n319));
  AND2_X1   g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n315), .ZN(new_n324));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n325), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(new_n315), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT79), .B1(new_n324), .B2(new_n325), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n330), .A2(new_n331), .A3(new_n316), .A4(new_n322), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n219), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n327), .A2(new_n332), .A3(new_n210), .A4(new_n218), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n314), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n327), .A2(new_n332), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341));
  INV_X1    g140(.A(new_n219), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n340), .A2(KEYINPUT80), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT80), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n335), .B2(KEYINPUT4), .ZN(new_n345));
  INV_X1    g144(.A(new_n222), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT70), .B1(new_n210), .B2(new_n218), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n346), .A2(new_n333), .A3(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n343), .B(new_n345), .C1(new_n348), .C2(new_n341), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT81), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n342), .B1(new_n333), .B2(KEYINPUT3), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n327), .A2(new_n332), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n338), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n350), .B1(new_n349), .B2(new_n354), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n339), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n341), .B1(new_n223), .B2(new_n333), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n340), .A2(KEYINPUT4), .A3(new_n342), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n354), .A2(new_n358), .A3(new_n314), .A4(new_n359), .ZN(new_n360));
  AOI211_X1 g159(.A(new_n312), .B(new_n313), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n313), .ZN(new_n362));
  INV_X1    g161(.A(new_n360), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n349), .A2(new_n354), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT81), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n363), .B1(new_n367), .B2(new_n339), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n362), .B1(new_n368), .B2(new_n312), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n357), .A2(new_n360), .ZN(new_n370));
  INV_X1    g169(.A(new_n312), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n361), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n274), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n274), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(G211gat), .A2(G218gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(G211gat), .A2(G218gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT72), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G211gat), .ZN(new_n383));
  INV_X1    g182(.A(G218gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT72), .ZN(new_n386));
  NAND2_X1  g185(.A1(G211gat), .A2(G218gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(G197gat), .A2(G204gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(G197gat), .A2(G204gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT22), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(new_n387), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n393), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT73), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n393), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n377), .A2(new_n379), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(KEYINPUT75), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n376), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n274), .A2(KEYINPUT75), .A3(new_n375), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT74), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n279), .B2(new_n248), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(new_n375), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n274), .A2(new_n378), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n412), .A2(KEYINPUT74), .A3(new_n374), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n408), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n394), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n389), .A2(KEYINPUT73), .A3(new_n393), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT73), .B1(new_n389), .B2(new_n393), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n401), .B(new_n404), .C1(new_n414), .C2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT77), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n274), .A2(KEYINPUT75), .A3(new_n375), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT75), .B1(new_n274), .B2(new_n375), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n379), .A2(KEYINPUT74), .ZN(new_n425));
  AOI211_X1 g224(.A(new_n409), .B(new_n375), .C1(new_n274), .C2(new_n378), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n400), .B1(new_n427), .B2(new_n399), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT77), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n404), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n420), .A2(new_n421), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT76), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n404), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n411), .A2(new_n413), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n418), .B1(new_n435), .B2(new_n424), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT76), .B1(new_n436), .B2(new_n400), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n404), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n431), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n373), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G228gat), .ZN(new_n442));
  INV_X1    g241(.A(G233gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n416), .B2(new_n417), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n397), .A2(KEYINPUT84), .A3(new_n398), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n415), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n378), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n340), .B1(new_n450), .B2(new_n352), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n353), .A2(new_n378), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT85), .B1(new_n399), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n399), .A2(new_n452), .A3(KEYINPUT85), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n445), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT3), .B1(new_n418), .B2(new_n378), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n444), .B1(new_n458), .B2(new_n340), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n353), .A2(KEYINPUT86), .A3(new_n378), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT86), .B1(new_n353), .B2(new_n378), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n460), .A2(new_n461), .A3(new_n418), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G22gat), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT3), .B1(new_n449), .B2(new_n378), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n454), .B(new_n455), .C1(new_n467), .C2(new_n340), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n463), .B1(new_n468), .B2(new_n445), .ZN(new_n469));
  INV_X1    g268(.A(G22gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G50gat), .ZN(new_n474));
  XOR2_X1   g273(.A(G78gat), .B(G106gat), .Z(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n470), .B1(new_n457), .B2(new_n464), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT87), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n466), .A2(new_n471), .A3(new_n478), .A4(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n308), .B1(new_n441), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n370), .B2(new_n371), .ZN(new_n485));
  AOI211_X1 g284(.A(KEYINPUT89), .B(new_n312), .C1(new_n357), .C2(new_n360), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n357), .A2(new_n312), .A3(new_n360), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n313), .ZN(new_n488));
  NOR3_X1   g287(.A1(new_n485), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n404), .A2(KEYINPUT38), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n427), .A2(new_n418), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n377), .A2(new_n379), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(new_n399), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n490), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n428), .B2(new_n492), .ZN(new_n497));
  NOR4_X1   g296(.A1(new_n436), .A2(KEYINPUT90), .A3(KEYINPUT37), .A4(new_n400), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n339), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n365), .B2(new_n366), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n371), .B(new_n362), .C1(new_n501), .C2(new_n363), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n429), .B1(new_n428), .B2(new_n404), .ZN(new_n503));
  NOR4_X1   g302(.A1(new_n436), .A2(KEYINPUT77), .A3(new_n400), .A4(new_n434), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT91), .B1(new_n489), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n372), .A2(KEYINPUT89), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n370), .A2(new_n484), .A3(new_n371), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(new_n369), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n502), .A2(new_n420), .A3(new_n430), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n499), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n433), .A2(KEYINPUT37), .A3(new_n437), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n434), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n497), .A2(new_n498), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT38), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n507), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n481), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT87), .B1(new_n469), .B2(new_n470), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n520), .A2(new_n476), .B1(new_n466), .B2(new_n471), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n351), .A2(new_n353), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n358), .A3(new_n359), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(new_n338), .ZN(new_n525));
  OR2_X1    g324(.A1(new_n525), .A2(KEYINPUT39), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n525), .B(KEYINPUT39), .C1(new_n338), .C2(new_n336), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n312), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT40), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT88), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT88), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n526), .A2(new_n527), .A3(new_n312), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n438), .A2(new_n439), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n533), .B1(new_n534), .B2(new_n431), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n485), .A2(new_n486), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n522), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n483), .B1(new_n518), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n302), .B1(new_n480), .B2(new_n481), .ZN(new_n539));
  INV_X1    g338(.A(new_n440), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT35), .B1(new_n510), .B2(new_n502), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n368), .A2(new_n312), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n502), .B1(new_n544), .B2(new_n488), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n540), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n542), .A2(new_n543), .B1(new_n546), .B2(KEYINPUT35), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G113gat), .B(G141gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(G197gat), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT11), .B(G169gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT12), .Z(new_n553));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT16), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(G1gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n556), .B1(G1gat), .B2(new_n554), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G8gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n559));
  XNOR2_X1  g358(.A(G43gat), .B(G50gat), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(KEYINPUT92), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(KEYINPUT92), .B2(new_n560), .ZN(new_n562));
  OR3_X1    g361(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n563), .A2(new_n564), .B1(G29gat), .B2(G36gat), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n564), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(new_n570), .B2(new_n563), .ZN(new_n572));
  INV_X1    g371(.A(new_n560), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n573), .A2(new_n559), .B1(G29gat), .B2(G36gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n562), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n558), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n577), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT13), .Z(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n558), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT17), .B1(new_n568), .B2(new_n575), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(new_n585), .B2(KEYINPUT95), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n584), .A2(KEYINPUT95), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n575), .B(new_n568), .C1(new_n587), .C2(KEYINPUT17), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n583), .B1(KEYINPUT18), .B2(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n590), .A2(KEYINPUT18), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n553), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n590), .A2(KEYINPUT18), .ZN(new_n594));
  INV_X1    g393(.A(new_n553), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n590), .A2(KEYINPUT18), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n583), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n548), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G99gat), .B(G106gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n576), .B1(KEYINPUT17), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G190gat), .B(G218gat), .Z(new_n614));
  NOR3_X1   g413(.A1(new_n576), .A2(KEYINPUT17), .A3(new_n610), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G134gat), .B(G162gat), .Z(new_n619));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n619), .B(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n618), .A2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G64gat), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n627), .A2(G57gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(G57gat), .ZN(new_n629));
  AND2_X1   g428(.A1(G71gat), .A2(G78gat), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n628), .A2(new_n629), .B1(KEYINPUT9), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G71gat), .B(G78gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n558), .B1(KEYINPUT21), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT98), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT97), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n635), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n633), .A2(KEYINPUT21), .ZN(new_n641));
  XNOR2_X1  g440(.A(G127gat), .B(G155gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(G183gat), .B(G211gat), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n626), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(G230gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n443), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT100), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n633), .B1(new_n658), .B2(new_n609), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n610), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT10), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n610), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n660), .A2(new_n656), .A3(new_n443), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n655), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n664), .A2(new_n665), .A3(new_n655), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n651), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(KEYINPUT101), .A3(new_n666), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n650), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n600), .A2(new_n373), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g476(.A1(new_n600), .A2(new_n440), .A3(new_n675), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT16), .B(G8gat), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT102), .Z(new_n682));
  AOI22_X1  g481(.A1(new_n680), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(G1325gat));
  NAND2_X1  g483(.A1(new_n600), .A2(new_n675), .ZN(new_n685));
  OAI21_X1  g484(.A(G15gat), .B1(new_n685), .B2(new_n308), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n302), .A2(G15gat), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT103), .ZN(G1326gat));
  NOR2_X1   g488(.A1(new_n685), .A2(new_n482), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT43), .B(G22gat), .Z(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(G1327gat));
  OAI21_X1  g491(.A(new_n626), .B1(new_n538), .B2(new_n547), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n598), .A2(new_n649), .A3(new_n673), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(G29gat), .A3(new_n545), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT45), .Z(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n518), .A2(new_n537), .ZN(new_n701));
  INV_X1    g500(.A(new_n483), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n545), .A2(new_n431), .A3(new_n534), .ZN(new_n705));
  INV_X1    g504(.A(new_n302), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n519), .B2(new_n521), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT35), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n510), .A2(new_n502), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT35), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n709), .A2(new_n539), .A3(new_n710), .A4(new_n540), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n704), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n708), .A2(new_n711), .A3(new_n704), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n703), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n626), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  AOI22_X1  g517(.A1(new_n715), .A2(new_n718), .B1(new_n693), .B2(KEYINPUT44), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n700), .B1(new_n719), .B2(new_n695), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n708), .A2(new_n711), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n716), .B1(new_n722), .B2(new_n626), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n708), .A2(new_n704), .A3(new_n711), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n712), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n717), .B1(new_n725), .B2(new_n703), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT105), .B(new_n696), .C1(new_n723), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n728), .B2(new_n545), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n699), .A2(new_n729), .ZN(G1328gat));
  OAI21_X1  g529(.A(G36gat), .B1(new_n728), .B2(new_n540), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n697), .A2(G36gat), .A3(new_n540), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT46), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1329gat));
  NOR3_X1   g533(.A1(new_n724), .A2(new_n538), .A3(new_n712), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n694), .A2(new_n716), .B1(new_n735), .B2(new_n717), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n696), .ZN(new_n737));
  OAI211_X1 g536(.A(KEYINPUT47), .B(G43gat), .C1(new_n737), .C2(new_n308), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n697), .A2(G43gat), .A3(new_n302), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT47), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(KEYINPUT106), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n308), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n720), .A2(new_n743), .A3(new_n727), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n744), .A2(G43gat), .B1(new_n739), .B2(KEYINPUT106), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n745), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g545(.A(G50gat), .B1(new_n737), .B2(new_n482), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n482), .A2(G50gat), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n697), .A2(KEYINPUT108), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT108), .B1(new_n697), .B2(new_n749), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n747), .A2(KEYINPUT48), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n697), .A2(new_n749), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n720), .A2(new_n522), .A3(new_n727), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(G50gat), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT109), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n752), .B(new_n759), .C1(new_n755), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1331gat));
  AND4_X1   g560(.A1(new_n599), .A2(new_n715), .A3(new_n650), .A4(new_n672), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n373), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n440), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT49), .B(G64gat), .Z(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(G1333gat));
  NAND2_X1  g567(.A1(new_n762), .A2(new_n743), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n302), .A2(G71gat), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n769), .A2(G71gat), .B1(new_n762), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n762), .A2(new_n522), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g573(.A1(new_n598), .A2(new_n648), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n719), .A2(new_n673), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n373), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n605), .B1(new_n778), .B2(KEYINPUT110), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(KEYINPUT110), .B2(new_n778), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n781));
  INV_X1    g580(.A(new_n626), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n715), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n715), .A2(KEYINPUT111), .A3(KEYINPUT51), .A4(new_n783), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n786), .A2(new_n787), .B1(new_n785), .B2(new_n784), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n672), .A2(new_n605), .A3(new_n373), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n780), .B1(new_n788), .B2(new_n789), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n736), .A2(new_n672), .A3(new_n775), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n791), .B2(new_n540), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n672), .A2(new_n606), .A3(new_n440), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n792), .B(new_n793), .C1(new_n788), .C2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n786), .A2(new_n787), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT51), .B1(new_n784), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n715), .A2(KEYINPUT112), .A3(new_n783), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n794), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n606), .B1(new_n777), .B2(new_n440), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n796), .B(KEYINPUT52), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n787), .A2(new_n786), .B1(new_n799), .B2(new_n800), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n792), .B1(new_n806), .B2(new_n794), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n796), .B1(new_n807), .B2(KEYINPUT52), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n795), .B1(new_n805), .B2(new_n808), .ZN(G1337gat));
  OAI21_X1  g608(.A(G99gat), .B1(new_n791), .B2(new_n308), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n673), .A2(G99gat), .A3(new_n302), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n810), .B1(new_n788), .B2(new_n811), .ZN(G1338gat));
  OAI21_X1  g611(.A(G106gat), .B1(new_n791), .B2(new_n482), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n673), .A2(G106gat), .A3(new_n482), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n806), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT53), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n813), .B(new_n817), .C1(new_n788), .C2(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1339gat));
  INV_X1    g618(.A(new_n664), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n662), .A2(new_n657), .A3(new_n663), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  XOR2_X1   g621(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n823));
  AOI21_X1  g622(.A(new_n654), .B1(new_n664), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n670), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n598), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT115), .B1(new_n580), .B2(new_n582), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n581), .B2(new_n589), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n580), .A2(KEYINPUT115), .A3(new_n582), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n552), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n597), .A3(new_n672), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n626), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n626), .A2(new_n827), .A3(new_n829), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n597), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n649), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n675), .A2(new_n599), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n840), .A2(new_n844), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n522), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n440), .A2(new_n545), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n706), .A3(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(new_n204), .A3(new_n599), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n840), .A2(new_n844), .A3(new_n841), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n844), .B1(new_n840), .B2(new_n841), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n373), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n541), .ZN(new_n855));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n598), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n850), .A2(new_n856), .ZN(G1340gat));
  NOR3_X1   g656(.A1(new_n849), .A2(new_n202), .A3(new_n673), .ZN(new_n858));
  AOI21_X1  g657(.A(G120gat), .B1(new_n855), .B2(new_n672), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  OAI21_X1  g659(.A(G127gat), .B1(new_n849), .B2(new_n649), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n855), .A2(new_n213), .A3(new_n648), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1342gat));
  NAND3_X1  g662(.A1(new_n855), .A2(new_n211), .A3(new_n626), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n849), .B2(new_n782), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  XNOR2_X1  g667(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n825), .A2(new_n869), .ZN(new_n870));
  AOI211_X1 g669(.A(new_n870), .B(new_n828), .C1(new_n593), .C2(new_n597), .ZN(new_n871));
  AND3_X1   g670(.A1(new_n834), .A2(new_n597), .A3(new_n672), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT118), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n598), .A2(new_n829), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n874), .B(new_n835), .C1(new_n875), .C2(new_n870), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n873), .A2(new_n782), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n839), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n648), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n841), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n522), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n843), .A2(new_n883), .A3(new_n522), .A4(new_n845), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n308), .A2(new_n848), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G141gat), .B1(new_n886), .B2(new_n599), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n854), .A2(KEYINPUT119), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n853), .A2(new_n889), .A3(new_n373), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n743), .A2(new_n482), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n440), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n599), .A2(G141gat), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n888), .A2(new_n890), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n887), .A2(new_n898), .A3(new_n895), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1344gat));
  OAI211_X1 g699(.A(new_n883), .B(new_n522), .C1(new_n879), .C2(new_n880), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n851), .A2(new_n852), .A3(new_n482), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n883), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n672), .ZN(new_n904));
  OAI21_X1  g703(.A(G148gat), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT59), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n882), .A2(new_n672), .A3(new_n884), .A4(new_n885), .ZN(new_n907));
  INV_X1    g706(.A(G148gat), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(KEYINPUT59), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n907), .A2(KEYINPUT120), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT120), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n888), .A2(new_n890), .A3(new_n893), .ZN(new_n913));
  OR3_X1    g712(.A1(new_n913), .A2(G148gat), .A3(new_n673), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(G1345gat));
  OAI21_X1  g714(.A(G155gat), .B1(new_n886), .B2(new_n649), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n649), .A2(G155gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n913), .B2(new_n917), .ZN(G1346gat));
  INV_X1    g717(.A(G162gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n886), .A2(new_n919), .A3(new_n782), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n913), .A2(new_n782), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n540), .A2(new_n373), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n302), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n847), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n926), .A2(new_n225), .A3(new_n599), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n853), .A2(KEYINPUT121), .A3(new_n545), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n843), .A2(new_n545), .A3(new_n845), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT121), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n707), .A2(new_n540), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n598), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n927), .B1(new_n934), .B2(new_n225), .ZN(G1348gat));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n673), .A2(G176gat), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n853), .A2(new_n482), .A3(new_n925), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n226), .B1(new_n939), .B2(new_n672), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G176gat), .B1(new_n926), .B2(new_n673), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n932), .A2(new_n933), .ZN(new_n943));
  INV_X1    g742(.A(new_n937), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n942), .B(KEYINPUT122), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n945), .ZN(G1349gat));
  NAND2_X1  g745(.A1(new_n648), .A2(new_n245), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n932), .A2(new_n933), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n238), .B1(new_n939), .B2(new_n648), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT60), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G183gat), .B1(new_n926), .B2(new_n649), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT60), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n952), .B(new_n953), .C1(new_n943), .C2(new_n947), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n954), .ZN(G1350gat));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n626), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n956), .A2(new_n957), .A3(G190gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n956), .B2(G190gat), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n626), .A2(new_n242), .ZN(new_n961));
  OAI22_X1  g760(.A1(new_n959), .A2(new_n960), .B1(new_n943), .B2(new_n961), .ZN(G1351gat));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n903), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT57), .B1(new_n846), .B2(new_n482), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(KEYINPUT124), .A3(new_n901), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n924), .A2(new_n743), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n964), .A2(new_n966), .A3(new_n598), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G197gat), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n892), .A2(new_n540), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n971), .B1(new_n928), .B2(new_n931), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n599), .A2(G197gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT123), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n973), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(G1352gat));
  NAND4_X1  g775(.A1(new_n964), .A2(new_n966), .A3(new_n672), .A4(new_n967), .ZN(new_n977));
  XOR2_X1   g776(.A(KEYINPUT125), .B(G204gat), .Z(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n673), .A2(new_n978), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n972), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n972), .A2(new_n983), .A3(new_n980), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n979), .A2(new_n982), .A3(new_n984), .ZN(G1353gat));
  NAND4_X1  g784(.A1(new_n965), .A2(new_n648), .A3(new_n901), .A4(new_n967), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  INV_X1    g787(.A(KEYINPUT126), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n649), .A2(G211gat), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n972), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n989), .B1(new_n972), .B2(new_n990), .ZN(new_n992));
  OAI22_X1  g791(.A1(new_n987), .A2(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  AOI21_X1  g792(.A(G218gat), .B1(new_n972), .B2(new_n626), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n782), .A2(new_n384), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(G1355gat));
endmodule


