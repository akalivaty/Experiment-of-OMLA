

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759;

  XNOR2_X1 U371 ( .A(n495), .B(n496), .ZN(n735) );
  XNOR2_X1 U372 ( .A(G119), .B(n350), .ZN(n419) );
  BUF_X1 U373 ( .A(G128), .Z(n350) );
  BUF_X1 U374 ( .A(G107), .Z(n351) );
  XNOR2_X1 U375 ( .A(n481), .B(KEYINPUT4), .ZN(n499) );
  XNOR2_X1 U376 ( .A(n551), .B(n361), .ZN(n366) );
  XOR2_X2 U377 ( .A(KEYINPUT78), .B(KEYINPUT34), .Z(n362) );
  XNOR2_X2 U378 ( .A(n365), .B(n629), .ZN(n631) );
  XNOR2_X2 U379 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X2 U380 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X2 U381 ( .A(n462), .B(KEYINPUT90), .ZN(n711) );
  INV_X1 U382 ( .A(n351), .ZN(n440) );
  NAND2_X2 U383 ( .A1(n396), .A2(n393), .ZN(n513) );
  INV_X2 U384 ( .A(G953), .ZN(n748) );
  NOR2_X1 U385 ( .A1(n593), .A2(n592), .ZN(n677) );
  NAND2_X1 U386 ( .A1(n523), .A2(n412), .ZN(n585) );
  NAND2_X1 U387 ( .A1(n563), .A2(n523), .ZN(n712) );
  XNOR2_X1 U388 ( .A(n735), .B(n506), .ZN(n630) );
  AND2_X1 U389 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U390 ( .A(n540), .B(n539), .ZN(n553) );
  AND2_X1 U391 ( .A1(n405), .A2(n404), .ZN(n385) );
  XNOR2_X1 U392 ( .A(n584), .B(n583), .ZN(n598) );
  XNOR2_X1 U393 ( .A(n544), .B(KEYINPUT33), .ZN(n730) );
  XNOR2_X1 U394 ( .A(n465), .B(n464), .ZN(n580) );
  BUF_X1 U395 ( .A(n589), .Z(n590) );
  BUF_X1 U396 ( .A(n699), .Z(n386) );
  XNOR2_X1 U397 ( .A(n415), .B(G119), .ZN(n384) );
  BUF_X1 U398 ( .A(n367), .Z(n352) );
  XNOR2_X1 U399 ( .A(n527), .B(n399), .ZN(n367) );
  INV_X1 U400 ( .A(n526), .ZN(n353) );
  NAND2_X1 U401 ( .A1(n375), .A2(n378), .ZN(n374) );
  NAND2_X1 U402 ( .A1(n401), .A2(n376), .ZN(n375) );
  XNOR2_X1 U403 ( .A(n389), .B(n388), .ZN(n595) );
  INV_X1 U404 ( .A(KEYINPUT47), .ZN(n388) );
  NAND2_X1 U405 ( .A1(n373), .A2(n370), .ZN(n381) );
  AND2_X1 U406 ( .A1(n377), .A2(n374), .ZN(n373) );
  AND2_X1 U407 ( .A1(n401), .A2(n372), .ZN(n371) );
  XNOR2_X1 U408 ( .A(G902), .B(KEYINPUT15), .ZN(n507) );
  NAND2_X1 U409 ( .A1(n509), .A2(n610), .ZN(n397) );
  XNOR2_X1 U410 ( .A(G122), .B(G104), .ZN(n493) );
  XNOR2_X1 U411 ( .A(n423), .B(n422), .ZN(n484) );
  NAND2_X1 U412 ( .A1(n748), .A2(G234), .ZN(n423) );
  XOR2_X1 U413 ( .A(G137), .B(G140), .Z(n437) );
  XNOR2_X1 U414 ( .A(n502), .B(G104), .ZN(n439) );
  XNOR2_X1 U415 ( .A(G110), .B(KEYINPUT69), .ZN(n502) );
  XNOR2_X1 U416 ( .A(n491), .B(n490), .ZN(n523) );
  NOR2_X1 U417 ( .A1(n386), .A2(n391), .ZN(n586) );
  NAND2_X1 U418 ( .A1(n698), .A2(n354), .ZN(n391) );
  OR2_X1 U419 ( .A1(n637), .A2(G902), .ZN(n460) );
  XNOR2_X1 U420 ( .A(n746), .B(G146), .ZN(n459) );
  XNOR2_X1 U421 ( .A(G137), .B(G116), .ZN(n452) );
  XNOR2_X1 U422 ( .A(n481), .B(n482), .ZN(n414) );
  INV_X1 U423 ( .A(KEYINPUT40), .ZN(n406) );
  XNOR2_X1 U424 ( .A(n582), .B(n581), .ZN(n583) );
  INV_X1 U425 ( .A(KEYINPUT70), .ZN(n581) );
  INV_X1 U426 ( .A(KEYINPUT46), .ZN(n378) );
  NAND2_X1 U427 ( .A1(n677), .A2(n355), .ZN(n389) );
  INV_X1 U428 ( .A(KEYINPUT67), .ZN(n390) );
  NOR2_X1 U429 ( .A1(n759), .A2(n378), .ZN(n372) );
  NAND2_X1 U430 ( .A1(n379), .A2(n378), .ZN(n377) );
  INV_X1 U431 ( .A(n385), .ZN(n379) );
  XNOR2_X1 U432 ( .A(G131), .B(G140), .ZN(n469) );
  XNOR2_X1 U433 ( .A(G113), .B(G143), .ZN(n473) );
  XNOR2_X1 U434 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n497) );
  XNOR2_X1 U435 ( .A(KEYINPUT76), .B(KEYINPUT88), .ZN(n501) );
  XNOR2_X1 U436 ( .A(n387), .B(n597), .ZN(n616) );
  NAND2_X1 U437 ( .A1(n381), .A2(n380), .ZN(n387) );
  AND2_X1 U438 ( .A1(n689), .A2(n356), .ZN(n380) );
  NAND2_X1 U439 ( .A1(n395), .A2(n507), .ZN(n394) );
  XNOR2_X1 U440 ( .A(n433), .B(n432), .ZN(n699) );
  AND2_X1 U441 ( .A1(n699), .A2(n698), .ZN(n541) );
  AND2_X1 U442 ( .A1(n616), .A2(n614), .ZN(n369) );
  XNOR2_X1 U443 ( .A(n475), .B(n418), .ZN(n747) );
  XNOR2_X1 U444 ( .A(G137), .B(G140), .ZN(n418) );
  XOR2_X1 U445 ( .A(KEYINPUT65), .B(n611), .Z(n612) );
  XNOR2_X1 U446 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U447 ( .A(n602), .B(KEYINPUT106), .ZN(n411) );
  INV_X1 U448 ( .A(KEYINPUT86), .ZN(n409) );
  OR2_X1 U449 ( .A1(n463), .A2(n382), .ZN(n465) );
  XNOR2_X1 U450 ( .A(n383), .B(KEYINPUT30), .ZN(n382) );
  AND2_X1 U451 ( .A1(n586), .A2(n702), .ZN(n573) );
  INV_X1 U452 ( .A(KEYINPUT22), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n459), .B(n458), .ZN(n637) );
  XNOR2_X1 U454 ( .A(n369), .B(n750), .ZN(n749) );
  XNOR2_X1 U455 ( .A(n488), .B(n487), .ZN(n625) );
  XNOR2_X1 U456 ( .A(n414), .B(n413), .ZN(n488) );
  NAND2_X1 U457 ( .A1(n403), .A2(n402), .ZN(n401) );
  NAND2_X1 U458 ( .A1(n591), .A2(n601), .ZN(n689) );
  XNOR2_X1 U459 ( .A(n410), .B(n408), .ZN(n591) );
  XNOR2_X1 U460 ( .A(n409), .B(KEYINPUT36), .ZN(n408) );
  NAND2_X1 U461 ( .A1(n411), .A2(n590), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n585), .B(n534), .ZN(n676) );
  INV_X1 U463 ( .A(n386), .ZN(n572) );
  OR2_X1 U464 ( .A1(n451), .A2(n450), .ZN(n354) );
  AND2_X1 U465 ( .A1(n710), .A2(n390), .ZN(n355) );
  XOR2_X1 U466 ( .A(n596), .B(KEYINPUT72), .Z(n356) );
  AND2_X1 U467 ( .A1(n407), .A2(n541), .ZN(n357) );
  AND2_X1 U468 ( .A1(n537), .A2(n588), .ZN(n358) );
  AND2_X1 U469 ( .A1(n528), .A2(n588), .ZN(n359) );
  AND2_X1 U470 ( .A1(n529), .A2(n557), .ZN(n360) );
  XOR2_X1 U471 ( .A(n550), .B(KEYINPUT77), .Z(n361) );
  XOR2_X1 U472 ( .A(KEYINPUT66), .B(KEYINPUT19), .Z(n363) );
  INV_X1 U473 ( .A(G122), .ZN(n642) );
  BUF_X1 U474 ( .A(n521), .Z(n364) );
  BUF_X1 U475 ( .A(n630), .Z(n365) );
  NAND2_X1 U476 ( .A1(n554), .A2(n366), .ZN(n556) );
  XNOR2_X1 U477 ( .A(n366), .B(G122), .ZN(G24) );
  NAND2_X1 U478 ( .A1(n367), .A2(n358), .ZN(n540) );
  NAND2_X1 U479 ( .A1(n352), .A2(n360), .ZN(n552) );
  NAND2_X1 U480 ( .A1(n352), .A2(n359), .ZN(n566) );
  XNOR2_X1 U481 ( .A(n368), .B(n497), .ZN(n498) );
  XNOR2_X1 U482 ( .A(n368), .B(KEYINPUT10), .ZN(n475) );
  XNOR2_X2 U483 ( .A(G146), .B(G125), .ZN(n368) );
  NAND2_X1 U484 ( .A1(n620), .A2(n369), .ZN(n692) );
  NAND2_X1 U485 ( .A1(n609), .A2(n369), .ZN(n613) );
  XNOR2_X1 U486 ( .A(n499), .B(n436), .ZN(n746) );
  NAND2_X1 U487 ( .A1(n385), .A2(n401), .ZN(n758) );
  NAND2_X1 U488 ( .A1(n371), .A2(n385), .ZN(n370) );
  INV_X1 U489 ( .A(n759), .ZN(n376) );
  INV_X1 U490 ( .A(n702), .ZN(n557) );
  NAND2_X1 U491 ( .A1(n702), .A2(n711), .ZN(n383) );
  XNOR2_X2 U492 ( .A(n384), .B(n456), .ZN(n496) );
  XNOR2_X2 U493 ( .A(n446), .B(n445), .ZN(n574) );
  XNOR2_X2 U494 ( .A(n574), .B(KEYINPUT1), .ZN(n601) );
  XNOR2_X1 U495 ( .A(n400), .B(n492), .ZN(n494) );
  XNOR2_X2 U496 ( .A(G116), .B(G107), .ZN(n400) );
  NAND2_X1 U497 ( .A1(n521), .A2(n416), .ZN(n522) );
  XNOR2_X1 U498 ( .A(n589), .B(n363), .ZN(n521) );
  AND2_X1 U499 ( .A1(n392), .A2(n397), .ZN(n396) );
  NAND2_X1 U500 ( .A1(n630), .A2(n509), .ZN(n392) );
  OR2_X1 U501 ( .A1(n630), .A2(n394), .ZN(n393) );
  INV_X1 U502 ( .A(n509), .ZN(n395) );
  XNOR2_X2 U503 ( .A(n398), .B(KEYINPUT87), .ZN(n589) );
  NAND2_X1 U504 ( .A1(n513), .A2(n711), .ZN(n398) );
  XNOR2_X1 U505 ( .A(n400), .B(n483), .ZN(n413) );
  NAND2_X1 U506 ( .A1(n598), .A2(n406), .ZN(n405) );
  NOR2_X1 U507 ( .A1(n585), .A2(n406), .ZN(n402) );
  INV_X1 U508 ( .A(n598), .ZN(n403) );
  NAND2_X1 U509 ( .A1(n585), .A2(n406), .ZN(n404) );
  INV_X1 U510 ( .A(n541), .ZN(n695) );
  AND2_X1 U511 ( .A1(n574), .A2(n354), .ZN(n407) );
  INV_X1 U512 ( .A(n523), .ZN(n562) );
  NAND2_X1 U513 ( .A1(n676), .A2(n586), .ZN(n587) );
  INV_X1 U514 ( .A(n563), .ZN(n412) );
  XNOR2_X2 U515 ( .A(G113), .B(KEYINPUT3), .ZN(n415) );
  INV_X1 U516 ( .A(n364), .ZN(n592) );
  XNOR2_X1 U517 ( .A(n570), .B(KEYINPUT45), .ZN(n619) );
  XNOR2_X2 U518 ( .A(n624), .B(n623), .ZN(n657) );
  NAND2_X1 U519 ( .A1(n622), .A2(n694), .ZN(n624) );
  AND2_X1 U520 ( .A1(n520), .A2(n519), .ZN(n416) );
  XOR2_X1 U521 ( .A(n525), .B(KEYINPUT100), .Z(n417) );
  INV_X1 U522 ( .A(KEYINPUT8), .ZN(n422) );
  XNOR2_X1 U523 ( .A(n441), .B(n440), .ZN(n442) );
  INV_X1 U524 ( .A(KEYINPUT7), .ZN(n483) );
  INV_X1 U525 ( .A(KEYINPUT74), .ZN(n464) );
  XOR2_X1 U526 ( .A(KEYINPUT23), .B(G110), .Z(n420) );
  XNOR2_X1 U527 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U528 ( .A(n747), .B(n421), .ZN(n427) );
  XOR2_X1 U529 ( .A(KEYINPUT24), .B(KEYINPUT80), .Z(n425) );
  NAND2_X1 U530 ( .A1(G221), .A2(n484), .ZN(n424) );
  XOR2_X1 U531 ( .A(n425), .B(n424), .Z(n426) );
  XNOR2_X1 U532 ( .A(n427), .B(n426), .ZN(n653) );
  INV_X1 U533 ( .A(G902), .ZN(n489) );
  NAND2_X1 U534 ( .A1(n653), .A2(n489), .ZN(n433) );
  XOR2_X1 U535 ( .A(KEYINPUT93), .B(KEYINPUT25), .Z(n431) );
  NAND2_X1 U536 ( .A1(n507), .A2(G234), .ZN(n428) );
  XNOR2_X1 U537 ( .A(n428), .B(KEYINPUT92), .ZN(n429) );
  XNOR2_X1 U538 ( .A(KEYINPUT20), .B(n429), .ZN(n434) );
  NAND2_X1 U539 ( .A1(G217), .A2(n434), .ZN(n430) );
  XOR2_X1 U540 ( .A(n431), .B(n430), .Z(n432) );
  NAND2_X1 U541 ( .A1(n434), .A2(G221), .ZN(n435) );
  XOR2_X1 U542 ( .A(KEYINPUT21), .B(n435), .Z(n698) );
  XNOR2_X2 U543 ( .A(G143), .B(G128), .ZN(n481) );
  XNOR2_X1 U544 ( .A(G134), .B(G131), .ZN(n436) );
  XNOR2_X1 U545 ( .A(G101), .B(n437), .ZN(n438) );
  XNOR2_X1 U546 ( .A(n439), .B(n438), .ZN(n443) );
  NAND2_X1 U547 ( .A1(G227), .A2(n748), .ZN(n441) );
  XNOR2_X1 U548 ( .A(n459), .B(n444), .ZN(n658) );
  NOR2_X1 U549 ( .A1(n658), .A2(G902), .ZN(n446) );
  INV_X1 U550 ( .A(G469), .ZN(n445) );
  NAND2_X1 U551 ( .A1(G237), .A2(G234), .ZN(n447) );
  XNOR2_X1 U552 ( .A(n447), .B(KEYINPUT14), .ZN(n520) );
  INV_X1 U553 ( .A(n520), .ZN(n724) );
  NAND2_X1 U554 ( .A1(G953), .A2(G902), .ZN(n514) );
  NOR2_X1 U555 ( .A1(n724), .A2(n514), .ZN(n448) );
  XNOR2_X1 U556 ( .A(n448), .B(KEYINPUT103), .ZN(n449) );
  NOR2_X1 U557 ( .A1(G900), .A2(n449), .ZN(n451) );
  NAND2_X1 U558 ( .A1(n748), .A2(G952), .ZN(n518) );
  NOR2_X1 U559 ( .A1(n518), .A2(n724), .ZN(n450) );
  XNOR2_X1 U560 ( .A(KEYINPUT75), .B(n357), .ZN(n463) );
  XOR2_X1 U561 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n453) );
  XNOR2_X1 U562 ( .A(n453), .B(n452), .ZN(n455) );
  NOR2_X1 U563 ( .A1(G953), .A2(G237), .ZN(n466) );
  NAND2_X1 U564 ( .A1(n466), .A2(G210), .ZN(n454) );
  XNOR2_X1 U565 ( .A(n455), .B(n454), .ZN(n457) );
  XNOR2_X1 U566 ( .A(G101), .B(KEYINPUT68), .ZN(n456) );
  XNOR2_X1 U567 ( .A(n496), .B(n457), .ZN(n458) );
  XNOR2_X2 U568 ( .A(n460), .B(G472), .ZN(n702) );
  INV_X1 U569 ( .A(G237), .ZN(n461) );
  NAND2_X1 U570 ( .A1(n489), .A2(n461), .ZN(n508) );
  NAND2_X1 U571 ( .A1(n508), .A2(G214), .ZN(n462) );
  INV_X1 U572 ( .A(n711), .ZN(n604) );
  XNOR2_X1 U573 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n479) );
  XOR2_X1 U574 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n468) );
  NAND2_X1 U575 ( .A1(G214), .A2(n466), .ZN(n467) );
  XNOR2_X1 U576 ( .A(n468), .B(n467), .ZN(n472) );
  XOR2_X1 U577 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n470) );
  XNOR2_X1 U578 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U579 ( .A(n472), .B(n471), .ZN(n477) );
  XNOR2_X1 U580 ( .A(n493), .B(n473), .ZN(n474) );
  XNOR2_X1 U581 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U582 ( .A(n477), .B(n476), .ZN(n646) );
  NOR2_X1 U583 ( .A1(G902), .A2(n646), .ZN(n478) );
  XNOR2_X1 U584 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U585 ( .A(n480), .B(G475), .ZN(n563) );
  XNOR2_X1 U586 ( .A(n642), .B(G134), .ZN(n482) );
  XOR2_X1 U587 ( .A(KEYINPUT98), .B(KEYINPUT9), .Z(n486) );
  NAND2_X1 U588 ( .A1(G217), .A2(n484), .ZN(n485) );
  XNOR2_X1 U589 ( .A(n486), .B(n485), .ZN(n487) );
  NAND2_X1 U590 ( .A1(n625), .A2(n489), .ZN(n491) );
  INV_X1 U591 ( .A(G478), .ZN(n490) );
  NAND2_X1 U592 ( .A1(n412), .A2(n562), .ZN(n547) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U595 ( .A(n499), .B(n498), .ZN(n505) );
  NAND2_X1 U596 ( .A1(n748), .A2(G224), .ZN(n500) );
  XNOR2_X1 U597 ( .A(n501), .B(n500), .ZN(n503) );
  XNOR2_X1 U598 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U599 ( .A(n505), .B(n504), .ZN(n506) );
  INV_X1 U600 ( .A(n507), .ZN(n610) );
  AND2_X1 U601 ( .A1(n508), .A2(G210), .ZN(n509) );
  BUF_X1 U602 ( .A(n513), .Z(n510) );
  INV_X1 U603 ( .A(n510), .ZN(n511) );
  NOR2_X1 U604 ( .A1(n547), .A2(n511), .ZN(n512) );
  NAND2_X1 U605 ( .A1(n580), .A2(n512), .ZN(n594) );
  XNOR2_X1 U606 ( .A(n594), .B(G143), .ZN(G45) );
  INV_X1 U607 ( .A(G898), .ZN(n516) );
  INV_X1 U608 ( .A(n514), .ZN(n515) );
  NAND2_X1 U609 ( .A1(n516), .A2(n515), .ZN(n517) );
  NAND2_X1 U610 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X2 U611 ( .A(n522), .B(KEYINPUT0), .ZN(n559) );
  INV_X1 U612 ( .A(n559), .ZN(n526) );
  INV_X1 U613 ( .A(n698), .ZN(n524) );
  OR2_X1 U614 ( .A1(n712), .A2(n524), .ZN(n525) );
  NAND2_X1 U615 ( .A1(n526), .A2(n417), .ZN(n527) );
  NOR2_X1 U616 ( .A1(n601), .A2(n572), .ZN(n528) );
  XNOR2_X1 U617 ( .A(n702), .B(KEYINPUT6), .ZN(n588) );
  XNOR2_X1 U618 ( .A(n566), .B(G101), .ZN(G3) );
  NOR2_X1 U619 ( .A1(n601), .A2(n386), .ZN(n529) );
  XNOR2_X1 U620 ( .A(n552), .B(G110), .ZN(G12) );
  XNOR2_X1 U621 ( .A(n559), .B(KEYINPUT91), .ZN(n545) );
  INV_X1 U622 ( .A(n545), .ZN(n532) );
  AND2_X1 U623 ( .A1(n574), .A2(n541), .ZN(n530) );
  NAND2_X1 U624 ( .A1(n530), .A2(n557), .ZN(n531) );
  OR2_X1 U625 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U626 ( .A(n533), .B(KEYINPUT94), .ZN(n667) );
  INV_X1 U627 ( .A(KEYINPUT102), .ZN(n534) );
  INV_X1 U628 ( .A(n676), .ZN(n681) );
  NOR2_X1 U629 ( .A1(n667), .A2(n681), .ZN(n535) );
  XOR2_X1 U630 ( .A(G104), .B(n535), .Z(G6) );
  NAND2_X1 U631 ( .A1(n601), .A2(n572), .ZN(n536) );
  XNOR2_X1 U632 ( .A(n536), .B(KEYINPUT101), .ZN(n537) );
  INV_X1 U633 ( .A(KEYINPUT79), .ZN(n538) );
  XNOR2_X1 U634 ( .A(n538), .B(KEYINPUT32), .ZN(n539) );
  XNOR2_X1 U635 ( .A(n553), .B(G119), .ZN(G21) );
  NAND2_X1 U636 ( .A1(n601), .A2(n541), .ZN(n558) );
  INV_X1 U637 ( .A(n558), .ZN(n543) );
  INV_X1 U638 ( .A(n588), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U640 ( .A1(n545), .A2(n730), .ZN(n546) );
  XNOR2_X1 U641 ( .A(n546), .B(n362), .ZN(n549) );
  INV_X1 U642 ( .A(n547), .ZN(n548) );
  NAND2_X1 U643 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U644 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n550) );
  INV_X1 U645 ( .A(KEYINPUT44), .ZN(n555) );
  XNOR2_X1 U646 ( .A(n556), .B(n555), .ZN(n569) );
  OR2_X1 U647 ( .A1(n558), .A2(n557), .ZN(n705) );
  OR2_X1 U648 ( .A1(n353), .A2(n705), .ZN(n561) );
  INV_X1 U649 ( .A(KEYINPUT31), .ZN(n560) );
  XNOR2_X1 U650 ( .A(n561), .B(n560), .ZN(n684) );
  NAND2_X1 U651 ( .A1(n667), .A2(n684), .ZN(n565) );
  NAND2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n685) );
  INV_X1 U653 ( .A(KEYINPUT99), .ZN(n564) );
  XNOR2_X1 U654 ( .A(n685), .B(n564), .ZN(n599) );
  NAND2_X1 U655 ( .A1(n599), .A2(n585), .ZN(n710) );
  NAND2_X1 U656 ( .A1(n565), .A2(n710), .ZN(n567) );
  AND2_X1 U657 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U658 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U659 ( .A1(n619), .A2(n610), .ZN(n571) );
  XNOR2_X1 U660 ( .A(n571), .B(KEYINPUT81), .ZN(n609) );
  XNOR2_X1 U661 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n579) );
  XNOR2_X1 U662 ( .A(KEYINPUT28), .B(n573), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n575), .A2(n574), .ZN(n593) );
  INV_X1 U664 ( .A(n593), .ZN(n577) );
  NOR2_X1 U665 ( .A1(n712), .A2(n604), .ZN(n717) );
  XOR2_X1 U666 ( .A(KEYINPUT38), .B(n510), .Z(n714) );
  NAND2_X1 U667 ( .A1(n717), .A2(n714), .ZN(n576) );
  XNOR2_X1 U668 ( .A(n576), .B(KEYINPUT41), .ZN(n729) );
  NAND2_X1 U669 ( .A1(n577), .A2(n729), .ZN(n578) );
  XNOR2_X1 U670 ( .A(n579), .B(n578), .ZN(n759) );
  NAND2_X1 U671 ( .A1(n580), .A2(n714), .ZN(n584) );
  XOR2_X1 U672 ( .A(KEYINPUT85), .B(KEYINPUT39), .Z(n582) );
  NOR2_X1 U673 ( .A1(n588), .A2(n587), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  INV_X1 U675 ( .A(KEYINPUT48), .ZN(n597) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U677 ( .A(n600), .B(KEYINPUT107), .ZN(n756) );
  INV_X1 U678 ( .A(n756), .ZN(n608) );
  INV_X1 U679 ( .A(n601), .ZN(n696) );
  NAND2_X1 U680 ( .A1(n696), .A2(n602), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n605), .B(KEYINPUT43), .ZN(n606) );
  NOR2_X1 U683 ( .A1(n606), .A2(n510), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT104), .ZN(n757) );
  NOR2_X1 U685 ( .A1(n608), .A2(n757), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n610), .A2(KEYINPUT2), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n622) );
  AND2_X1 U688 ( .A1(n614), .A2(KEYINPUT2), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n618) );
  INV_X1 U690 ( .A(KEYINPUT82), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n618), .B(n617), .ZN(n621) );
  BUF_X1 U692 ( .A(n619), .Z(n620) );
  NAND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n694) );
  INV_X1 U694 ( .A(KEYINPUT64), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n657), .A2(G478), .ZN(n626) );
  XOR2_X1 U696 ( .A(n626), .B(n625), .Z(n628) );
  INV_X1 U697 ( .A(G952), .ZN(n627) );
  NAND2_X1 U698 ( .A1(n627), .A2(G953), .ZN(n649) );
  INV_X1 U699 ( .A(n649), .ZN(n665) );
  NOR2_X1 U700 ( .A1(n628), .A2(n665), .ZN(G63) );
  NAND2_X1 U701 ( .A1(n657), .A2(G210), .ZN(n632) );
  XNOR2_X1 U702 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n633), .A2(n649), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G51) );
  NAND2_X1 U707 ( .A1(n657), .A2(G472), .ZN(n639) );
  XOR2_X1 U708 ( .A(KEYINPUT108), .B(KEYINPUT62), .Z(n636) );
  XNOR2_X1 U709 ( .A(n639), .B(n638), .ZN(n640) );
  NAND2_X1 U710 ( .A1(n640), .A2(n649), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U712 ( .A1(n657), .A2(G475), .ZN(n648) );
  XNOR2_X1 U713 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n644) );
  XNOR2_X1 U714 ( .A(KEYINPUT59), .B(KEYINPUT89), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n648), .B(n647), .ZN(n650) );
  NAND2_X1 U717 ( .A1(n650), .A2(n649), .ZN(n652) );
  XOR2_X1 U718 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n651) );
  XNOR2_X1 U719 ( .A(n652), .B(n651), .ZN(G60) );
  NAND2_X1 U720 ( .A1(n657), .A2(G217), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n653), .B(KEYINPUT125), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X1 U723 ( .A1(n656), .A2(n665), .ZN(G66) );
  NAND2_X1 U724 ( .A1(n657), .A2(G469), .ZN(n664) );
  XNOR2_X1 U725 ( .A(n658), .B(KEYINPUT120), .ZN(n662) );
  XOR2_X1 U726 ( .A(KEYINPUT119), .B(KEYINPUT121), .Z(n660) );
  XNOR2_X1 U727 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n664), .B(n663), .ZN(n666) );
  NOR2_X1 U731 ( .A1(n666), .A2(n665), .ZN(G54) );
  NOR2_X1 U732 ( .A1(n667), .A2(n685), .ZN(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT110), .B(KEYINPUT27), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n669), .B(n668), .ZN(n670) );
  XOR2_X1 U735 ( .A(n670), .B(KEYINPUT26), .Z(n672) );
  XNOR2_X1 U736 ( .A(n351), .B(KEYINPUT109), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n672), .B(n671), .ZN(G9) );
  XOR2_X1 U738 ( .A(n350), .B(KEYINPUT29), .Z(n675) );
  INV_X1 U739 ( .A(n685), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n677), .A2(n673), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n675), .B(n674), .ZN(G30) );
  XOR2_X1 U742 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n679) );
  NAND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U744 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U745 ( .A(G146), .B(n680), .ZN(G48) );
  NOR2_X1 U746 ( .A1(n681), .A2(n684), .ZN(n683) );
  XNOR2_X1 U747 ( .A(G113), .B(KEYINPUT113), .ZN(n682) );
  XNOR2_X1 U748 ( .A(n683), .B(n682), .ZN(G15) );
  NOR2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  XOR2_X1 U750 ( .A(G116), .B(n686), .Z(G18) );
  XOR2_X1 U751 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n688) );
  XNOR2_X1 U752 ( .A(G125), .B(KEYINPUT37), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n688), .B(n687), .ZN(n690) );
  XOR2_X1 U754 ( .A(n690), .B(n689), .Z(G27) );
  INV_X1 U755 ( .A(KEYINPUT2), .ZN(n691) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  AND2_X1 U757 ( .A1(n694), .A2(n693), .ZN(n728) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U759 ( .A(n697), .B(KEYINPUT50), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n386), .A2(n698), .ZN(n700) );
  XOR2_X1 U761 ( .A(KEYINPUT49), .B(n700), .Z(n701) );
  NOR2_X1 U762 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U765 ( .A(KEYINPUT51), .B(n707), .Z(n708) );
  NAND2_X1 U766 ( .A1(n729), .A2(n708), .ZN(n709) );
  XNOR2_X1 U767 ( .A(n709), .B(KEYINPUT116), .ZN(n721) );
  NAND2_X1 U768 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n715) );
  AND2_X1 U770 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U772 ( .A(KEYINPUT117), .B(n718), .ZN(n719) );
  NAND2_X1 U773 ( .A1(n719), .A2(n730), .ZN(n720) );
  NAND2_X1 U774 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U775 ( .A(KEYINPUT52), .B(n722), .Z(n723) );
  NOR2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U777 ( .A1(n725), .A2(G952), .ZN(n726) );
  XOR2_X1 U778 ( .A(KEYINPUT118), .B(n726), .Z(n727) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U782 ( .A1(n733), .A2(G953), .ZN(n734) );
  XNOR2_X1 U783 ( .A(n734), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U784 ( .A(G110), .B(KEYINPUT127), .ZN(n736) );
  XNOR2_X1 U785 ( .A(n735), .B(n736), .ZN(n738) );
  NOR2_X1 U786 ( .A1(G898), .A2(n748), .ZN(n737) );
  NOR2_X1 U787 ( .A1(n738), .A2(n737), .ZN(n745) );
  NAND2_X1 U788 ( .A1(n620), .A2(n748), .ZN(n743) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n739) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n739), .ZN(n740) );
  NAND2_X1 U791 ( .A1(n740), .A2(G898), .ZN(n741) );
  XNOR2_X1 U792 ( .A(n741), .B(KEYINPUT126), .ZN(n742) );
  NAND2_X1 U793 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U794 ( .A(n745), .B(n744), .ZN(G69) );
  XNOR2_X1 U795 ( .A(n747), .B(n746), .ZN(n750) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n755) );
  INV_X1 U797 ( .A(n750), .ZN(n751) );
  XNOR2_X1 U798 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n753), .A2(G953), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n755), .A2(n754), .ZN(G72) );
  XNOR2_X1 U802 ( .A(G134), .B(n756), .ZN(G36) );
  XOR2_X1 U803 ( .A(G140), .B(n757), .Z(G42) );
  XOR2_X1 U804 ( .A(G131), .B(n758), .Z(G33) );
  XOR2_X1 U805 ( .A(G137), .B(n759), .Z(G39) );
endmodule

