//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT68), .ZN(new_n468));
  AOI22_X1  g043(.A1(G2105), .A2(new_n465), .B1(new_n468), .B2(G101), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(new_n459), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT67), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n466), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT70), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n480), .B(new_n481), .ZN(new_n482));
  OAI211_X1 g057(.A(G2105), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT69), .A3(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n475), .A2(G136), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n482), .A2(new_n485), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  AND4_X1   g068(.A1(new_n466), .A2(new_n493), .A3(new_n460), .A4(new_n462), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n470), .B1(new_n459), .B2(G2104), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(new_n460), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n496), .A2(G138), .A3(new_n466), .A4(new_n471), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n494), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n466), .A2(G114), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n483), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n498), .A2(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n504), .A2(new_n508), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(G166));
  AND2_X1   g088(.A1(new_n504), .A2(new_n508), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G89), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G651), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n518), .A2(new_n520), .A3(G51), .A4(G543), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT5), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G543), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n523), .A2(new_n525), .A3(G63), .A4(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n521), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n527), .B1(new_n521), .B2(new_n526), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n515), .B(new_n517), .C1(new_n528), .C2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(new_n504), .A2(G64), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n506), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n504), .A2(new_n508), .A3(G90), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n508), .A2(G52), .A3(G543), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(new_n523), .A2(new_n525), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  INV_X1    g115(.A(G68), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n522), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT72), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  OAI221_X1 g119(.A(new_n544), .B1(new_n541), .B2(new_n522), .C1(new_n539), .C2(new_n540), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(G651), .A3(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n508), .A2(G543), .ZN(new_n547));
  AOI22_X1  g122(.A1(G81), .A2(new_n514), .B1(new_n547), .B2(G43), .ZN(new_n548));
  AND2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND3_X1  g130(.A1(new_n504), .A2(new_n508), .A3(KEYINPUT73), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT73), .B1(new_n504), .B2(new_n508), .ZN(new_n558));
  OAI21_X1  g133(.A(G91), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n506), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n518), .A2(new_n520), .A3(G53), .A4(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n559), .A2(new_n561), .A3(new_n563), .ZN(G299));
  INV_X1    g139(.A(G171), .ZN(G301));
  OAI221_X1 g140(.A(new_n509), .B1(new_n510), .B2(new_n511), .C1(new_n505), .C2(new_n506), .ZN(G303));
  INV_X1    g141(.A(KEYINPUT73), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n510), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(new_n556), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n547), .A2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n569), .A2(G86), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n539), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(G651), .A2(new_n577), .B1(new_n547), .B2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G305));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n508), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n510), .A2(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n504), .A2(G60), .ZN(new_n584));
  NAND2_X1  g159(.A1(G72), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n506), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  OAI21_X1  g164(.A(G92), .B1(new_n557), .B2(new_n558), .ZN(new_n590));
  XNOR2_X1  g165(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n539), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(G651), .A2(new_n595), .B1(new_n547), .B2(G54), .ZN(new_n596));
  INV_X1    g171(.A(new_n591), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n569), .A2(G92), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n592), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n589), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n589), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g187(.A(new_n463), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n468), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT75), .B(KEYINPUT13), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n620));
  INV_X1    g195(.A(G135), .ZN(new_n621));
  INV_X1    g196(.A(G123), .ZN(new_n622));
  OAI221_X1 g197(.A(new_n620), .B1(new_n474), .B2(new_n621), .C1(new_n622), .C2(new_n483), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2427), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT15), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2435), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT77), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n634), .B(new_n637), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n630), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G14), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2084), .B(G2090), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n642), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT78), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n644), .A2(new_n645), .ZN(new_n651));
  AOI21_X1  g226(.A(KEYINPUT18), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n649), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n656), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT20), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n661), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n658), .A2(new_n660), .A3(new_n662), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n664), .C2(new_n663), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n669), .B(new_n674), .ZN(G229));
  XNOR2_X1  g250(.A(KEYINPUT85), .B(KEYINPUT36), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT34), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G22), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G166), .B2(new_n678), .ZN(new_n680));
  INV_X1    g255(.A(G1971), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n570), .A2(G16), .A3(new_n571), .A4(new_n572), .ZN(new_n683));
  OR2_X1    g258(.A1(G16), .A2(G23), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n685), .B1(new_n683), .B2(new_n684), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n678), .A2(G6), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G305), .B2(G16), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n677), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n692), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n691), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n686), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(new_n687), .ZN(new_n698));
  NAND4_X1  g273(.A1(new_n696), .A2(KEYINPUT34), .A3(new_n698), .A4(new_n682), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT81), .B(G29), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(G25), .ZN(new_n702));
  OR2_X1    g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n703), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n704));
  INV_X1    g279(.A(G131), .ZN(new_n705));
  INV_X1    g280(.A(G119), .ZN(new_n706));
  OAI221_X1 g281(.A(new_n704), .B1(new_n474), .B2(new_n705), .C1(new_n706), .C2(new_n483), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(KEYINPUT82), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n484), .A2(G119), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n475), .A2(G131), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .A4(new_n704), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n701), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n702), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n716), .B(new_n702), .C1(new_n713), .C2(new_n714), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G24), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n587), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT83), .B(G1986), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n722), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n720), .B(new_n724), .C1(new_n587), .C2(G16), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT84), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n676), .B1(new_n700), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n676), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n727), .B(new_n730), .C1(new_n694), .C2(new_n699), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n701), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n714), .A2(G35), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n733), .A2(new_n737), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G2090), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n678), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n678), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G1966), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(KEYINPUT93), .A3(G1966), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n701), .A2(G27), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n701), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(G2078), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n739), .B2(G2090), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n745), .A2(G1966), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT30), .B(G28), .Z(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n741), .A2(new_n750), .A3(new_n754), .A4(new_n759), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT24), .B(G34), .Z(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n701), .ZN(new_n762));
  AOI22_X1  g337(.A1(G160), .A2(G29), .B1(KEYINPUT89), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(KEYINPUT89), .B2(new_n762), .ZN(new_n764));
  INV_X1    g339(.A(G2084), .ZN(new_n765));
  NOR2_X1   g340(.A1(G5), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G171), .B2(G16), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(G1961), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n475), .A2(G140), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT86), .ZN(new_n771));
  INV_X1    g346(.A(G128), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n483), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT87), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n466), .A2(G116), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n771), .B(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G29), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n714), .A2(KEYINPUT28), .A3(G26), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(KEYINPUT28), .B1(new_n714), .B2(G26), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G2067), .Z(new_n783));
  NOR4_X1   g358(.A1(new_n732), .A2(new_n760), .A3(new_n769), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n549), .A2(new_n678), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n678), .B2(G19), .ZN(new_n786));
  INV_X1    g361(.A(G1341), .ZN(new_n787));
  OAI22_X1  g362(.A1(new_n786), .A2(new_n787), .B1(G1961), .B2(new_n767), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n787), .B2(new_n786), .ZN(new_n789));
  OR2_X1    g364(.A1(G29), .A2(G33), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n475), .A2(G139), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  AOI22_X1  g368(.A1(new_n613), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT88), .Z(new_n795));
  OAI211_X1 g370(.A(new_n791), .B(new_n793), .C1(new_n795), .C2(new_n466), .ZN(new_n796));
  INV_X1    g371(.A(G29), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n790), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G2072), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n678), .A2(KEYINPUT23), .A3(G20), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n802));
  INV_X1    g377(.A(G20), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G16), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n801), .B(new_n804), .C1(new_n604), .C2(new_n678), .ZN(new_n805));
  INV_X1    g380(.A(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n752), .A2(G2078), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n789), .A2(new_n800), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n678), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n600), .B2(new_n678), .ZN(new_n812));
  INV_X1    g387(.A(G1348), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n798), .A2(new_n799), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n784), .A2(new_n810), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n764), .A2(new_n765), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n623), .A2(new_n714), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n797), .A2(G32), .ZN(new_n819));
  AOI22_X1  g394(.A1(G129), .A2(new_n484), .B1(new_n475), .B2(G141), .ZN(new_n820));
  NAND3_X1  g395(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT90), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT26), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n468), .A2(G105), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n819), .B1(new_n825), .B2(new_n797), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT27), .B(G1996), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT91), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n826), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NOR4_X1   g405(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n830), .ZN(G311));
  INV_X1    g406(.A(new_n816), .ZN(new_n832));
  INV_X1    g407(.A(new_n817), .ZN(new_n833));
  INV_X1    g408(.A(new_n818), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n829), .ZN(G150));
  XNOR2_X1  g410(.A(KEYINPUT96), .B(G55), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n547), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n514), .A2(G93), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n523), .A2(new_n525), .A3(G67), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(KEYINPUT95), .B1(new_n841), .B2(G651), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT95), .ZN(new_n843));
  AOI211_X1 g418(.A(new_n843), .B(new_n506), .C1(new_n839), .C2(new_n840), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n837), .B(new_n838), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G860), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT37), .Z(new_n850));
  INV_X1    g425(.A(new_n549), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n846), .B2(new_n847), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n549), .A2(new_n845), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT39), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n600), .A2(G559), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT38), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n850), .B1(new_n858), .B2(G860), .ZN(G145));
  XOR2_X1   g434(.A(new_n477), .B(new_n623), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G162), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n777), .B(new_n713), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n796), .A2(G164), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n615), .B(KEYINPUT98), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n796), .A2(G164), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n869), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n871), .A2(new_n862), .A3(new_n867), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n484), .A2(G130), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n475), .A2(G142), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n466), .A2(G118), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n825), .B(new_n877), .ZN(new_n878));
  AND3_X1   g453(.A1(new_n870), .A2(new_n872), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n878), .B1(new_n870), .B2(new_n872), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n861), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n870), .A2(new_n872), .ZN(new_n882));
  INV_X1    g457(.A(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n870), .A2(new_n872), .A3(new_n878), .ZN(new_n885));
  INV_X1    g460(.A(new_n861), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT99), .B(G37), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n854), .B(new_n609), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n599), .A2(new_n604), .ZN(new_n894));
  NAND4_X1  g469(.A1(G299), .A2(new_n592), .A3(new_n596), .A4(new_n598), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT100), .B1(new_n894), .B2(new_n895), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n599), .B2(new_n604), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n896), .A2(new_n899), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n893), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n577), .A2(G651), .ZN(new_n910));
  INV_X1    g485(.A(G48), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n581), .ZN(new_n912));
  INV_X1    g487(.A(G86), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(new_n568), .B2(new_n556), .ZN(new_n914));
  OAI21_X1  g489(.A(G166), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n574), .A2(G303), .A3(new_n578), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n919));
  INV_X1    g494(.A(new_n586), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n514), .A2(G85), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n547), .A2(G47), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT101), .B1(new_n583), .B2(new_n586), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(G288), .A2(new_n925), .A3(new_n924), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n918), .A2(KEYINPUT102), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT102), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n917), .B(new_n930), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n927), .A2(new_n928), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT42), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n909), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n908), .A2(new_n934), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G868), .ZN(new_n939));
  INV_X1    g514(.A(G868), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n848), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n892), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n940), .B1(new_n936), .B2(new_n937), .ZN(new_n943));
  INV_X1    g518(.A(new_n941), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n943), .A2(KEYINPUT103), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n942), .A2(new_n945), .ZN(G295));
  NAND2_X1  g521(.A1(new_n939), .A2(new_n941), .ZN(G331));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(new_n534), .B2(new_n537), .ZN(new_n949));
  INV_X1    g524(.A(G64), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n533), .B1(new_n539), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(G651), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n952), .A2(KEYINPUT104), .A3(new_n536), .A4(new_n535), .ZN(new_n953));
  NAND3_X1  g528(.A1(G286), .A2(new_n949), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G286), .B1(new_n949), .B2(new_n953), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n852), .A2(new_n853), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n949), .A2(new_n953), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G168), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n954), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n843), .B1(new_n963), .B2(new_n506), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n841), .A2(KEYINPUT95), .A3(G651), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT97), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n837), .A4(new_n838), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n549), .B1(new_n962), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n549), .A2(new_n845), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n961), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n958), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n974), .B1(new_n896), .B2(new_n899), .ZN(new_n975));
  AOI211_X1 g550(.A(KEYINPUT106), .B(KEYINPUT41), .C1(new_n894), .C2(new_n895), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n896), .A2(new_n901), .ZN(new_n978));
  INV_X1    g553(.A(new_n902), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(KEYINPUT41), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n973), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n958), .A2(new_n896), .A3(new_n971), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n933), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT105), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n906), .B2(new_n972), .ZN(new_n985));
  INV_X1    g560(.A(new_n933), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n903), .A2(new_n905), .B1(new_n958), .B2(new_n971), .ZN(new_n988));
  NOR4_X1   g563(.A1(new_n988), .A2(new_n982), .A3(new_n933), .A4(KEYINPUT105), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n889), .B(new_n983), .C1(new_n987), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n958), .A2(new_n896), .A3(new_n971), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n978), .A2(new_n979), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n904), .B1(new_n995), .B2(new_n899), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n986), .B(new_n994), .C1(new_n996), .C2(new_n973), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT105), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n985), .A2(new_n984), .A3(new_n986), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G37), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n933), .B1(new_n988), .B2(new_n982), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1000), .A2(KEYINPUT43), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n992), .A2(new_n993), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1000), .A2(new_n991), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1006));
  AND4_X1   g581(.A1(KEYINPUT107), .A2(new_n1005), .A3(KEYINPUT44), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n993), .B1(new_n990), .B2(KEYINPUT43), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT107), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1004), .B1(new_n1007), .B2(new_n1009), .ZN(G397));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n498), .B2(new_n502), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n469), .A2(G40), .A3(new_n476), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT108), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n825), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT109), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n777), .B(G2067), .Z(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n1017), .B2(new_n825), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1016), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n713), .A2(new_n716), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n717), .B1(new_n708), .B2(new_n712), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1016), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1019), .A2(new_n1028), .A3(new_n825), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1021), .A2(new_n1024), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(new_n587), .B(G1986), .Z(new_n1031));
  AOI21_X1  g606(.A(new_n1030), .B1(new_n1016), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n1033));
  OAI211_X1 g608(.A(KEYINPUT45), .B(new_n1011), .C1(new_n498), .C2(new_n502), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n1014), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1012), .A2(KEYINPUT115), .A3(new_n1013), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(new_n1015), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1015), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1011), .C1(new_n498), .C2(new_n502), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  OAI22_X1  g619(.A1(new_n1039), .A2(G1966), .B1(G2084), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1033), .B(G8), .C1(new_n1045), .C2(G286), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G168), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1044), .A2(G2084), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1014), .A2(new_n1036), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1034), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1038), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n1041), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1966), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1050), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT51), .B(new_n1049), .C1(new_n1056), .C2(new_n1047), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT123), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1056), .A2(KEYINPUT123), .A3(new_n1049), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1046), .B(new_n1057), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1014), .A2(new_n1041), .A3(new_n1034), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n681), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT110), .B(G2090), .Z(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1044), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G8), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(G303), .A2(G8), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1068), .B(KEYINPUT55), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  XNOR2_X1  g646(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n1072));
  XOR2_X1   g647(.A(KEYINPUT112), .B(G1981), .Z(new_n1073));
  NOR2_X1   g648(.A1(G305), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1981), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n514), .A2(G86), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1075), .B1(new_n578), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1072), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(new_n1047), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT114), .B(new_n1072), .C1(new_n1074), .C2(new_n1077), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT111), .ZN(new_n1087));
  INV_X1    g662(.A(G1976), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1087), .B1(G288), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n919), .A2(KEYINPUT111), .A3(G1976), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1084), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT52), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(G288), .B2(new_n1088), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1084), .A2(new_n1089), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1086), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1071), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1044), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1040), .A2(KEYINPUT119), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1961), .ZN(new_n1103));
  OR2_X1    g678(.A1(new_n1062), .A2(G2078), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1102), .A2(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G2078), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1039), .A2(KEYINPUT53), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1108), .A3(G301), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(KEYINPUT53), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1041), .B2(KEYINPUT125), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1015), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1111), .A2(new_n1034), .A3(new_n1014), .A4(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1106), .A2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(KEYINPUT54), .B(new_n1109), .C1(new_n1115), .C2(G301), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1106), .A2(G301), .A3(new_n1114), .ZN(new_n1118));
  AOI21_X1  g693(.A(G301), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1061), .A2(new_n1098), .A3(new_n1116), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1102), .A2(new_n813), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1012), .A2(new_n1015), .A3(G2067), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1122), .A2(KEYINPUT120), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n1126));
  AOI21_X1  g701(.A(G1348), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1127), .B2(new_n1123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n599), .B1(new_n1129), .B2(KEYINPUT60), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT60), .ZN(new_n1131));
  AOI211_X1 g706(.A(new_n1131), .B(new_n600), .C1(new_n1125), .C2(new_n1128), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1130), .A2(new_n1132), .B1(KEYINPUT60), .B2(new_n1129), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT58), .B(G1341), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1062), .A2(G1996), .B1(new_n1083), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n549), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT59), .Z(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT56), .B(G2072), .Z(new_n1139));
  OR2_X1    g714(.A1(new_n1062), .A2(new_n1139), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1044), .A2(KEYINPUT117), .A3(new_n806), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT117), .B1(new_n1044), .B2(new_n806), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n559), .A2(new_n561), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT57), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(G299), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1147), .B(new_n1140), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT61), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1149), .A2(new_n1153), .A3(new_n1150), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1138), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1133), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1125), .A2(new_n600), .A3(new_n1128), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1149), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1159), .B2(new_n1150), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1150), .ZN(new_n1161));
  AOI211_X1 g736(.A(KEYINPUT121), .B(new_n1161), .C1(new_n1158), .C2(new_n1149), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1121), .B1(new_n1156), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1061), .A2(KEYINPUT62), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1045), .A2(new_n1058), .A3(new_n1048), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT123), .B1(new_n1056), .B2(new_n1049), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1168), .A2(new_n1169), .A3(new_n1046), .A4(new_n1057), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1165), .A2(new_n1119), .A3(new_n1098), .A4(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1095), .A2(new_n1070), .A3(new_n1067), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1074), .B1(new_n1173), .B2(new_n919), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1084), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT63), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1056), .A2(new_n1047), .A3(G286), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1097), .B2(new_n1179), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1070), .A2(KEYINPUT116), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1067), .A2(new_n1181), .ZN(new_n1182));
  AND4_X1   g757(.A1(KEYINPUT63), .A2(new_n1086), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1067), .A2(new_n1181), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1182), .A2(new_n1183), .A3(new_n1178), .A4(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1176), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1171), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1032), .B1(new_n1164), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1189));
  OR2_X1    g764(.A1(new_n1030), .A2(new_n1189), .ZN(new_n1190));
  NOR4_X1   g765(.A1(new_n1014), .A2(G1986), .A3(G290), .A4(new_n1015), .ZN(new_n1191));
  XOR2_X1   g766(.A(new_n1191), .B(KEYINPUT48), .Z(new_n1192));
  NAND2_X1  g767(.A1(new_n1030), .A2(new_n1189), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1022), .A2(new_n825), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1016), .ZN(new_n1196));
  NAND2_X1  g771(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1019), .A2(new_n1197), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1019), .A2(new_n1197), .ZN(new_n1199));
  OAI221_X1 g774(.A(new_n1196), .B1(KEYINPUT126), .B2(KEYINPUT46), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT47), .ZN(new_n1201));
  NAND4_X1  g776(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .A4(new_n1029), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(G2067), .B2(new_n777), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1203), .A2(new_n1016), .ZN(new_n1204));
  AND3_X1   g779(.A1(new_n1194), .A2(new_n1201), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1188), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(G227), .ZN(new_n1208));
  NAND3_X1  g782(.A1(new_n890), .A2(new_n640), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g783(.A(G229), .ZN(new_n1210));
  NAND4_X1  g784(.A1(new_n992), .A2(new_n1003), .A3(G319), .A4(new_n1210), .ZN(new_n1211));
  NOR2_X1   g785(.A1(new_n1209), .A2(new_n1211), .ZN(G308));
  OR2_X1    g786(.A1(new_n1209), .A2(new_n1211), .ZN(G225));
endmodule


