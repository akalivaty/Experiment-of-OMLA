

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588;

  INV_X1 U322 ( .A(n390), .ZN(n339) );
  XNOR2_X1 U323 ( .A(n340), .B(n339), .ZN(n352) );
  OR2_X1 U324 ( .A1(n578), .A2(KEYINPUT41), .ZN(n355) );
  XNOR2_X1 U325 ( .A(n352), .B(n351), .ZN(n354) );
  XNOR2_X1 U326 ( .A(n357), .B(KEYINPUT65), .ZN(n529) );
  XNOR2_X1 U327 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U328 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  INV_X1 U329 ( .A(KEYINPUT117), .ZN(n454) );
  XOR2_X1 U330 ( .A(G120GAT), .B(KEYINPUT0), .Z(n291) );
  XNOR2_X1 U331 ( .A(G113GAT), .B(G134GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n441) );
  XOR2_X1 U333 ( .A(G15GAT), .B(G127GAT), .Z(n319) );
  XOR2_X1 U334 ( .A(n441), .B(n319), .Z(n293) );
  NAND2_X1 U335 ( .A1(G227GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U336 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U337 ( .A(G71GAT), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U338 ( .A(KEYINPUT86), .B(KEYINPUT20), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U340 ( .A(n297), .B(n296), .Z(n306) );
  XNOR2_X1 U341 ( .A(KEYINPUT18), .B(KEYINPUT88), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n298), .B(KEYINPUT17), .ZN(n299) );
  XOR2_X1 U343 ( .A(n299), .B(KEYINPUT87), .Z(n301) );
  XNOR2_X1 U344 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n318) );
  XOR2_X1 U346 ( .A(G183GAT), .B(G99GAT), .Z(n303) );
  XNOR2_X1 U347 ( .A(G43GAT), .B(G190GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n318), .B(n304), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n527) );
  XOR2_X1 U351 ( .A(G36GAT), .B(G190GAT), .Z(n382) );
  XOR2_X1 U352 ( .A(KEYINPUT95), .B(n382), .Z(n308) );
  NAND2_X1 U353 ( .A1(G226GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n310) );
  XNOR2_X1 U355 ( .A(G8GAT), .B(G183GAT), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n309), .B(G211GAT), .ZN(n334) );
  XOR2_X1 U357 ( .A(n310), .B(n334), .Z(n316) );
  XOR2_X1 U358 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n312) );
  XNOR2_X1 U359 ( .A(G197GAT), .B(G218GAT), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n423) );
  XOR2_X1 U361 ( .A(G64GAT), .B(G92GAT), .Z(n314) );
  XNOR2_X1 U362 ( .A(G176GAT), .B(G204GAT), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n337) );
  XNOR2_X1 U364 ( .A(n423), .B(n337), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U366 ( .A(n318), .B(n317), .Z(n517) );
  XNOR2_X1 U367 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n409) );
  XOR2_X1 U368 ( .A(G22GAT), .B(G155GAT), .Z(n417) );
  XOR2_X1 U369 ( .A(G64GAT), .B(n417), .Z(n321) );
  XNOR2_X1 U370 ( .A(n319), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U372 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n323) );
  NAND2_X1 U373 ( .A1(G231GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U375 ( .A(n325), .B(n324), .Z(n327) );
  XOR2_X1 U376 ( .A(G1GAT), .B(KEYINPUT72), .Z(n367) );
  XNOR2_X1 U377 ( .A(n367), .B(KEYINPUT84), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n329) );
  XNOR2_X1 U380 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n331), .B(n330), .Z(n336) );
  XOR2_X1 U383 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n333) );
  XNOR2_X1 U384 ( .A(G71GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n338) );
  XNOR2_X1 U386 ( .A(n338), .B(n334), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n582) );
  XNOR2_X1 U388 ( .A(n582), .B(KEYINPUT107), .ZN(n558) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U390 ( .A(G99GAT), .B(G85GAT), .Z(n390) );
  XNOR2_X1 U391 ( .A(G106GAT), .B(G78GAT), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n341), .B(G148GAT), .ZN(n428) );
  INV_X1 U393 ( .A(KEYINPUT33), .ZN(n342) );
  NAND2_X1 U394 ( .A1(KEYINPUT74), .A2(n342), .ZN(n345) );
  INV_X1 U395 ( .A(KEYINPUT74), .ZN(n343) );
  NAND2_X1 U396 ( .A1(n343), .A2(KEYINPUT33), .ZN(n344) );
  NAND2_X1 U397 ( .A1(n345), .A2(n344), .ZN(n347) );
  XNOR2_X1 U398 ( .A(G120GAT), .B(KEYINPUT32), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n428), .B(n348), .ZN(n350) );
  XOR2_X1 U401 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n351) );
  NAND2_X1 U403 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n578) );
  NAND2_X1 U405 ( .A1(n578), .A2(KEYINPUT41), .ZN(n356) );
  NAND2_X1 U406 ( .A1(n356), .A2(n355), .ZN(n357) );
  XOR2_X1 U407 ( .A(G197GAT), .B(G22GAT), .Z(n359) );
  XNOR2_X1 U408 ( .A(G15GAT), .B(G141GAT), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U410 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n361) );
  XNOR2_X1 U411 ( .A(G8GAT), .B(KEYINPUT71), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U413 ( .A(n363), .B(n362), .ZN(n376) );
  XOR2_X1 U414 ( .A(G113GAT), .B(G50GAT), .Z(n365) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G36GAT), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U417 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U419 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U420 ( .A(n370), .B(KEYINPUT70), .Z(n374) );
  XOR2_X1 U421 ( .A(G29GAT), .B(G43GAT), .Z(n372) );
  XNOR2_X1 U422 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n371) );
  XNOR2_X1 U423 ( .A(n372), .B(n371), .ZN(n394) );
  XNOR2_X1 U424 ( .A(n394), .B(KEYINPUT69), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U426 ( .A(n376), .B(n375), .ZN(n573) );
  NAND2_X1 U427 ( .A1(n529), .A2(n573), .ZN(n378) );
  XNOR2_X1 U428 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n378), .B(n377), .ZN(n399) );
  XOR2_X1 U430 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n380) );
  XNOR2_X1 U431 ( .A(KEYINPUT77), .B(KEYINPUT10), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n386) );
  XNOR2_X1 U433 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n381) );
  XNOR2_X1 U434 ( .A(n381), .B(G162GAT), .ZN(n420) );
  XOR2_X1 U435 ( .A(n382), .B(n420), .Z(n384) );
  NAND2_X1 U436 ( .A1(G232GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n398) );
  XOR2_X1 U439 ( .A(KEYINPUT11), .B(G92GAT), .Z(n388) );
  XNOR2_X1 U440 ( .A(G106GAT), .B(G218GAT), .ZN(n387) );
  XNOR2_X1 U441 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U442 ( .A(n389), .B(KEYINPUT79), .Z(n392) );
  XNOR2_X1 U443 ( .A(G134GAT), .B(n390), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U445 ( .A(n393), .B(KEYINPUT78), .Z(n396) );
  XNOR2_X1 U446 ( .A(n394), .B(KEYINPUT80), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U448 ( .A(n398), .B(n397), .ZN(n553) );
  NAND2_X1 U449 ( .A1(n399), .A2(n553), .ZN(n400) );
  NOR2_X1 U450 ( .A1(n558), .A2(n400), .ZN(n401) );
  XNOR2_X1 U451 ( .A(n401), .B(KEYINPUT47), .ZN(n407) );
  XNOR2_X1 U452 ( .A(n553), .B(KEYINPUT36), .ZN(n584) );
  NOR2_X1 U453 ( .A1(n582), .A2(n584), .ZN(n403) );
  XNOR2_X1 U454 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n402) );
  XNOR2_X1 U455 ( .A(n403), .B(n402), .ZN(n405) );
  NOR2_X1 U456 ( .A1(n573), .A2(n578), .ZN(n404) );
  NAND2_X1 U457 ( .A1(n405), .A2(n404), .ZN(n406) );
  NAND2_X1 U458 ( .A1(n407), .A2(n406), .ZN(n408) );
  XOR2_X1 U459 ( .A(n409), .B(n408), .Z(n524) );
  NOR2_X1 U460 ( .A1(n517), .A2(n524), .ZN(n411) );
  XNOR2_X1 U461 ( .A(KEYINPUT54), .B(KEYINPUT116), .ZN(n410) );
  NAND2_X1 U462 ( .A1(n411), .A2(n410), .ZN(n413) );
  OR2_X1 U463 ( .A1(n411), .A2(n410), .ZN(n412) );
  NAND2_X1 U464 ( .A1(n413), .A2(n412), .ZN(n569) );
  XOR2_X1 U465 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n415) );
  XNOR2_X1 U466 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U468 ( .A(n416), .B(G204GAT), .Z(n419) );
  XNOR2_X1 U469 ( .A(n417), .B(G211GAT), .ZN(n418) );
  XNOR2_X1 U470 ( .A(n419), .B(n418), .ZN(n432) );
  XOR2_X1 U471 ( .A(n420), .B(KEYINPUT23), .Z(n422) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U473 ( .A(n422), .B(n421), .ZN(n424) );
  XOR2_X1 U474 ( .A(n424), .B(n423), .Z(n430) );
  XOR2_X1 U475 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n426) );
  XNOR2_X1 U476 ( .A(KEYINPUT3), .B(KEYINPUT92), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U478 ( .A(G141GAT), .B(n427), .Z(n445) );
  XNOR2_X1 U479 ( .A(n445), .B(n428), .ZN(n429) );
  XNOR2_X1 U480 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U481 ( .A(n432), .B(n431), .Z(n466) );
  XOR2_X1 U482 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n434) );
  XNOR2_X1 U483 ( .A(KEYINPUT1), .B(KEYINPUT94), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U485 ( .A(G85GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U486 ( .A(G29GAT), .B(G127GAT), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U488 ( .A(G57GAT), .B(G155GAT), .Z(n438) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(G148GAT), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U491 ( .A(n440), .B(n439), .Z(n447) );
  XOR2_X1 U492 ( .A(n441), .B(KEYINPUT5), .Z(n443) );
  NAND2_X1 U493 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U497 ( .A(n449), .B(n448), .ZN(n568) );
  INV_X1 U498 ( .A(n568), .ZN(n460) );
  NOR2_X1 U499 ( .A1(n466), .A2(n460), .ZN(n450) );
  AND2_X1 U500 ( .A1(n569), .A2(n450), .ZN(n451) );
  XNOR2_X1 U501 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NOR2_X1 U502 ( .A1(n527), .A2(n452), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n454), .B(n453), .ZN(n563) );
  NAND2_X1 U504 ( .A1(n563), .A2(n529), .ZN(n458) );
  XOR2_X1 U505 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n456) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT119), .Z(n455) );
  INV_X1 U507 ( .A(n573), .ZN(n543) );
  NOR2_X1 U508 ( .A1(n578), .A2(n543), .ZN(n491) );
  XNOR2_X1 U509 ( .A(n466), .B(KEYINPUT68), .ZN(n459) );
  XNOR2_X1 U510 ( .A(n459), .B(KEYINPUT28), .ZN(n485) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n517), .Z(n463) );
  NAND2_X1 U512 ( .A1(n460), .A2(n463), .ZN(n523) );
  NOR2_X1 U513 ( .A1(n485), .A2(n523), .ZN(n461) );
  NAND2_X1 U514 ( .A1(n527), .A2(n461), .ZN(n472) );
  NAND2_X1 U515 ( .A1(n466), .A2(n527), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT26), .ZN(n571) );
  INV_X1 U517 ( .A(n571), .ZN(n541) );
  AND2_X1 U518 ( .A1(n541), .A2(n463), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT96), .B(n464), .Z(n469) );
  NOR2_X1 U520 ( .A1(n527), .A2(n517), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT25), .B(n467), .ZN(n468) );
  NAND2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n568), .A2(n470), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n472), .A2(n471), .ZN(n488) );
  INV_X1 U526 ( .A(n553), .ZN(n562) );
  NOR2_X1 U527 ( .A1(n562), .A2(n582), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n473), .B(KEYINPUT16), .ZN(n474) );
  XOR2_X1 U529 ( .A(KEYINPUT85), .B(n474), .Z(n475) );
  AND2_X1 U530 ( .A1(n488), .A2(n475), .ZN(n502) );
  NAND2_X1 U531 ( .A1(n491), .A2(n502), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT97), .B(n476), .Z(n486) );
  NOR2_X1 U533 ( .A1(n568), .A2(n486), .ZN(n478) );
  XNOR2_X1 U534 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U536 ( .A(G1GAT), .B(n479), .Z(G1324GAT) );
  NOR2_X1 U537 ( .A1(n517), .A2(n486), .ZN(n481) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n527), .A2(n486), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n484), .ZN(G1326GAT) );
  INV_X1 U544 ( .A(n485), .ZN(n525) );
  NOR2_X1 U545 ( .A1(n525), .A2(n486), .ZN(n487) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  NAND2_X1 U547 ( .A1(n582), .A2(n488), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n584), .A2(n489), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT37), .B(n490), .Z(n514) );
  NAND2_X1 U550 ( .A1(n514), .A2(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(KEYINPUT38), .B(n492), .ZN(n499) );
  NOR2_X1 U552 ( .A1(n499), .A2(n568), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n493), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n517), .A2(n499), .ZN(n495) );
  XOR2_X1 U556 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  XNOR2_X1 U557 ( .A(KEYINPUT101), .B(KEYINPUT40), .ZN(n497) );
  NOR2_X1 U558 ( .A1(n527), .A2(n499), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(n498), .ZN(G1330GAT) );
  NOR2_X1 U561 ( .A1(n499), .A2(n525), .ZN(n500) );
  XOR2_X1 U562 ( .A(G50GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U563 ( .A(KEYINPUT102), .B(n501), .ZN(G1331GAT) );
  INV_X1 U564 ( .A(n529), .ZN(n545) );
  NOR2_X1 U565 ( .A1(n573), .A2(n545), .ZN(n513) );
  NAND2_X1 U566 ( .A1(n513), .A2(n502), .ZN(n503) );
  XOR2_X1 U567 ( .A(KEYINPUT103), .B(n503), .Z(n510) );
  NOR2_X1 U568 ( .A1(n568), .A2(n510), .ZN(n505) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n506), .Z(G1332GAT) );
  NOR2_X1 U572 ( .A1(n517), .A2(n510), .ZN(n507) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n527), .A2(n510), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(KEYINPUT105), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  NOR2_X1 U577 ( .A1(n525), .A2(n510), .ZN(n512) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n568), .A2(n520), .ZN(n515) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n515), .Z(n516) );
  XNOR2_X1 U583 ( .A(KEYINPUT106), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n520), .ZN(n518) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n527), .A2(n520), .ZN(n519) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n525), .A2(n520), .ZN(n521) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(n521), .Z(n522) );
  XNOR2_X1 U590 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n524), .A2(n523), .ZN(n542) );
  NAND2_X1 U592 ( .A1(n542), .A2(n525), .ZN(n526) );
  NOR2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n573), .A2(n537), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G113GAT), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT49), .B(KEYINPUT109), .Z(n531) );
  NAND2_X1 U597 ( .A1(n537), .A2(n529), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U599 ( .A(G120GAT), .B(n532), .Z(G1341GAT) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(KEYINPUT111), .ZN(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT110), .B(KEYINPUT50), .Z(n534) );
  NAND2_X1 U602 ( .A1(n537), .A2(n558), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT51), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U606 ( .A1(n537), .A2(n562), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n552) );
  NOR2_X1 U610 ( .A1(n543), .A2(n552), .ZN(n544) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n552), .ZN(n547) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n582), .A2(n552), .ZN(n550) );
  XNOR2_X1 U617 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(KEYINPUT115), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n573), .A2(n563), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n558), .A2(n563), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT121), .B(n561), .Z(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n577) );
  XOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .Z(n575) );
  NAND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(KEYINPUT122), .B(n572), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n573), .A2(n581), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(n577), .B(n576), .Z(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U644 ( .A1(n578), .A2(n581), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  INV_X1 U646 ( .A(n581), .ZN(n585) );
  OR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XOR2_X1 U652 ( .A(G218GAT), .B(n588), .Z(G1355GAT) );
endmodule

