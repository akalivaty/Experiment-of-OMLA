

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779;

  OR2_X1 U381 ( .A1(n748), .A2(G902), .ZN(n410) );
  NAND2_X1 U382 ( .A1(G214), .A2(n482), .ZN(n711) );
  XNOR2_X1 U383 ( .A(n495), .B(n494), .ZN(n743) );
  XNOR2_X1 U384 ( .A(G902), .B(KEYINPUT15), .ZN(n637) );
  AND2_X2 U385 ( .A1(n729), .A2(n426), .ZN(n392) );
  NAND2_X2 U386 ( .A1(n362), .A2(n447), .ZN(n614) );
  OR2_X2 U387 ( .A1(n695), .A2(n694), .ZN(n620) );
  NOR2_X2 U388 ( .A1(n694), .A2(n379), .ZN(n569) );
  AND2_X2 U389 ( .A1(n426), .A2(n443), .ZN(n400) );
  AND2_X2 U390 ( .A1(n380), .A2(n452), .ZN(n362) );
  XNOR2_X2 U391 ( .A(n389), .B(KEYINPUT78), .ZN(n735) );
  NAND2_X1 U392 ( .A1(n361), .A2(n393), .ZN(n390) );
  NAND2_X1 U393 ( .A1(n392), .A2(n375), .ZN(n361) );
  XNOR2_X2 U394 ( .A(n473), .B(G134), .ZN(n532) );
  NOR2_X1 U395 ( .A1(G953), .A2(G237), .ZN(n517) );
  XNOR2_X1 U396 ( .A(G119), .B(G128), .ZN(n500) );
  XNOR2_X1 U397 ( .A(G104), .B(G101), .ZN(n487) );
  INV_X1 U398 ( .A(G953), .ZN(n767) );
  NAND2_X1 U399 ( .A1(n558), .A2(n559), .ZN(n684) );
  AND2_X2 U400 ( .A1(n710), .A2(n438), .ZN(n416) );
  NOR2_X2 U401 ( .A1(n608), .A2(n594), .ZN(n595) );
  XNOR2_X2 U402 ( .A(n591), .B(KEYINPUT0), .ZN(n608) );
  NOR2_X1 U403 ( .A1(n624), .A2(n704), .ZN(n623) );
  INV_X1 U404 ( .A(n565), .ZN(n551) );
  INV_X2 U405 ( .A(G101), .ZN(n430) );
  AND2_X1 U406 ( .A1(n642), .A2(n691), .ZN(n729) );
  AND2_X1 U407 ( .A1(n602), .A2(n415), .ZN(n633) );
  NAND2_X1 U408 ( .A1(n566), .A2(n551), .ZN(n553) );
  BUF_X1 U409 ( .A(n544), .Z(n545) );
  XOR2_X1 U410 ( .A(G116), .B(G107), .Z(n529) );
  BUF_X1 U411 ( .A(n729), .Z(n363) );
  XNOR2_X1 U412 ( .A(n583), .B(KEYINPUT87), .ZN(n642) );
  NOR2_X1 U413 ( .A1(n567), .A2(n437), .ZN(n436) );
  XNOR2_X1 U414 ( .A(n465), .B(KEYINPUT30), .ZN(n567) );
  NAND2_X1 U415 ( .A1(n596), .A2(n711), .ZN(n465) );
  XNOR2_X1 U416 ( .A(n379), .B(KEYINPUT1), .ZN(n695) );
  NAND2_X2 U417 ( .A1(n407), .A2(n404), .ZN(n379) );
  XNOR2_X1 U418 ( .A(n527), .B(n526), .ZN(n566) );
  XNOR2_X1 U419 ( .A(n425), .B(n423), .ZN(n644) );
  XNOR2_X1 U420 ( .A(n531), .B(n533), .ZN(n425) );
  XNOR2_X1 U421 ( .A(n521), .B(n499), .ZN(n440) );
  XNOR2_X1 U422 ( .A(n424), .B(n529), .ZN(n423) );
  XNOR2_X1 U423 ( .A(n530), .B(G122), .ZN(n424) );
  XOR2_X1 U424 ( .A(G122), .B(G104), .Z(n523) );
  INV_X2 U425 ( .A(n414), .ZN(n581) );
  XNOR2_X2 U426 ( .A(n495), .B(n401), .ZN(n647) );
  XNOR2_X2 U427 ( .A(n753), .B(n481), .ZN(n665) );
  XNOR2_X2 U428 ( .A(n581), .B(KEYINPUT38), .ZN(n710) );
  AND2_X1 U429 ( .A1(n397), .A2(n671), .ZN(n634) );
  NAND2_X1 U430 ( .A1(n606), .A2(n605), .ZN(n635) );
  XNOR2_X1 U431 ( .A(n620), .B(n609), .ZN(n610) );
  XNOR2_X1 U432 ( .A(n497), .B(n498), .ZN(n521) );
  INV_X1 U433 ( .A(n568), .ZN(n438) );
  NOR2_X1 U434 ( .A1(G902), .A2(n657), .ZN(n527) );
  NAND2_X1 U435 ( .A1(n446), .A2(n444), .ZN(n443) );
  NAND2_X1 U436 ( .A1(n637), .A2(KEYINPUT66), .ZN(n446) );
  NAND2_X1 U437 ( .A1(n638), .A2(n445), .ZN(n444) );
  NAND2_X1 U438 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n445) );
  XNOR2_X1 U439 ( .A(G137), .B(G116), .ZN(n464) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n475) );
  XOR2_X1 U441 ( .A(KEYINPUT18), .B(KEYINPUT89), .Z(n476) );
  NAND2_X1 U442 ( .A1(n385), .A2(n381), .ZN(n636) );
  NAND2_X1 U443 ( .A1(n386), .A2(n411), .ZN(n385) );
  NAND2_X1 U444 ( .A1(n629), .A2(n612), .ZN(n451) );
  NAND2_X1 U445 ( .A1(n610), .A2(n612), .ZN(n452) );
  NOR2_X1 U446 ( .A1(n629), .A2(n421), .ZN(n577) );
  OR2_X1 U447 ( .A1(n687), .A2(n546), .ZN(n421) );
  NAND2_X1 U448 ( .A1(n449), .A2(n450), .ZN(n447) );
  NAND2_X1 U449 ( .A1(n496), .A2(G902), .ZN(n408) );
  XNOR2_X1 U450 ( .A(n522), .B(n441), .ZN(n657) );
  XNOR2_X1 U451 ( .A(n442), .B(n521), .ZN(n441) );
  INV_X1 U452 ( .A(KEYINPUT74), .ZN(n477) );
  INV_X1 U453 ( .A(KEYINPUT36), .ZN(n419) );
  NAND2_X1 U454 ( .A1(n365), .A2(n378), .ZN(n571) );
  INV_X1 U455 ( .A(n615), .ZN(n378) );
  NOR2_X1 U456 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U457 ( .A1(G953), .A2(G902), .ZN(n586) );
  AND2_X1 U458 ( .A1(n634), .A2(n607), .ZN(n387) );
  NAND2_X1 U459 ( .A1(n635), .A2(n634), .ZN(n411) );
  NAND2_X1 U460 ( .A1(n635), .A2(n607), .ZN(n383) );
  OR2_X1 U461 ( .A1(G237), .A2(G902), .ZN(n482) );
  XNOR2_X1 U462 ( .A(n524), .B(n525), .ZN(n442) );
  XNOR2_X1 U463 ( .A(G113), .B(G143), .ZN(n525) );
  NAND2_X1 U464 ( .A1(n443), .A2(n374), .ZN(n399) );
  NOR2_X1 U465 ( .A1(n566), .A2(n565), .ZN(n592) );
  AND2_X1 U466 ( .A1(n377), .A2(n369), .ZN(n568) );
  XNOR2_X1 U467 ( .A(n469), .B(KEYINPUT109), .ZN(n377) );
  XNOR2_X1 U468 ( .A(n402), .B(n367), .ZN(n401) );
  INV_X1 U469 ( .A(n440), .ZN(n766) );
  XOR2_X1 U470 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n530) );
  XNOR2_X1 U471 ( .A(KEYINPUT92), .B(G107), .ZN(n486) );
  XOR2_X1 U472 ( .A(KEYINPUT14), .B(n466), .Z(n723) );
  NAND2_X1 U473 ( .A1(G234), .A2(G237), .ZN(n466) );
  NAND2_X1 U474 ( .A1(n447), .A2(n372), .ZN(n718) );
  INV_X1 U475 ( .A(KEYINPUT34), .ZN(n613) );
  NAND2_X1 U476 ( .A1(n699), .A2(n698), .ZN(n694) );
  BUF_X1 U477 ( .A(n608), .Z(n624) );
  OR2_X1 U478 ( .A1(n743), .A2(n405), .ZN(n404) );
  AND2_X1 U479 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U480 ( .A1(G469), .A2(n406), .ZN(n405) );
  XNOR2_X1 U481 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U482 ( .A(n550), .B(KEYINPUT112), .ZN(n775) );
  NAND2_X1 U483 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n549) );
  XNOR2_X1 U485 ( .A(n553), .B(n422), .ZN(n687) );
  INV_X1 U486 ( .A(n571), .ZN(n683) );
  XNOR2_X1 U487 ( .A(n606), .B(G110), .ZN(G12) );
  XOR2_X1 U488 ( .A(n368), .B(n516), .Z(n364) );
  AND2_X1 U489 ( .A1(n570), .A2(n418), .ZN(n365) );
  XNOR2_X1 U490 ( .A(n512), .B(n511), .ZN(n366) );
  XOR2_X1 U491 ( .A(n463), .B(n462), .Z(n367) );
  XOR2_X1 U492 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n368) );
  OR2_X1 U493 ( .A1(n723), .A2(n470), .ZN(n369) );
  NOR2_X1 U494 ( .A1(n719), .A2(n718), .ZN(n370) );
  AND2_X1 U495 ( .A1(n642), .A2(n641), .ZN(n371) );
  AND2_X1 U496 ( .A1(n452), .A2(n451), .ZN(n372) );
  XNOR2_X1 U497 ( .A(G140), .B(G137), .ZN(n499) );
  INV_X1 U498 ( .A(G902), .ZN(n406) );
  XNOR2_X1 U499 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n373) );
  NAND2_X1 U500 ( .A1(n639), .A2(n731), .ZN(n374) );
  AND2_X1 U501 ( .A1(n638), .A2(KEYINPUT66), .ZN(n375) );
  BUF_X1 U502 ( .A(n663), .Z(n747) );
  NOR2_X2 U503 ( .A1(n778), .A2(n779), .ZN(n543) );
  NAND2_X1 U504 ( .A1(n376), .A2(n628), .ZN(n561) );
  INV_X1 U505 ( .A(n684), .ZN(n376) );
  NOR2_X1 U506 ( .A1(n567), .A2(n568), .ZN(n570) );
  XNOR2_X1 U507 ( .A(n595), .B(KEYINPUT22), .ZN(n602) );
  NAND2_X1 U508 ( .A1(n394), .A2(n399), .ZN(n393) );
  XNOR2_X1 U509 ( .A(n379), .B(KEYINPUT111), .ZN(n557) );
  NOR2_X1 U510 ( .A1(n625), .A2(n379), .ZN(n626) );
  AND2_X1 U511 ( .A1(n448), .A2(n451), .ZN(n380) );
  NAND2_X1 U512 ( .A1(n382), .A2(n619), .ZN(n381) );
  NAND2_X1 U513 ( .A1(n384), .A2(n383), .ZN(n382) );
  NOR2_X1 U514 ( .A1(n654), .A2(n412), .ZN(n384) );
  NAND2_X1 U515 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U516 ( .A1(n413), .A2(n412), .ZN(n388) );
  NAND2_X1 U517 ( .A1(n390), .A2(n735), .ZN(n643) );
  NAND2_X1 U518 ( .A1(n371), .A2(n426), .ZN(n389) );
  XNOR2_X2 U519 ( .A(n636), .B(n373), .ZN(n426) );
  NAND2_X1 U520 ( .A1(n400), .A2(n729), .ZN(n394) );
  NAND2_X1 U521 ( .A1(n395), .A2(n590), .ZN(n591) );
  AND2_X1 U522 ( .A1(n395), .A2(n557), .ZN(n559) );
  XNOR2_X1 U523 ( .A(n555), .B(n556), .ZN(n395) );
  XNOR2_X2 U524 ( .A(n396), .B(KEYINPUT16), .ZN(n427) );
  XNOR2_X1 U525 ( .A(n396), .B(n403), .ZN(n402) );
  XNOR2_X2 U526 ( .A(n429), .B(n428), .ZN(n396) );
  NAND2_X1 U527 ( .A1(n398), .A2(n628), .ZN(n397) );
  NAND2_X1 U528 ( .A1(n689), .A2(n675), .ZN(n398) );
  XNOR2_X1 U529 ( .A(n623), .B(n622), .ZN(n689) );
  NAND2_X1 U530 ( .A1(n647), .A2(n406), .ZN(n431) );
  XNOR2_X1 U531 ( .A(n464), .B(KEYINPUT77), .ZN(n403) );
  XNOR2_X2 U532 ( .A(n764), .B(G146), .ZN(n495) );
  XNOR2_X2 U533 ( .A(n532), .B(n457), .ZN(n764) );
  NAND2_X1 U534 ( .A1(n743), .A2(n496), .ZN(n409) );
  XNOR2_X2 U535 ( .A(n410), .B(n366), .ZN(n699) );
  INV_X1 U536 ( .A(KEYINPUT44), .ZN(n412) );
  INV_X1 U537 ( .A(n654), .ZN(n413) );
  NAND2_X1 U538 ( .A1(n414), .A2(n711), .ZN(n555) );
  XNOR2_X2 U539 ( .A(n485), .B(n453), .ZN(n414) );
  AND2_X1 U540 ( .A1(n414), .A2(n569), .ZN(n418) );
  XNOR2_X1 U541 ( .A(n474), .B(n497), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n535), .B(KEYINPUT40), .ZN(n778) );
  BUF_X1 U543 ( .A(n695), .Z(n415) );
  NAND2_X1 U544 ( .A1(n416), .A2(n569), .ZN(n437) );
  INV_X1 U545 ( .A(n539), .ZN(n596) );
  XNOR2_X1 U546 ( .A(n544), .B(KEYINPUT103), .ZN(n539) );
  NAND2_X1 U547 ( .A1(n577), .A2(n547), .ZN(n420) );
  NOR2_X1 U548 ( .A1(n585), .A2(n553), .ZN(n535) );
  XNOR2_X1 U549 ( .A(n417), .B(n433), .ZN(n432) );
  NAND2_X1 U550 ( .A1(n434), .A2(n435), .ZN(n417) );
  NAND2_X1 U551 ( .A1(n598), .A2(n597), .ZN(n606) );
  XNOR2_X2 U552 ( .A(n618), .B(n617), .ZN(n654) );
  XNOR2_X2 U553 ( .A(n427), .B(n471), .ZN(n753) );
  AND2_X1 U554 ( .A1(n576), .A2(n775), .ZN(n435) );
  INV_X1 U555 ( .A(KEYINPUT107), .ZN(n422) );
  INV_X1 U556 ( .A(n426), .ZN(n732) );
  OR2_X1 U557 ( .A1(n732), .A2(G953), .ZN(n756) );
  XNOR2_X2 U558 ( .A(KEYINPUT3), .B(G119), .ZN(n428) );
  XNOR2_X2 U559 ( .A(n430), .B(G113), .ZN(n429) );
  XNOR2_X2 U560 ( .A(n431), .B(G472), .ZN(n544) );
  NAND2_X1 U561 ( .A1(n432), .A2(n692), .ZN(n583) );
  INV_X1 U562 ( .A(KEYINPUT48), .ZN(n433) );
  XNOR2_X1 U563 ( .A(n543), .B(KEYINPUT46), .ZN(n434) );
  XNOR2_X1 U564 ( .A(n436), .B(KEYINPUT39), .ZN(n585) );
  XNOR2_X1 U565 ( .A(n439), .B(n440), .ZN(n748) );
  XNOR2_X1 U566 ( .A(n506), .B(n509), .ZN(n439) );
  XNOR2_X2 U567 ( .A(G143), .B(G128), .ZN(n473) );
  INV_X1 U568 ( .A(n608), .ZN(n448) );
  NOR2_X1 U569 ( .A1(n629), .A2(n612), .ZN(n449) );
  INV_X1 U570 ( .A(n610), .ZN(n450) );
  XNOR2_X1 U571 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X2 U572 ( .A(KEYINPUT100), .B(n554), .ZN(n628) );
  XOR2_X1 U573 ( .A(n484), .B(n483), .Z(n453) );
  AND2_X1 U574 ( .A1(n646), .A2(n651), .ZN(G63) );
  XNOR2_X1 U575 ( .A(KEYINPUT81), .B(n615), .ZN(n455) );
  NAND2_X1 U576 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U577 ( .A(KEYINPUT99), .ZN(n552) );
  AND2_X1 U578 ( .A1(n600), .A2(n629), .ZN(n601) );
  INV_X1 U579 ( .A(n752), .ZN(n651) );
  XNOR2_X1 U580 ( .A(KEYINPUT4), .B(G131), .ZN(n456) );
  XNOR2_X1 U581 ( .A(n456), .B(KEYINPUT72), .ZN(n457) );
  NAND2_X1 U582 ( .A1(n517), .A2(G210), .ZN(n463) );
  INV_X1 U583 ( .A(KEYINPUT95), .ZN(n458) );
  NAND2_X1 U584 ( .A1(KEYINPUT5), .A2(n458), .ZN(n461) );
  INV_X1 U585 ( .A(KEYINPUT5), .ZN(n459) );
  NAND2_X1 U586 ( .A1(n459), .A2(KEYINPUT95), .ZN(n460) );
  NAND2_X1 U587 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U588 ( .A1(n723), .A2(n586), .ZN(n467) );
  XOR2_X1 U589 ( .A(KEYINPUT108), .B(n467), .Z(n468) );
  NOR2_X1 U590 ( .A1(G900), .A2(n468), .ZN(n469) );
  INV_X1 U591 ( .A(G952), .ZN(n724) );
  NOR2_X1 U592 ( .A1(G953), .A2(n724), .ZN(n588) );
  INV_X1 U593 ( .A(n588), .ZN(n470) );
  XOR2_X1 U594 ( .A(n529), .B(n523), .Z(n471) );
  XNOR2_X1 U595 ( .A(G146), .B(G125), .ZN(n497) );
  NAND2_X1 U596 ( .A1(G224), .A2(n767), .ZN(n472) );
  XNOR2_X1 U597 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U598 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U599 ( .A(n477), .B(G110), .ZN(n491) );
  XNOR2_X1 U600 ( .A(n478), .B(n491), .ZN(n479) );
  XNOR2_X1 U601 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U602 ( .A1(n665), .A2(n637), .ZN(n485) );
  XOR2_X1 U603 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n484) );
  NAND2_X1 U604 ( .A1(G210), .A2(n482), .ZN(n483) );
  XNOR2_X1 U605 ( .A(n487), .B(n486), .ZN(n490) );
  NAND2_X1 U606 ( .A1(n767), .A2(G227), .ZN(n488) );
  XNOR2_X1 U607 ( .A(n488), .B(KEYINPUT80), .ZN(n489) );
  XNOR2_X1 U608 ( .A(n490), .B(n489), .ZN(n493) );
  XNOR2_X1 U609 ( .A(n491), .B(n499), .ZN(n492) );
  XNOR2_X1 U610 ( .A(n493), .B(n492), .ZN(n494) );
  INV_X1 U611 ( .A(G469), .ZN(n496) );
  XNOR2_X1 U612 ( .A(KEYINPUT71), .B(KEYINPUT10), .ZN(n498) );
  XOR2_X1 U613 ( .A(KEYINPUT79), .B(G110), .Z(n501) );
  XNOR2_X1 U614 ( .A(n501), .B(n500), .ZN(n505) );
  XOR2_X1 U615 ( .A(KEYINPUT24), .B(KEYINPUT73), .Z(n503) );
  XNOR2_X1 U616 ( .A(KEYINPUT93), .B(KEYINPUT23), .ZN(n502) );
  XNOR2_X1 U617 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U618 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U619 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n508) );
  NAND2_X1 U620 ( .A1(G234), .A2(n767), .ZN(n507) );
  XNOR2_X1 U621 ( .A(n508), .B(n507), .ZN(n528) );
  NAND2_X1 U622 ( .A1(G221), .A2(n528), .ZN(n509) );
  XOR2_X1 U623 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n512) );
  NAND2_X1 U624 ( .A1(G234), .A2(n637), .ZN(n510) );
  XNOR2_X1 U625 ( .A(KEYINPUT20), .B(n510), .ZN(n513) );
  NAND2_X1 U626 ( .A1(n513), .A2(G217), .ZN(n511) );
  NAND2_X1 U627 ( .A1(n513), .A2(G221), .ZN(n515) );
  INV_X1 U628 ( .A(KEYINPUT21), .ZN(n514) );
  XNOR2_X1 U629 ( .A(n515), .B(n514), .ZN(n698) );
  XNOR2_X1 U630 ( .A(G131), .B(G140), .ZN(n516) );
  XOR2_X1 U631 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n519) );
  NAND2_X1 U632 ( .A1(G214), .A2(n517), .ZN(n518) );
  XNOR2_X1 U633 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U634 ( .A(n364), .B(n520), .ZN(n522) );
  INV_X1 U635 ( .A(n523), .ZN(n524) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(G475), .ZN(n526) );
  NAND2_X1 U637 ( .A1(G217), .A2(n528), .ZN(n531) );
  INV_X1 U638 ( .A(n532), .ZN(n533) );
  NAND2_X1 U639 ( .A1(n644), .A2(n406), .ZN(n534) );
  XNOR2_X2 U640 ( .A(n534), .B(G478), .ZN(n565) );
  NAND2_X1 U641 ( .A1(n711), .A2(n710), .ZN(n715) );
  INV_X1 U642 ( .A(n592), .ZN(n713) );
  NOR2_X1 U643 ( .A1(n715), .A2(n713), .ZN(n536) );
  XNOR2_X1 U644 ( .A(n536), .B(KEYINPUT41), .ZN(n708) );
  INV_X1 U645 ( .A(n698), .ZN(n537) );
  NOR2_X1 U646 ( .A1(n568), .A2(n537), .ZN(n538) );
  INV_X1 U647 ( .A(n699), .ZN(n630) );
  NAND2_X1 U648 ( .A1(n538), .A2(n630), .ZN(n546) );
  NOR2_X1 U649 ( .A1(n539), .A2(n546), .ZN(n540) );
  XNOR2_X1 U650 ( .A(n540), .B(KEYINPUT28), .ZN(n558) );
  NAND2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n541) );
  NOR2_X1 U652 ( .A1(n708), .A2(n541), .ZN(n542) );
  XNOR2_X1 U653 ( .A(n542), .B(KEYINPUT42), .ZN(n779) );
  XNOR2_X1 U654 ( .A(n545), .B(KEYINPUT6), .ZN(n629) );
  INV_X1 U655 ( .A(n555), .ZN(n547) );
  INV_X1 U656 ( .A(n415), .ZN(n548) );
  OR2_X2 U657 ( .A1(n566), .A2(n551), .ZN(n674) );
  XNOR2_X2 U658 ( .A(n674), .B(n552), .ZN(n584) );
  NAND2_X1 U659 ( .A1(n553), .A2(n584), .ZN(n554) );
  XOR2_X1 U660 ( .A(KEYINPUT19), .B(KEYINPUT69), .Z(n556) );
  INV_X1 U661 ( .A(KEYINPUT83), .ZN(n560) );
  INV_X1 U662 ( .A(KEYINPUT47), .ZN(n562) );
  XNOR2_X1 U663 ( .A(n563), .B(n562), .ZN(n574) );
  NAND2_X1 U664 ( .A1(n628), .A2(n684), .ZN(n564) );
  NAND2_X1 U665 ( .A1(KEYINPUT83), .A2(n564), .ZN(n572) );
  NAND2_X1 U666 ( .A1(n566), .A2(n565), .ZN(n615) );
  NAND2_X1 U667 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U668 ( .A(n575), .B(KEYINPUT76), .ZN(n576) );
  NAND2_X1 U669 ( .A1(n577), .A2(n711), .ZN(n578) );
  XOR2_X1 U670 ( .A(n578), .B(KEYINPUT110), .Z(n579) );
  NAND2_X1 U671 ( .A1(n579), .A2(n415), .ZN(n580) );
  XNOR2_X1 U672 ( .A(n580), .B(KEYINPUT43), .ZN(n582) );
  NAND2_X1 U673 ( .A1(n582), .A2(n581), .ZN(n692) );
  OR2_X1 U674 ( .A1(n585), .A2(n584), .ZN(n691) );
  NOR2_X1 U675 ( .A1(G898), .A2(n586), .ZN(n587) );
  NOR2_X1 U676 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U677 ( .A1(n723), .A2(n589), .ZN(n590) );
  NAND2_X1 U678 ( .A1(n592), .A2(n698), .ZN(n593) );
  XOR2_X1 U679 ( .A(KEYINPUT101), .B(n593), .Z(n594) );
  XNOR2_X1 U680 ( .A(n633), .B(KEYINPUT104), .ZN(n598) );
  NOR2_X1 U681 ( .A1(n596), .A2(n699), .ZN(n597) );
  NOR2_X1 U682 ( .A1(n695), .A2(n699), .ZN(n599) );
  XNOR2_X1 U683 ( .A(KEYINPUT102), .B(n599), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n604) );
  INV_X1 U685 ( .A(KEYINPUT32), .ZN(n603) );
  XNOR2_X1 U686 ( .A(n604), .B(n603), .ZN(n777) );
  INV_X1 U687 ( .A(n777), .ZN(n605) );
  INV_X1 U688 ( .A(KEYINPUT67), .ZN(n607) );
  INV_X1 U689 ( .A(KEYINPUT105), .ZN(n609) );
  XNOR2_X1 U690 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n611), .B(KEYINPUT75), .ZN(n612) );
  XNOR2_X1 U692 ( .A(n614), .B(n613), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n616), .A2(n455), .ZN(n618) );
  XNOR2_X1 U694 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n617) );
  OR2_X1 U695 ( .A1(KEYINPUT67), .A2(KEYINPUT44), .ZN(n619) );
  INV_X1 U696 ( .A(n620), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n621), .A2(n545), .ZN(n704) );
  XNOR2_X1 U698 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n622) );
  INV_X1 U699 ( .A(n624), .ZN(n627) );
  OR2_X1 U700 ( .A1(n694), .A2(n545), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n675) );
  INV_X1 U702 ( .A(n628), .ZN(n714) );
  INV_X1 U703 ( .A(n629), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n671) );
  INV_X1 U706 ( .A(KEYINPUT2), .ZN(n731) );
  INV_X1 U707 ( .A(n637), .ZN(n638) );
  INV_X1 U708 ( .A(KEYINPUT66), .ZN(n639) );
  NAND2_X1 U709 ( .A1(KEYINPUT2), .A2(n691), .ZN(n640) );
  XOR2_X1 U710 ( .A(KEYINPUT82), .B(n640), .Z(n641) );
  XNOR2_X2 U711 ( .A(n643), .B(KEYINPUT65), .ZN(n663) );
  NAND2_X1 U712 ( .A1(n747), .A2(G478), .ZN(n645) );
  AND2_X1 U713 ( .A1(n724), .A2(G953), .ZN(n752) );
  NAND2_X1 U714 ( .A1(n663), .A2(G472), .ZN(n649) );
  XOR2_X1 U715 ( .A(KEYINPUT62), .B(n647), .Z(n648) );
  XNOR2_X1 U716 ( .A(n649), .B(n648), .ZN(n650) );
  INV_X1 U717 ( .A(n650), .ZN(n652) );
  NAND2_X1 U718 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U720 ( .A(n654), .B(G122), .Z(G24) );
  NAND2_X1 U721 ( .A1(n663), .A2(G475), .ZN(n659) );
  XOR2_X1 U722 ( .A(KEYINPUT68), .B(KEYINPUT88), .Z(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(KEYINPUT59), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n659), .B(n658), .ZN(n660) );
  NOR2_X2 U725 ( .A1(n660), .A2(n752), .ZN(n662) );
  XNOR2_X1 U726 ( .A(KEYINPUT70), .B(KEYINPUT60), .ZN(n661) );
  XNOR2_X1 U727 ( .A(n662), .B(n661), .ZN(G60) );
  NAND2_X1 U728 ( .A1(n663), .A2(G210), .ZN(n667) );
  XNOR2_X1 U729 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n667), .B(n666), .ZN(n668) );
  NOR2_X2 U732 ( .A1(n668), .A2(n752), .ZN(n670) );
  XNOR2_X1 U733 ( .A(KEYINPUT120), .B(KEYINPUT56), .ZN(n669) );
  XNOR2_X1 U734 ( .A(n670), .B(n669), .ZN(G51) );
  XNOR2_X1 U735 ( .A(G101), .B(n671), .ZN(G3) );
  NOR2_X1 U736 ( .A1(n675), .A2(n687), .ZN(n673) );
  XNOR2_X1 U737 ( .A(G104), .B(KEYINPUT113), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n673), .B(n672), .ZN(G6) );
  NOR2_X1 U739 ( .A1(n675), .A2(n674), .ZN(n680) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n677) );
  XNOR2_X1 U741 ( .A(G107), .B(KEYINPUT26), .ZN(n676) );
  XNOR2_X1 U742 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U743 ( .A(KEYINPUT114), .B(n678), .ZN(n679) );
  XNOR2_X1 U744 ( .A(n680), .B(n679), .ZN(G9) );
  NOR2_X1 U745 ( .A1(n684), .A2(n674), .ZN(n682) );
  XNOR2_X1 U746 ( .A(G128), .B(KEYINPUT29), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n682), .B(n681), .ZN(G30) );
  XOR2_X1 U748 ( .A(G143), .B(n683), .Z(G45) );
  NOR2_X1 U749 ( .A1(n687), .A2(n684), .ZN(n685) );
  XOR2_X1 U750 ( .A(KEYINPUT116), .B(n685), .Z(n686) );
  XNOR2_X1 U751 ( .A(G146), .B(n686), .ZN(G48) );
  NOR2_X1 U752 ( .A1(n689), .A2(n687), .ZN(n688) );
  XOR2_X1 U753 ( .A(G113), .B(n688), .Z(G15) );
  NOR2_X1 U754 ( .A1(n689), .A2(n674), .ZN(n690) );
  XOR2_X1 U755 ( .A(G116), .B(n690), .Z(G18) );
  XNOR2_X1 U756 ( .A(G134), .B(n691), .ZN(G36) );
  XNOR2_X1 U757 ( .A(G140), .B(n692), .ZN(G42) );
  NOR2_X1 U758 ( .A1(n708), .A2(n718), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n693), .A2(G953), .ZN(n728) );
  XNOR2_X1 U760 ( .A(KEYINPUT51), .B(KEYINPUT118), .ZN(n707) );
  NAND2_X1 U761 ( .A1(n415), .A2(n694), .ZN(n696) );
  XOR2_X1 U762 ( .A(KEYINPUT117), .B(n696), .Z(n697) );
  XNOR2_X1 U763 ( .A(n697), .B(KEYINPUT50), .ZN(n703) );
  NOR2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U765 ( .A(KEYINPUT49), .B(n700), .Z(n701) );
  NOR2_X1 U766 ( .A1(n545), .A2(n701), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n705) );
  NAND2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U769 ( .A(n707), .B(n706), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n720) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n719) );
  NOR2_X1 U775 ( .A1(n720), .A2(n370), .ZN(n721) );
  XNOR2_X1 U776 ( .A(n721), .B(KEYINPUT52), .ZN(n722) );
  XNOR2_X1 U777 ( .A(n722), .B(KEYINPUT119), .ZN(n726) );
  NOR2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U780 ( .A1(n728), .A2(n727), .ZN(n739) );
  NOR2_X1 U781 ( .A1(KEYINPUT2), .A2(n363), .ZN(n730) );
  XNOR2_X1 U782 ( .A(KEYINPUT85), .B(n730), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n734), .A2(n733), .ZN(n737) );
  INV_X1 U785 ( .A(n735), .ZN(n736) );
  NOR2_X1 U786 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U787 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U788 ( .A(n740), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U789 ( .A1(n747), .A2(G469), .ZN(n745) );
  XOR2_X1 U790 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n741) );
  XOR2_X1 U791 ( .A(n741), .B(KEYINPUT121), .Z(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(n744) );
  XNOR2_X1 U793 ( .A(n745), .B(n744), .ZN(n746) );
  NOR2_X1 U794 ( .A1(n752), .A2(n746), .ZN(G54) );
  NAND2_X1 U795 ( .A1(n747), .A2(G217), .ZN(n750) );
  XNOR2_X1 U796 ( .A(n748), .B(KEYINPUT122), .ZN(n749) );
  XNOR2_X1 U797 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U798 ( .A1(n752), .A2(n751), .ZN(G66) );
  XNOR2_X1 U799 ( .A(n753), .B(G110), .ZN(n755) );
  NOR2_X1 U800 ( .A1(n767), .A2(G898), .ZN(n754) );
  NOR2_X1 U801 ( .A1(n755), .A2(n754), .ZN(n763) );
  XNOR2_X1 U802 ( .A(n756), .B(KEYINPUT124), .ZN(n761) );
  XOR2_X1 U803 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n758) );
  NAND2_X1 U804 ( .A1(G224), .A2(G953), .ZN(n757) );
  XNOR2_X1 U805 ( .A(n758), .B(n757), .ZN(n759) );
  NAND2_X1 U806 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U808 ( .A(n763), .B(n762), .ZN(G69) );
  XNOR2_X1 U809 ( .A(n764), .B(KEYINPUT125), .ZN(n765) );
  XNOR2_X1 U810 ( .A(n766), .B(n765), .ZN(n770) );
  XOR2_X1 U811 ( .A(n770), .B(n363), .Z(n768) );
  NAND2_X1 U812 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U813 ( .A(n769), .B(KEYINPUT126), .ZN(n774) );
  XNOR2_X1 U814 ( .A(G227), .B(n770), .ZN(n771) );
  NAND2_X1 U815 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U816 ( .A1(G953), .A2(n772), .ZN(n773) );
  NAND2_X1 U817 ( .A1(n774), .A2(n773), .ZN(G72) );
  XOR2_X1 U818 ( .A(n775), .B(G125), .Z(n776) );
  XNOR2_X1 U819 ( .A(KEYINPUT37), .B(n776), .ZN(G27) );
  XOR2_X1 U820 ( .A(G119), .B(n777), .Z(G21) );
  XOR2_X1 U821 ( .A(n778), .B(G131), .Z(G33) );
  XOR2_X1 U822 ( .A(G137), .B(n779), .Z(G39) );
endmodule

