//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969;
  AND2_X1   g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n209), .B1(new_n215), .B2(KEYINPUT82), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT82), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(new_n212), .B2(new_n214), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n208), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n206), .A2(KEYINPUT15), .ZN(new_n220));
  INV_X1    g019(.A(new_n215), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n207), .A4(new_n209), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT17), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT96), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n226), .A2(G85gat), .A3(G92gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n226), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(G99gat), .B(G106gat), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G92gat), .ZN(new_n234));
  AND2_X1   g033(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT97), .A2(G85gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G99gat), .ZN(new_n238));
  INV_X1    g037(.A(G106gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT8), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n231), .A2(new_n233), .A3(new_n237), .A4(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n237), .A2(new_n229), .A3(new_n240), .A4(new_n230), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n232), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n219), .A2(new_n222), .A3(KEYINPUT17), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT98), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n202), .A2(KEYINPUT41), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n241), .A2(new_n243), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n223), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n246), .A2(KEYINPUT98), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(G134gat), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n249), .A2(new_n255), .A3(new_n251), .A4(new_n252), .ZN(new_n256));
  XNOR2_X1  g055(.A(G190gat), .B(G218gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n254), .B2(new_n256), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n205), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n204), .A3(new_n259), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT92), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT91), .ZN(new_n268));
  INV_X1    g067(.A(G64gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G57gat), .ZN(new_n270));
  INV_X1    g069(.A(G57gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G64gat), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n270), .A2(new_n272), .A3(new_n268), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n267), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(G71gat), .A2(G78gat), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT90), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(KEYINPUT90), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n277), .A2(new_n278), .B1(G71gat), .B2(G78gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(G71gat), .A2(G78gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n270), .A2(new_n272), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n275), .A2(new_n279), .B1(new_n267), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n283), .A2(KEYINPUT21), .ZN(new_n284));
  INV_X1    g083(.A(G15gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G22gat), .ZN(new_n286));
  INV_X1    g085(.A(G22gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G15gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT16), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(G1gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n290), .B(KEYINPUT84), .C1(G1gat), .C2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G8gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n290), .B(KEYINPUT83), .C1(G1gat), .C2(new_n291), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n292), .A2(new_n293), .A3(G8gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OR3_X1    g098(.A1(new_n284), .A2(new_n299), .A3(KEYINPUT95), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT95), .B1(new_n284), .B2(new_n299), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n300), .A2(KEYINPUT20), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT20), .B1(new_n300), .B2(new_n301), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n274), .A2(new_n273), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT92), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n266), .B(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n279), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n267), .A2(new_n282), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G231gat), .A2(G233gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  OR3_X1    g112(.A1(new_n302), .A2(new_n303), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n313), .B1(new_n302), .B2(new_n303), .ZN(new_n315));
  XOR2_X1   g114(.A(G183gat), .B(G211gat), .Z(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G127gat), .B(G155gat), .Z(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  AND3_X1   g119(.A1(new_n314), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n314), .B2(new_n315), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT100), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n241), .A4(new_n243), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n250), .A2(new_n283), .A3(KEYINPUT100), .A4(KEYINPUT10), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n244), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n329), .A2(new_n332), .B1(G230gat), .B2(G233gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(G230gat), .A2(G233gat), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n330), .B2(new_n325), .ZN(new_n335));
  XNOR2_X1  g134(.A(G120gat), .B(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(G176gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G204gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n333), .A2(new_n335), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n334), .B(KEYINPUT101), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n344), .B1(new_n329), .B2(new_n332), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n340), .B1(new_n345), .B2(new_n335), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n265), .A2(new_n323), .A3(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n292), .A2(new_n293), .A3(G8gat), .ZN(new_n350));
  AOI21_X1  g149(.A(G8gat), .B1(new_n292), .B2(new_n293), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n225), .A2(new_n352), .A3(new_n297), .A4(new_n245), .ZN(new_n353));
  NAND2_X1  g152(.A1(G229gat), .A2(G233gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT85), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n299), .A2(new_n223), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT88), .B1(new_n299), .B2(new_n223), .ZN(new_n358));
  INV_X1    g157(.A(new_n223), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n352), .A2(new_n359), .A3(new_n360), .A4(new_n297), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n355), .B(KEYINPUT13), .Z(new_n363));
  AOI22_X1  g162(.A1(new_n357), .A2(KEYINPUT18), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT18), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n366), .A2(KEYINPUT86), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(KEYINPUT86), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n365), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT87), .ZN(new_n370));
  XNOR2_X1  g169(.A(G113gat), .B(G141gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n371), .B(G197gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT11), .ZN(new_n373));
  INV_X1    g172(.A(G169gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT12), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n373), .B(G169gat), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT12), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n364), .B(new_n369), .C1(new_n370), .C2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n362), .A2(new_n363), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n353), .A2(KEYINPUT18), .A3(new_n355), .A4(new_n356), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n369), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n380), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n370), .A3(new_n383), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT89), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n381), .A2(new_n387), .A3(KEYINPUT89), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(KEYINPUT74), .B(G197gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(new_n339), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT22), .ZN(new_n396));
  INV_X1    g195(.A(G211gat), .ZN(new_n397));
  INV_X1    g196(.A(G218gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(G211gat), .B(G218gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n401), .A3(new_n399), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G141gat), .B(G148gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT2), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT76), .B(G162gat), .ZN(new_n415));
  INV_X1    g214(.A(G155gat), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT2), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n407), .A2(new_n418), .A3(new_n408), .ZN(new_n419));
  AND2_X1   g218(.A1(G155gat), .A2(G162gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(G155gat), .A2(G162gat), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT75), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n423), .A3(new_n411), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n414), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n406), .B1(KEYINPUT29), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n414), .A2(new_n424), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT29), .B1(new_n403), .B2(new_n404), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(KEYINPUT3), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n430), .A3(new_n287), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n287), .B1(new_n427), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT31), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n433), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT31), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n431), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n430), .A2(KEYINPUT81), .ZN(new_n438));
  XOR2_X1   g237(.A(G78gat), .B(G106gat), .Z(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(G50gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT80), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n438), .A2(G228gat), .A3(G233gat), .A4(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n438), .A2(G228gat), .A3(G233gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n441), .ZN(new_n445));
  AND4_X1   g244(.A1(new_n434), .A2(new_n437), .A3(new_n443), .A4(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n437), .A2(new_n434), .B1(new_n445), .B2(new_n443), .ZN(new_n447));
  OR2_X1    g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449));
  XNOR2_X1  g248(.A(G15gat), .B(G43gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(G71gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G99gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT72), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n453), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT26), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n374), .A3(new_n337), .ZN(new_n461));
  OAI211_X1 g260(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G183gat), .A2(G190gat), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(G183gat), .ZN(new_n468));
  INV_X1    g267(.A(G183gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT27), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT28), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(G190gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n466), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n473), .A2(new_n468), .A3(new_n470), .A4(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(KEYINPUT66), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479));
  AOI21_X1  g278(.A(G190gat), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT28), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n465), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G113gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(G120gat), .ZN(new_n484));
  INV_X1    g283(.A(G120gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(G113gat), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT1), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(G127gat), .B(G134gat), .Z(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(G127gat), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n490), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(G127gat), .B(G134gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(KEYINPUT69), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n493), .B2(new_n487), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT25), .ZN(new_n495));
  NOR2_X1   g294(.A1(G183gat), .A2(G190gat), .ZN(new_n496));
  AND2_X1   g295(.A1(G183gat), .A2(G190gat), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(KEYINPUT24), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n464), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n464), .A2(KEYINPUT65), .A3(new_n499), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OR3_X1    g303(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n505), .A2(new_n506), .B1(G169gat), .B2(G176gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n495), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n498), .A2(new_n500), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n498), .A2(KEYINPUT64), .A3(new_n500), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(new_n495), .A3(new_n507), .A4(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n482), .A2(new_n494), .A3(new_n509), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT70), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n482), .A2(new_n509), .A3(new_n514), .ZN(new_n517));
  INV_X1    g316(.A(new_n494), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G190gat), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n469), .A2(KEYINPUT27), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(KEYINPUT66), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n479), .B1(new_n468), .B2(new_n470), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n472), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n475), .A3(new_n476), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n508), .B1(new_n525), .B2(new_n465), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(new_n527), .A3(new_n494), .A4(new_n514), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n516), .A2(new_n519), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G227gat), .A2(G233gat), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n529), .A2(KEYINPUT71), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT71), .B1(new_n529), .B2(new_n531), .ZN(new_n533));
  OAI211_X1 g332(.A(KEYINPUT32), .B(new_n455), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n449), .A2(KEYINPUT32), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n531), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n529), .A2(KEYINPUT71), .A3(new_n531), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n534), .B1(new_n540), .B2(new_n452), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n516), .A2(new_n519), .A3(new_n528), .A4(new_n530), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT34), .Z(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n534), .B(new_n543), .C1(new_n540), .C2(new_n452), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(KEYINPUT73), .A3(new_n544), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n448), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n414), .A2(new_n494), .A3(new_n424), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT78), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n410), .B1(new_n419), .B2(new_n422), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n413), .B1(new_n417), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n556), .A2(KEYINPUT78), .A3(new_n551), .A4(new_n494), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n414), .A2(new_n494), .A3(new_n424), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT4), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n554), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G225gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT77), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n425), .B1(new_n414), .B2(new_n424), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n425), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n518), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT5), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n428), .A2(new_n518), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n558), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n569), .B1(new_n571), .B2(new_n562), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n426), .A2(new_n564), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n573), .A2(new_n518), .B1(new_n559), .B2(new_n552), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n562), .A2(KEYINPUT5), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n568), .A2(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT79), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n578));
  XNOR2_X1  g377(.A(G1gat), .B(G29gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT0), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G57gat), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(G85gat), .Z(new_n582));
  NOR4_X1   g381(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n572), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n574), .A2(new_n575), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n577), .B1(new_n589), .B2(new_n578), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT6), .B1(new_n576), .B2(new_n582), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n589), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G8gat), .B(G36gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(new_n269), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(new_n234), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT29), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n517), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G226gat), .ZN(new_n599));
  INV_X1    g398(.A(G233gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n526), .B2(new_n514), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n405), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n601), .B1(new_n517), .B2(new_n597), .ZN(new_n607));
  NOR3_X1   g406(.A1(new_n607), .A2(new_n604), .A3(new_n406), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n596), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n603), .A2(new_n405), .A3(new_n605), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n406), .B1(new_n607), .B2(new_n604), .ZN(new_n611));
  INV_X1    g410(.A(new_n596), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n609), .A2(KEYINPUT30), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT30), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n610), .A2(new_n611), .A3(new_n615), .A4(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n593), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT35), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n614), .A2(new_n616), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT79), .B1(new_n622), .B2(KEYINPUT6), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n623), .A2(new_n583), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n624), .B2(new_n592), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n446), .A2(new_n447), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n625), .A2(new_n545), .A3(new_n547), .A4(new_n626), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n550), .A2(new_n620), .B1(new_n627), .B2(new_n619), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n548), .A2(KEYINPUT36), .A3(new_n549), .ZN(new_n629));
  INV_X1    g428(.A(new_n613), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT37), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n606), .B2(new_n608), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n610), .A2(KEYINPUT37), .A3(new_n611), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n612), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n630), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n606), .A2(new_n608), .A3(new_n631), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT37), .B1(new_n610), .B2(new_n611), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n596), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT38), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n636), .A2(new_n624), .A3(new_n640), .A4(new_n592), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n559), .A2(new_n552), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n567), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n562), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT39), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n588), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n644), .B(KEYINPUT39), .C1(new_n562), .C2(new_n571), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n646), .A2(KEYINPUT40), .A3(new_n647), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n621), .A2(new_n589), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n641), .A2(new_n652), .A3(new_n626), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n448), .A2(new_n618), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT36), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n545), .A2(new_n655), .A3(new_n547), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n629), .A2(new_n653), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  AOI211_X1 g456(.A(new_n349), .B(new_n393), .C1(new_n628), .C2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n593), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g460(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n621), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n663), .B1(new_n289), .B2(new_n295), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n295), .B1(new_n658), .B2(new_n621), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT42), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(KEYINPUT42), .B2(new_n664), .ZN(G1325gat));
  AND2_X1   g466(.A1(new_n545), .A2(new_n547), .ZN(new_n668));
  AOI21_X1  g467(.A(G15gat), .B1(new_n658), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n629), .A2(new_n656), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n670), .A2(new_n285), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n658), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n658), .A2(new_n448), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND2_X1  g474(.A1(new_n262), .A2(new_n264), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n550), .A2(new_n620), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n627), .A2(new_n619), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n657), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n323), .A2(new_n347), .ZN(new_n680));
  AND4_X1   g479(.A1(new_n676), .A2(new_n679), .A3(new_n392), .A4(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n210), .A3(new_n659), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT45), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n676), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n265), .B1(new_n628), .B2(new_n657), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n388), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n323), .A2(new_n347), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n659), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n683), .B1(new_n210), .B2(new_n693), .ZN(G1328gat));
  NAND3_X1  g493(.A1(new_n681), .A2(new_n211), .A3(new_n621), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n681), .A2(KEYINPUT102), .A3(new_n211), .A4(new_n621), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n689), .A2(new_n621), .A3(new_n691), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G36gat), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n697), .A2(new_n699), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n702), .B(new_n704), .C1(new_n698), .C2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(new_n670), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT44), .B(new_n265), .C1(new_n628), .C2(new_n657), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n687), .B1(new_n679), .B2(new_n676), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n707), .B(new_n691), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT106), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n689), .A2(new_n712), .A3(new_n707), .A4(new_n691), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n713), .A3(G43gat), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n686), .A2(new_n668), .A3(new_n392), .A4(new_n680), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT105), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n681), .A2(new_n718), .A3(new_n719), .A4(new_n668), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n715), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n714), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n717), .A2(new_n720), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n710), .A2(G43gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT107), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n722), .A2(new_n726), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1330gat));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n689), .A2(new_n448), .A3(new_n691), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G50gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n734), .B2(KEYINPUT109), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n626), .A2(G50gat), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT108), .Z(new_n737));
  AOI22_X1  g536(.A1(new_n733), .A2(G50gat), .B1(new_n681), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n735), .B(new_n738), .ZN(G1331gat));
  INV_X1    g538(.A(new_n323), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n676), .A2(new_n740), .A3(new_n348), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n679), .A2(new_n690), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n593), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(new_n271), .ZN(G1332gat));
  NAND2_X1  g543(.A1(new_n742), .A2(KEYINPUT110), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT110), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n679), .A2(new_n746), .A3(new_n690), .A4(new_n741), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n617), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  INV_X1    g553(.A(G71gat), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n748), .B2(new_n707), .ZN(new_n756));
  INV_X1    g555(.A(new_n742), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n668), .A2(new_n755), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(KEYINPUT50), .ZN(G1334gat));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n748), .B2(new_n448), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g562(.A(KEYINPUT112), .B(new_n626), .C1(new_n745), .C2(new_n747), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT111), .B1(new_n762), .B2(new_n764), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n767), .A2(G78gat), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(G78gat), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(G1335gat));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n740), .A2(new_n690), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n684), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n773), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT51), .B1(new_n686), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  MUX2_X1   g576(.A(new_n774), .B(new_n777), .S(KEYINPUT113), .Z(new_n778));
  OR2_X1    g577(.A1(new_n235), .A2(new_n236), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n659), .A2(new_n779), .A3(new_n347), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n689), .A2(new_n347), .A3(new_n775), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n593), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n778), .A2(new_n780), .B1(new_n779), .B2(new_n782), .ZN(G1336gat));
  NOR3_X1   g582(.A1(new_n348), .A2(new_n617), .A3(G92gat), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n777), .A2(KEYINPUT114), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(G92gat), .B1(new_n781), .B2(new_n617), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT114), .B1(new_n777), .B2(new_n785), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT52), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n778), .B2(new_n785), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(G1337gat));
  OAI21_X1  g592(.A(G99gat), .B1(new_n781), .B2(new_n670), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n668), .A2(new_n238), .A3(new_n347), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n778), .B2(new_n795), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n448), .A2(new_n239), .A3(new_n347), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n778), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G106gat), .B1(new_n781), .B2(new_n626), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n797), .B(KEYINPUT116), .Z(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n774), .B2(new_n776), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n798), .A2(new_n801), .B1(new_n804), .B2(new_n800), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n329), .A2(new_n332), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n334), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n329), .A2(new_n344), .A3(new_n332), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n808), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT54), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n807), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n329), .A2(new_n344), .A3(new_n332), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT117), .B1(new_n816), .B2(new_n333), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n818), .B1(new_n811), .B2(new_n808), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(KEYINPUT118), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n345), .A2(new_n818), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n340), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n806), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT55), .B(new_n823), .C1(new_n815), .C2(new_n820), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n342), .B(new_n388), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n384), .A2(new_n385), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n353), .A2(new_n356), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n829), .A2(new_n355), .B1(new_n362), .B2(new_n363), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n375), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n347), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n676), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n342), .B(new_n831), .C1(new_n825), .C2(new_n826), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n265), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n740), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n349), .A2(new_n388), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n593), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n668), .A2(new_n626), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n617), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n393), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n837), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n659), .A3(new_n550), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT120), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n838), .A2(new_n847), .A3(new_n550), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n621), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n483), .A3(new_n388), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n843), .A2(new_n850), .ZN(G1340gat));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n485), .A3(new_n347), .ZN(new_n852));
  OAI21_X1  g651(.A(G120gat), .B1(new_n841), .B2(new_n348), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1341gat));
  NAND2_X1  g653(.A1(new_n846), .A2(new_n848), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n323), .A3(new_n617), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT121), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n849), .A2(new_n858), .A3(new_n323), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n490), .A3(new_n859), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n841), .A2(new_n490), .A3(new_n740), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(G1342gat));
  NOR2_X1   g661(.A1(new_n265), .A2(G134gat), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n838), .A2(new_n847), .A3(new_n550), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n847), .B1(new_n838), .B2(new_n550), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n617), .B(new_n863), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n841), .B2(new_n265), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n855), .A2(new_n869), .A3(new_n617), .A4(new_n863), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT122), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n867), .A2(new_n870), .A3(new_n873), .A4(new_n868), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(new_n837), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n342), .B(new_n392), .C1(new_n825), .C2(new_n826), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n832), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n265), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT123), .ZN(new_n880));
  INV_X1    g679(.A(new_n835), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n676), .B1(new_n877), .B2(new_n832), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n876), .B1(new_n885), .B2(new_n740), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT57), .B1(new_n886), .B2(new_n626), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n626), .B1(new_n836), .B2(new_n837), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n670), .A2(new_n659), .A3(new_n617), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(G141gat), .B1(new_n893), .B2(new_n393), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n888), .A2(new_n892), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(G141gat), .A3(new_n393), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(KEYINPUT58), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n887), .A2(new_n388), .A3(new_n890), .A4(new_n892), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n896), .B1(new_n900), .B2(G141gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(G1344gat));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n903), .B(G148gat), .C1(new_n893), .C2(new_n348), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n626), .A2(KEYINPUT57), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n740), .B1(new_n882), .B2(new_n835), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n349), .A2(new_n392), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n844), .A2(new_n448), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n347), .ZN(new_n912));
  OAI21_X1  g711(.A(G148gat), .B1(new_n912), .B2(new_n891), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT59), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n904), .A2(new_n914), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n895), .A2(G148gat), .A3(new_n348), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1345gat));
  OAI21_X1  g716(.A(G155gat), .B1(new_n893), .B2(new_n740), .ZN(new_n918));
  INV_X1    g717(.A(new_n895), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n416), .A3(new_n323), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n918), .A2(new_n920), .ZN(G1346gat));
  NAND3_X1  g720(.A1(new_n919), .A2(new_n415), .A3(new_n676), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n893), .A2(new_n265), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n415), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n659), .A2(new_n617), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n844), .A2(new_n550), .A3(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n374), .A3(new_n388), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n925), .B(KEYINPUT124), .Z(new_n929));
  AND3_X1   g728(.A1(new_n844), .A2(new_n840), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(new_n392), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n374), .ZN(G1348gat));
  AOI21_X1  g731(.A(G176gat), .B1(new_n927), .B2(new_n347), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n348), .A2(new_n337), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n930), .B2(new_n934), .ZN(G1349gat));
  AOI21_X1  g734(.A(new_n469), .B1(new_n930), .B2(new_n323), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n926), .A2(new_n740), .A3(new_n471), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g738(.A(new_n520), .B1(new_n930), .B2(new_n676), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT61), .Z(new_n941));
  NAND3_X1  g740(.A1(new_n927), .A2(new_n520), .A3(new_n676), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1351gat));
  AND3_X1   g742(.A1(new_n888), .A2(new_n670), .A3(new_n925), .ZN(new_n944));
  XNOR2_X1  g743(.A(KEYINPUT125), .B(G197gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n944), .A2(new_n388), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n907), .A2(new_n908), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n905), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n929), .A2(new_n670), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n949), .B(new_n950), .C1(new_n889), .C2(new_n888), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n393), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n947), .B1(new_n952), .B2(new_n945), .ZN(G1352gat));
  NAND3_X1  g752(.A1(new_n944), .A2(new_n339), .A3(new_n347), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  AND3_X1   g754(.A1(new_n911), .A2(new_n347), .A3(new_n950), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n955), .B1(new_n339), .B2(new_n956), .ZN(G1353gat));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n951), .B2(new_n740), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n911), .A2(KEYINPUT127), .A3(new_n323), .A4(new_n950), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(G211gat), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n944), .A2(new_n397), .A3(new_n323), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1354gat));
  NOR3_X1   g766(.A1(new_n951), .A2(new_n398), .A3(new_n265), .ZN(new_n968));
  AOI21_X1  g767(.A(G218gat), .B1(new_n944), .B2(new_n676), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(new_n969), .ZN(G1355gat));
endmodule


