

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U552 ( .A(KEYINPUT92), .B(n659), .Z(n714) );
  NOR2_X1 U553 ( .A1(G2104), .A2(n536), .ZN(n882) );
  INV_X1 U554 ( .A(G2105), .ZN(n536) );
  NOR2_X1 U555 ( .A1(n696), .A2(n695), .ZN(n698) );
  NOR2_X2 U556 ( .A1(n574), .A2(n521), .ZN(n604) );
  XNOR2_X2 U557 ( .A(n533), .B(n532), .ZN(n722) );
  NOR2_X1 U558 ( .A1(n658), .A2(n959), .ZN(n625) );
  XNOR2_X1 U559 ( .A(n625), .B(KEYINPUT26), .ZN(n626) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n666) );
  BUF_X1 U561 ( .A(n658), .Z(n671) );
  AND2_X1 U562 ( .A1(n710), .A2(n690), .ZN(n696) );
  NOR2_X1 U563 ( .A1(G164), .A2(n622), .ZN(n624) );
  INV_X1 U564 ( .A(KEYINPUT101), .ZN(n697) );
  NAND2_X1 U565 ( .A1(n624), .A2(n623), .ZN(n658) );
  INV_X1 U566 ( .A(KEYINPUT103), .ZN(n718) );
  INV_X1 U567 ( .A(KEYINPUT73), .ZN(n610) );
  XNOR2_X1 U568 ( .A(n610), .B(KEYINPUT13), .ZN(n611) );
  NOR2_X1 U569 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U570 ( .A1(G651), .A2(G543), .ZN(n814) );
  XNOR2_X1 U571 ( .A(n612), .B(n611), .ZN(n616) );
  AND2_X1 U572 ( .A1(n536), .A2(G2104), .ZN(n879) );
  NAND2_X1 U573 ( .A1(n618), .A2(n617), .ZN(n983) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n574) );
  INV_X1 U575 ( .A(G651), .ZN(n521) );
  NAND2_X1 U576 ( .A1(G73), .A2(n604), .ZN(n519) );
  XOR2_X1 U577 ( .A(KEYINPUT2), .B(n519), .Z(n528) );
  NAND2_X1 U578 ( .A1(n814), .A2(G86), .ZN(n520) );
  XNOR2_X1 U579 ( .A(n520), .B(KEYINPUT84), .ZN(n525) );
  NOR2_X1 U580 ( .A1(G543), .A2(n521), .ZN(n523) );
  XNOR2_X1 U581 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n522) );
  XNOR2_X2 U582 ( .A(n523), .B(n522), .ZN(n817) );
  NAND2_X1 U583 ( .A1(G61), .A2(n817), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U585 ( .A(KEYINPUT85), .B(n526), .Z(n527) );
  NOR2_X1 U586 ( .A1(n528), .A2(n527), .ZN(n531) );
  NOR2_X1 U587 ( .A1(G651), .A2(n574), .ZN(n529) );
  XNOR2_X2 U588 ( .A(KEYINPUT64), .B(n529), .ZN(n812) );
  NAND2_X1 U589 ( .A1(G48), .A2(n812), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n531), .A2(n530), .ZN(G305) );
  XNOR2_X1 U591 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n533) );
  NOR2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  NAND2_X1 U593 ( .A1(G138), .A2(n722), .ZN(n535) );
  NAND2_X1 U594 ( .A1(G102), .A2(n879), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G126), .A2(n882), .ZN(n538) );
  AND2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U598 ( .A1(G114), .A2(n883), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U600 ( .A1(n540), .A2(n539), .ZN(G164) );
  NAND2_X1 U601 ( .A1(G91), .A2(n814), .ZN(n542) );
  NAND2_X1 U602 ( .A1(G65), .A2(n817), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n604), .A2(G78), .ZN(n543) );
  XOR2_X1 U605 ( .A(KEYINPUT68), .B(n543), .Z(n544) );
  NOR2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U607 ( .A1(G53), .A2(n812), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(G299) );
  NAND2_X1 U609 ( .A1(G64), .A2(n817), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G52), .A2(n812), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G77), .A2(n604), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G90), .A2(n814), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  NOR2_X1 U616 ( .A1(n554), .A2(n553), .ZN(G171) );
  NAND2_X1 U617 ( .A1(G89), .A2(n814), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT75), .B(n555), .Z(n556) );
  XNOR2_X1 U619 ( .A(n556), .B(KEYINPUT4), .ZN(n558) );
  NAND2_X1 U620 ( .A1(G76), .A2(n604), .ZN(n557) );
  NAND2_X1 U621 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U623 ( .A1(n817), .A2(G63), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n560), .B(KEYINPUT76), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G51), .A2(n812), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U629 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G88), .A2(n814), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G62), .A2(n817), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n604), .A2(G75), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT86), .B(n569), .Z(n570) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U637 ( .A1(G50), .A2(n812), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(G303) );
  INV_X1 U639 ( .A(G303), .ZN(G166) );
  NAND2_X1 U640 ( .A1(G87), .A2(n574), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n817), .A2(n577), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n812), .A2(G49), .ZN(n578) );
  XOR2_X1 U645 ( .A(KEYINPUT83), .B(n578), .Z(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(G288) );
  INV_X1 U647 ( .A(KEYINPUT66), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G137), .A2(n722), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G113), .A2(n883), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U651 ( .A1(n583), .A2(n584), .ZN(n586) );
  OR2_X1 U652 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n882), .A2(G125), .ZN(n587) );
  AND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n623) );
  NAND2_X1 U656 ( .A1(G101), .A2(n879), .ZN(n589) );
  XOR2_X1 U657 ( .A(n589), .B(KEYINPUT23), .Z(n619) );
  AND2_X1 U658 ( .A1(n623), .A2(n619), .ZN(G160) );
  NAND2_X1 U659 ( .A1(G72), .A2(n604), .ZN(n591) );
  NAND2_X1 U660 ( .A1(G85), .A2(n814), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G60), .A2(n817), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G47), .A2(n812), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n594) );
  OR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(G290) );
  XNOR2_X1 U666 ( .A(G1981), .B(G305), .ZN(n980) );
  NAND2_X1 U667 ( .A1(G92), .A2(n814), .ZN(n597) );
  NAND2_X1 U668 ( .A1(G66), .A2(n817), .ZN(n596) );
  NAND2_X1 U669 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U670 ( .A(KEYINPUT74), .B(n598), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G79), .A2(n604), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G54), .A2(n812), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U674 ( .A(KEYINPUT15), .B(n603), .Z(n903) );
  NAND2_X1 U675 ( .A1(n604), .A2(G68), .ZN(n606) );
  INV_X1 U676 ( .A(KEYINPUT72), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n606), .B(n605), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n814), .A2(G81), .ZN(n607) );
  XOR2_X1 U679 ( .A(KEYINPUT12), .B(n607), .Z(n608) );
  NOR2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U681 ( .A1(G56), .A2(n817), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n613), .B(KEYINPUT14), .ZN(n614) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n614), .ZN(n615) );
  NOR2_X1 U684 ( .A1(n616), .A2(n615), .ZN(n618) );
  NAND2_X1 U685 ( .A1(G43), .A2(n812), .ZN(n617) );
  INV_X1 U686 ( .A(G1384), .ZN(n621) );
  AND2_X1 U687 ( .A1(n619), .A2(G40), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n622) );
  INV_X1 U689 ( .A(G1996), .ZN(n959) );
  INV_X1 U690 ( .A(n626), .ZN(n628) );
  NAND2_X1 U691 ( .A1(n671), .A2(G1341), .ZN(n627) );
  NAND2_X1 U692 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U693 ( .A1(n983), .A2(n629), .ZN(n630) );
  OR2_X1 U694 ( .A1(n903), .A2(n630), .ZN(n637) );
  NAND2_X1 U695 ( .A1(n903), .A2(n630), .ZN(n635) );
  INV_X1 U696 ( .A(n658), .ZN(n652) );
  AND2_X1 U697 ( .A1(n652), .A2(G2067), .ZN(n631) );
  XNOR2_X1 U698 ( .A(n631), .B(KEYINPUT95), .ZN(n633) );
  NAND2_X1 U699 ( .A1(n671), .A2(G1348), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U702 ( .A1(n637), .A2(n636), .ZN(n639) );
  INV_X1 U703 ( .A(KEYINPUT96), .ZN(n638) );
  XNOR2_X1 U704 ( .A(n639), .B(n638), .ZN(n645) );
  NAND2_X1 U705 ( .A1(n652), .A2(G2072), .ZN(n640) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(n640), .Z(n642) );
  NAND2_X1 U707 ( .A1(G1956), .A2(n671), .ZN(n641) );
  NAND2_X1 U708 ( .A1(n642), .A2(n641), .ZN(n646) );
  NOR2_X1 U709 ( .A1(G299), .A2(n646), .ZN(n643) );
  XOR2_X1 U710 ( .A(KEYINPUT97), .B(n643), .Z(n644) );
  NOR2_X1 U711 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U712 ( .A1(G299), .A2(n646), .ZN(n647) );
  XOR2_X1 U713 ( .A(KEYINPUT28), .B(n647), .Z(n648) );
  NOR2_X1 U714 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U715 ( .A(n650), .B(KEYINPUT29), .ZN(n657) );
  NOR2_X1 U716 ( .A1(n652), .A2(G1961), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(KEYINPUT93), .ZN(n654) );
  XNOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .ZN(n961) );
  NAND2_X1 U719 ( .A1(n652), .A2(n961), .ZN(n653) );
  NAND2_X1 U720 ( .A1(n654), .A2(n653), .ZN(n663) );
  AND2_X1 U721 ( .A1(n663), .A2(G171), .ZN(n655) );
  XOR2_X1 U722 ( .A(KEYINPUT94), .B(n655), .Z(n656) );
  NAND2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n669) );
  NAND2_X1 U724 ( .A1(n658), .A2(G8), .ZN(n659) );
  INV_X1 U725 ( .A(n714), .ZN(n688) );
  NOR2_X1 U726 ( .A1(n688), .A2(G1966), .ZN(n684) );
  NOR2_X1 U727 ( .A1(G2084), .A2(n671), .ZN(n681) );
  NOR2_X1 U728 ( .A1(n684), .A2(n681), .ZN(n660) );
  NAND2_X1 U729 ( .A1(G8), .A2(n660), .ZN(n661) );
  XNOR2_X1 U730 ( .A(KEYINPUT30), .B(n661), .ZN(n662) );
  NOR2_X1 U731 ( .A1(G168), .A2(n662), .ZN(n665) );
  NOR2_X1 U732 ( .A1(G171), .A2(n663), .ZN(n664) );
  NOR2_X1 U733 ( .A1(n665), .A2(n664), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n682) );
  NAND2_X1 U736 ( .A1(n682), .A2(G286), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(KEYINPUT98), .ZN(n678) );
  NOR2_X1 U738 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U739 ( .A(KEYINPUT99), .B(n672), .ZN(n675) );
  NOR2_X1 U740 ( .A1(n688), .A2(G1971), .ZN(n673) );
  NOR2_X1 U741 ( .A1(G166), .A2(n673), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(KEYINPUT100), .B(n676), .ZN(n677) );
  NAND2_X1 U744 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U745 ( .A1(n679), .A2(G8), .ZN(n680) );
  XNOR2_X1 U746 ( .A(n680), .B(KEYINPUT32), .ZN(n710) );
  NAND2_X1 U747 ( .A1(G8), .A2(n681), .ZN(n686) );
  INV_X1 U748 ( .A(n682), .ZN(n683) );
  NOR2_X1 U749 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n686), .A2(n685), .ZN(n709) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n986) );
  INV_X1 U752 ( .A(n986), .ZN(n687) );
  OR2_X1 U753 ( .A1(n688), .A2(n687), .ZN(n692) );
  INV_X1 U754 ( .A(n692), .ZN(n689) );
  AND2_X1 U755 ( .A1(n709), .A2(n689), .ZN(n690) );
  NOR2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n700) );
  NOR2_X1 U757 ( .A1(G1971), .A2(G303), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n700), .A2(n691), .ZN(n993) );
  OR2_X1 U759 ( .A1(n692), .A2(n993), .ZN(n694) );
  INV_X1 U760 ( .A(KEYINPUT33), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U762 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X1 U763 ( .A1(n980), .A2(n699), .ZN(n704) );
  NAND2_X1 U764 ( .A1(n700), .A2(KEYINPUT33), .ZN(n701) );
  XOR2_X1 U765 ( .A(KEYINPUT102), .B(n701), .Z(n702) );
  NAND2_X1 U766 ( .A1(n702), .A2(n714), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n708) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n705), .B(KEYINPUT24), .ZN(n706) );
  NAND2_X1 U770 ( .A1(n706), .A2(n714), .ZN(n707) );
  NAND2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n717) );
  AND2_X1 U772 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U773 ( .A1(G166), .A2(G8), .ZN(n711) );
  NOR2_X1 U774 ( .A1(G2090), .A2(n711), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U777 ( .A1(n717), .A2(n716), .ZN(n719) );
  XNOR2_X1 U778 ( .A(n719), .B(n718), .ZN(n754) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n721) );
  NAND2_X1 U780 ( .A1(G160), .A2(G40), .ZN(n720) );
  NOR2_X1 U781 ( .A1(n721), .A2(n720), .ZN(n770) );
  XNOR2_X1 U782 ( .A(KEYINPUT37), .B(G2067), .ZN(n767) );
  NAND2_X1 U783 ( .A1(G140), .A2(n722), .ZN(n724) );
  NAND2_X1 U784 ( .A1(G104), .A2(n879), .ZN(n723) );
  NAND2_X1 U785 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U786 ( .A(KEYINPUT34), .B(n725), .ZN(n731) );
  NAND2_X1 U787 ( .A1(n883), .A2(G116), .ZN(n726) );
  XNOR2_X1 U788 ( .A(n726), .B(KEYINPUT88), .ZN(n728) );
  NAND2_X1 U789 ( .A1(G128), .A2(n882), .ZN(n727) );
  NAND2_X1 U790 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U791 ( .A(n729), .B(KEYINPUT35), .Z(n730) );
  NOR2_X1 U792 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U793 ( .A(KEYINPUT36), .B(n732), .Z(n733) );
  XNOR2_X1 U794 ( .A(KEYINPUT89), .B(n733), .ZN(n896) );
  NOR2_X1 U795 ( .A1(n767), .A2(n896), .ZN(n949) );
  NAND2_X1 U796 ( .A1(n770), .A2(n949), .ZN(n765) );
  NAND2_X1 U797 ( .A1(G119), .A2(n882), .ZN(n735) );
  NAND2_X1 U798 ( .A1(G107), .A2(n883), .ZN(n734) );
  NAND2_X1 U799 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U800 ( .A(KEYINPUT90), .B(n736), .ZN(n739) );
  NAND2_X1 U801 ( .A1(G95), .A2(n879), .ZN(n737) );
  XNOR2_X1 U802 ( .A(KEYINPUT91), .B(n737), .ZN(n738) );
  NOR2_X1 U803 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U804 ( .A1(n722), .A2(G131), .ZN(n740) );
  NAND2_X1 U805 ( .A1(n741), .A2(n740), .ZN(n891) );
  AND2_X1 U806 ( .A1(n891), .A2(G1991), .ZN(n750) );
  NAND2_X1 U807 ( .A1(G141), .A2(n722), .ZN(n743) );
  NAND2_X1 U808 ( .A1(G129), .A2(n882), .ZN(n742) );
  NAND2_X1 U809 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U810 ( .A1(n879), .A2(G105), .ZN(n744) );
  XOR2_X1 U811 ( .A(KEYINPUT38), .B(n744), .Z(n745) );
  NOR2_X1 U812 ( .A1(n746), .A2(n745), .ZN(n748) );
  NAND2_X1 U813 ( .A1(n883), .A2(G117), .ZN(n747) );
  NAND2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n876) );
  AND2_X1 U815 ( .A1(G1996), .A2(n876), .ZN(n749) );
  NOR2_X1 U816 ( .A1(n750), .A2(n749), .ZN(n939) );
  INV_X1 U817 ( .A(n770), .ZN(n751) );
  NOR2_X1 U818 ( .A1(n939), .A2(n751), .ZN(n761) );
  INV_X1 U819 ( .A(n761), .ZN(n752) );
  NAND2_X1 U820 ( .A1(n765), .A2(n752), .ZN(n753) );
  NOR2_X1 U821 ( .A1(n754), .A2(n753), .ZN(n756) );
  XNOR2_X1 U822 ( .A(G1986), .B(G290), .ZN(n995) );
  NAND2_X1 U823 ( .A1(n995), .A2(n770), .ZN(n755) );
  NAND2_X1 U824 ( .A1(n756), .A2(n755), .ZN(n773) );
  XOR2_X1 U825 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n757) );
  XNOR2_X1 U826 ( .A(KEYINPUT105), .B(n757), .ZN(n764) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n876), .ZN(n937) );
  NOR2_X1 U828 ( .A1(n891), .A2(G1991), .ZN(n758) );
  XNOR2_X1 U829 ( .A(n758), .B(KEYINPUT104), .ZN(n942) );
  NOR2_X1 U830 ( .A1(G1986), .A2(G290), .ZN(n759) );
  NOR2_X1 U831 ( .A1(n942), .A2(n759), .ZN(n760) );
  NOR2_X1 U832 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U833 ( .A1(n937), .A2(n762), .ZN(n763) );
  XNOR2_X1 U834 ( .A(n764), .B(n763), .ZN(n766) );
  NAND2_X1 U835 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U836 ( .A1(n767), .A2(n896), .ZN(n953) );
  NAND2_X1 U837 ( .A1(n768), .A2(n953), .ZN(n769) );
  XOR2_X1 U838 ( .A(KEYINPUT107), .B(n769), .Z(n771) );
  NAND2_X1 U839 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U840 ( .A1(n773), .A2(n772), .ZN(n775) );
  XNOR2_X1 U841 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n774) );
  XNOR2_X1 U842 ( .A(n775), .B(n774), .ZN(G329) );
  XOR2_X1 U843 ( .A(G2443), .B(G2446), .Z(n777) );
  XNOR2_X1 U844 ( .A(G2427), .B(G2451), .ZN(n776) );
  XNOR2_X1 U845 ( .A(n777), .B(n776), .ZN(n783) );
  XOR2_X1 U846 ( .A(G2430), .B(G2454), .Z(n779) );
  XNOR2_X1 U847 ( .A(G1341), .B(G1348), .ZN(n778) );
  XNOR2_X1 U848 ( .A(n779), .B(n778), .ZN(n781) );
  XOR2_X1 U849 ( .A(G2435), .B(G2438), .Z(n780) );
  XNOR2_X1 U850 ( .A(n781), .B(n780), .ZN(n782) );
  XOR2_X1 U851 ( .A(n783), .B(n782), .Z(n784) );
  AND2_X1 U852 ( .A1(G14), .A2(n784), .ZN(G401) );
  AND2_X1 U853 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U854 ( .A(G57), .ZN(G237) );
  INV_X1 U855 ( .A(G132), .ZN(G219) );
  INV_X1 U856 ( .A(G82), .ZN(G220) );
  XOR2_X1 U857 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n786) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n785) );
  XNOR2_X1 U859 ( .A(n786), .B(n785), .ZN(G223) );
  XOR2_X1 U860 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n788) );
  INV_X1 U861 ( .A(G223), .ZN(n850) );
  NAND2_X1 U862 ( .A1(G567), .A2(n850), .ZN(n787) );
  XNOR2_X1 U863 ( .A(n788), .B(n787), .ZN(G234) );
  INV_X1 U864 ( .A(G860), .ZN(n794) );
  OR2_X1 U865 ( .A1(n983), .A2(n794), .ZN(G153) );
  INV_X1 U866 ( .A(G171), .ZN(G301) );
  NAND2_X1 U867 ( .A1(G868), .A2(G301), .ZN(n790) );
  INV_X1 U868 ( .A(n903), .ZN(n988) );
  INV_X1 U869 ( .A(G868), .ZN(n834) );
  NAND2_X1 U870 ( .A1(n988), .A2(n834), .ZN(n789) );
  NAND2_X1 U871 ( .A1(n790), .A2(n789), .ZN(G284) );
  XNOR2_X1 U872 ( .A(KEYINPUT77), .B(G868), .ZN(n791) );
  NOR2_X1 U873 ( .A1(G286), .A2(n791), .ZN(n793) );
  NOR2_X1 U874 ( .A1(G868), .A2(G299), .ZN(n792) );
  NOR2_X1 U875 ( .A1(n793), .A2(n792), .ZN(G297) );
  NAND2_X1 U876 ( .A1(n794), .A2(G559), .ZN(n795) );
  NAND2_X1 U877 ( .A1(n795), .A2(n903), .ZN(n796) );
  XNOR2_X1 U878 ( .A(n796), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U879 ( .A1(G868), .A2(n983), .ZN(n797) );
  XOR2_X1 U880 ( .A(KEYINPUT78), .B(n797), .Z(n800) );
  NOR2_X1 U881 ( .A1(n988), .A2(G559), .ZN(n798) );
  NAND2_X1 U882 ( .A1(G868), .A2(n798), .ZN(n799) );
  NAND2_X1 U883 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U884 ( .A(KEYINPUT79), .B(n801), .ZN(G282) );
  NAND2_X1 U885 ( .A1(n882), .A2(G123), .ZN(n802) );
  XNOR2_X1 U886 ( .A(n802), .B(KEYINPUT18), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G111), .A2(n883), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U889 ( .A1(G135), .A2(n722), .ZN(n806) );
  NAND2_X1 U890 ( .A1(G99), .A2(n879), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U892 ( .A1(n808), .A2(n807), .ZN(n941) );
  XNOR2_X1 U893 ( .A(n941), .B(G2096), .ZN(n809) );
  XNOR2_X1 U894 ( .A(n809), .B(KEYINPUT80), .ZN(n811) );
  INV_X1 U895 ( .A(G2100), .ZN(n810) );
  NAND2_X1 U896 ( .A1(n811), .A2(n810), .ZN(G156) );
  NAND2_X1 U897 ( .A1(n812), .A2(G55), .ZN(n813) );
  XNOR2_X1 U898 ( .A(n813), .B(KEYINPUT82), .ZN(n822) );
  NAND2_X1 U899 ( .A1(G80), .A2(n604), .ZN(n816) );
  NAND2_X1 U900 ( .A1(G93), .A2(n814), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n816), .A2(n815), .ZN(n820) );
  NAND2_X1 U902 ( .A1(G67), .A2(n817), .ZN(n818) );
  XNOR2_X1 U903 ( .A(KEYINPUT81), .B(n818), .ZN(n819) );
  NOR2_X1 U904 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U905 ( .A1(n822), .A2(n821), .ZN(n835) );
  NAND2_X1 U906 ( .A1(n903), .A2(G559), .ZN(n832) );
  XNOR2_X1 U907 ( .A(n983), .B(n832), .ZN(n823) );
  NOR2_X1 U908 ( .A1(G860), .A2(n823), .ZN(n824) );
  XOR2_X1 U909 ( .A(n835), .B(n824), .Z(G145) );
  XNOR2_X1 U910 ( .A(KEYINPUT87), .B(G290), .ZN(n825) );
  XNOR2_X1 U911 ( .A(n825), .B(G305), .ZN(n826) );
  XNOR2_X1 U912 ( .A(KEYINPUT19), .B(n826), .ZN(n828) );
  XNOR2_X1 U913 ( .A(G299), .B(G166), .ZN(n827) );
  XNOR2_X1 U914 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U915 ( .A(n829), .B(G288), .ZN(n830) );
  XNOR2_X1 U916 ( .A(n830), .B(n835), .ZN(n831) );
  XNOR2_X1 U917 ( .A(n831), .B(n983), .ZN(n900) );
  XOR2_X1 U918 ( .A(n900), .B(n832), .Z(n833) );
  NAND2_X1 U919 ( .A1(G868), .A2(n833), .ZN(n837) );
  NAND2_X1 U920 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U921 ( .A1(n837), .A2(n836), .ZN(G295) );
  NAND2_X1 U922 ( .A1(G2078), .A2(G2084), .ZN(n838) );
  XOR2_X1 U923 ( .A(KEYINPUT20), .B(n838), .Z(n839) );
  NAND2_X1 U924 ( .A1(G2090), .A2(n839), .ZN(n840) );
  XNOR2_X1 U925 ( .A(KEYINPUT21), .B(n840), .ZN(n841) );
  NAND2_X1 U926 ( .A1(n841), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U927 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U928 ( .A1(G220), .A2(G219), .ZN(n842) );
  XOR2_X1 U929 ( .A(KEYINPUT22), .B(n842), .Z(n843) );
  NOR2_X1 U930 ( .A1(G218), .A2(n843), .ZN(n844) );
  NAND2_X1 U931 ( .A1(G96), .A2(n844), .ZN(n856) );
  NAND2_X1 U932 ( .A1(n856), .A2(G2106), .ZN(n848) );
  NAND2_X1 U933 ( .A1(G69), .A2(G120), .ZN(n845) );
  NOR2_X1 U934 ( .A1(G237), .A2(n845), .ZN(n846) );
  NAND2_X1 U935 ( .A1(G108), .A2(n846), .ZN(n857) );
  NAND2_X1 U936 ( .A1(n857), .A2(G567), .ZN(n847) );
  NAND2_X1 U937 ( .A1(n848), .A2(n847), .ZN(n931) );
  NAND2_X1 U938 ( .A1(G483), .A2(G661), .ZN(n849) );
  NOR2_X1 U939 ( .A1(n931), .A2(n849), .ZN(n855) );
  NAND2_X1 U940 ( .A1(n855), .A2(G36), .ZN(G176) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n850), .ZN(G217) );
  NAND2_X1 U942 ( .A1(G15), .A2(G2), .ZN(n851) );
  XNOR2_X1 U943 ( .A(KEYINPUT109), .B(n851), .ZN(n852) );
  NAND2_X1 U944 ( .A1(n852), .A2(G661), .ZN(n853) );
  XNOR2_X1 U945 ( .A(KEYINPUT110), .B(n853), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n854) );
  NAND2_X1 U947 ( .A1(n855), .A2(n854), .ZN(G188) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G96), .ZN(G221) );
  INV_X1 U951 ( .A(G69), .ZN(G235) );
  NOR2_X1 U952 ( .A1(n857), .A2(n856), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  NAND2_X1 U954 ( .A1(G100), .A2(n879), .ZN(n859) );
  NAND2_X1 U955 ( .A1(G112), .A2(n883), .ZN(n858) );
  NAND2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U957 ( .A1(n882), .A2(G124), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U959 ( .A1(G136), .A2(n722), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(KEYINPUT113), .B(n863), .Z(n864) );
  NOR2_X1 U962 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U963 ( .A1(G130), .A2(n882), .ZN(n867) );
  NAND2_X1 U964 ( .A1(G118), .A2(n883), .ZN(n866) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U966 ( .A1(G142), .A2(n722), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G106), .A2(n879), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(KEYINPUT45), .B(n870), .Z(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n895) );
  XOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n874) );
  XNOR2_X1 U972 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U974 ( .A(n875), .B(n941), .Z(n878) );
  XOR2_X1 U975 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n890) );
  NAND2_X1 U977 ( .A1(G139), .A2(n722), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G103), .A2(n879), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n889) );
  NAND2_X1 U980 ( .A1(G127), .A2(n882), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G115), .A2(n883), .ZN(n884) );
  NAND2_X1 U982 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n886), .Z(n887) );
  XNOR2_X1 U984 ( .A(KEYINPUT114), .B(n887), .ZN(n888) );
  NOR2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n932) );
  XOR2_X1 U986 ( .A(n890), .B(n932), .Z(n893) );
  XOR2_X1 U987 ( .A(G160), .B(n891), .Z(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n896), .B(G162), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U992 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U993 ( .A(KEYINPUT117), .B(n900), .Z(n902) );
  XNOR2_X1 U994 ( .A(G171), .B(G286), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n902), .B(n901), .ZN(n904) );
  XNOR2_X1 U996 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U997 ( .A1(G37), .A2(n905), .ZN(G397) );
  XOR2_X1 U998 ( .A(KEYINPUT43), .B(G2678), .Z(n907) );
  XNOR2_X1 U999 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1001 ( .A(KEYINPUT42), .B(G2090), .Z(n909) );
  XNOR2_X1 U1002 ( .A(G2067), .B(G2072), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1004 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1005 ( .A(G2096), .B(G2100), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n913), .B(n912), .ZN(n915) );
  XOR2_X1 U1007 ( .A(G2078), .B(G2084), .Z(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(G227) );
  XOR2_X1 U1009 ( .A(G1976), .B(G1971), .Z(n917) );
  XNOR2_X1 U1010 ( .A(G1981), .B(G1966), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1012 ( .A(n918), .B(KEYINPUT41), .Z(n920) );
  XNOR2_X1 U1013 ( .A(G1996), .B(G1991), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n920), .B(n919), .ZN(n924) );
  XOR2_X1 U1015 ( .A(G2474), .B(G1961), .Z(n922) );
  XNOR2_X1 U1016 ( .A(G1986), .B(G1956), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(n924), .B(n923), .ZN(G229) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n931), .ZN(n928) );
  NOR2_X1 U1020 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1022 ( .A1(G397), .A2(n926), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(G395), .A2(n929), .ZN(n930) );
  XOR2_X1 U1025 ( .A(KEYINPUT118), .B(n930), .Z(G225) );
  XNOR2_X1 U1026 ( .A(KEYINPUT119), .B(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(n931), .ZN(G319) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1029 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1030 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT50), .B(n935), .Z(n952) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n938), .Z(n947) );
  XNOR2_X1 U1036 ( .A(G160), .B(G2084), .ZN(n940) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n945) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT120), .B(n943), .Z(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT121), .B(n950), .ZN(n951) );
  NOR2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n954) );
  NAND2_X1 U1045 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n955), .ZN(n956) );
  NAND2_X1 U1047 ( .A1(n956), .A2(G29), .ZN(n1032) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G33), .B(G2072), .ZN(n957) );
  NOR2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n966) );
  XNOR2_X1 U1051 ( .A(G32), .B(n959), .ZN(n960) );
  NAND2_X1 U1052 ( .A1(n960), .A2(G28), .ZN(n964) );
  XOR2_X1 U1053 ( .A(G27), .B(n961), .Z(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT122), .B(n962), .ZN(n963) );
  NOR2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(G25), .B(G1991), .ZN(n967) );
  NOR2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1059 ( .A(KEYINPUT53), .B(n969), .Z(n972) );
  XOR2_X1 U1060 ( .A(G34), .B(KEYINPUT54), .Z(n970) );
  XNOR2_X1 U1061 ( .A(G2084), .B(n970), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G35), .B(G2090), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1065 ( .A(KEYINPUT123), .B(n975), .Z(n976) );
  NOR2_X1 U1066 ( .A1(G29), .A2(n976), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(KEYINPUT55), .B(n977), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n978), .A2(G11), .ZN(n1030) );
  XNOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .ZN(n1003) );
  XOR2_X1 U1070 ( .A(G168), .B(G1966), .Z(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1072 ( .A(KEYINPUT57), .B(n981), .Z(n1001) );
  XNOR2_X1 U1073 ( .A(G299), .B(G1956), .ZN(n985) );
  XOR2_X1 U1074 ( .A(G1341), .B(KEYINPUT125), .Z(n982) );
  XNOR2_X1 U1075 ( .A(n983), .B(n982), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n999) );
  XNOR2_X1 U1078 ( .A(n988), .B(G1348), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G301), .B(G1961), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT124), .B(n991), .ZN(n997) );
  NAND2_X1 U1082 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1028) );
  INV_X1 U1089 ( .A(G16), .ZN(n1026) );
  XOR2_X1 U1090 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n1024) );
  XOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .Z(n1004) );
  XNOR2_X1 U1092 ( .A(G4), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(G20), .B(G1956), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(KEYINPUT60), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G23), .B(G1976), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(G1986), .B(G24), .Z(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G1966), .B(G21), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(G5), .B(G1961), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(n1024), .B(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1114 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(n1033), .B(KEYINPUT62), .ZN(n1034) );
  XNOR2_X1 U1117 ( .A(KEYINPUT127), .B(n1034), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

