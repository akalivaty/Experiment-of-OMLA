

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  XNOR2_X1 U320 ( .A(n300), .B(n299), .ZN(n305) );
  XOR2_X1 U321 ( .A(n334), .B(n418), .Z(n288) );
  XOR2_X1 U322 ( .A(G148GAT), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U323 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n296) );
  INV_X1 U324 ( .A(KEYINPUT32), .ZN(n371) );
  XNOR2_X1 U325 ( .A(n372), .B(n371), .ZN(n373) );
  NOR2_X1 U326 ( .A1(n577), .A2(n478), .ZN(n479) );
  XNOR2_X1 U327 ( .A(n295), .B(n294), .ZN(n300) );
  XNOR2_X1 U328 ( .A(n374), .B(n373), .ZN(n376) );
  NAND2_X1 U329 ( .A1(n462), .A2(n461), .ZN(n475) );
  XNOR2_X1 U330 ( .A(KEYINPUT104), .B(n483), .ZN(n490) );
  XNOR2_X1 U331 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U332 ( .A(n447), .B(n446), .ZN(G1349GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT22), .B(G106GAT), .Z(n290) );
  XOR2_X1 U334 ( .A(G141GAT), .B(G22GAT), .Z(n385) );
  XNOR2_X1 U335 ( .A(n385), .B(n363), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U337 ( .A(n291), .B(G218GAT), .Z(n295) );
  XOR2_X1 U338 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n293) );
  XNOR2_X1 U339 ( .A(KEYINPUT24), .B(KEYINPUT87), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U341 ( .A(KEYINPUT73), .B(G162GAT), .Z(n334) );
  XNOR2_X1 U342 ( .A(n296), .B(KEYINPUT2), .ZN(n418) );
  NAND2_X1 U343 ( .A1(G228GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n288), .B(n297), .ZN(n298) );
  XNOR2_X1 U345 ( .A(G50GAT), .B(n298), .ZN(n299) );
  XOR2_X1 U346 ( .A(KEYINPUT88), .B(G204GAT), .Z(n302) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(G211GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n304) );
  XOR2_X1 U349 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n303) );
  XOR2_X1 U350 ( .A(n304), .B(n303), .Z(n311) );
  XOR2_X1 U351 ( .A(n305), .B(n311), .Z(n454) );
  XOR2_X1 U352 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n307) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G8GAT), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n307), .B(n306), .ZN(n309) );
  XOR2_X1 U355 ( .A(G36GAT), .B(G92GAT), .Z(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n315) );
  XOR2_X1 U357 ( .A(G64GAT), .B(KEYINPUT77), .Z(n313) );
  XNOR2_X1 U358 ( .A(G190GAT), .B(G218GAT), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n310), .B(KEYINPUT75), .ZN(n338) );
  XNOR2_X1 U360 ( .A(n311), .B(n338), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n317) );
  NAND2_X1 U363 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n323) );
  XNOR2_X1 U365 ( .A(G183GAT), .B(KEYINPUT83), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n318), .B(G176GAT), .ZN(n319) );
  XOR2_X1 U367 ( .A(n319), .B(KEYINPUT17), .Z(n321) );
  XNOR2_X1 U368 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n320) );
  XOR2_X1 U369 ( .A(n321), .B(n320), .Z(n442) );
  INV_X1 U370 ( .A(n442), .ZN(n322) );
  XOR2_X2 U371 ( .A(n323), .B(n322), .Z(n511) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n324), .B(G29GAT), .ZN(n325) );
  XOR2_X1 U374 ( .A(n325), .B(KEYINPUT7), .Z(n327) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(G50GAT), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n389) );
  XOR2_X1 U377 ( .A(KEYINPUT71), .B(G92GAT), .Z(n329) );
  XNOR2_X1 U378 ( .A(G99GAT), .B(G85GAT), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(n330), .ZN(n375) );
  XOR2_X1 U381 ( .A(n389), .B(n375), .Z(n342) );
  XOR2_X1 U382 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n332) );
  XNOR2_X1 U383 ( .A(G134GAT), .B(KEYINPUT74), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n334), .B(n333), .Z(n336) );
  NAND2_X1 U386 ( .A1(G232GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U388 ( .A(n337), .B(KEYINPUT9), .Z(n340) );
  XNOR2_X1 U389 ( .A(n338), .B(KEYINPUT10), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U391 ( .A(n342), .B(n341), .ZN(n552) );
  XOR2_X1 U392 ( .A(G78GAT), .B(G155GAT), .Z(n344) );
  XNOR2_X1 U393 ( .A(G15GAT), .B(G183GAT), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U395 ( .A(n345), .B(G211GAT), .Z(n347) );
  XOR2_X1 U396 ( .A(G1GAT), .B(G8GAT), .Z(n384) );
  XNOR2_X1 U397 ( .A(G22GAT), .B(n384), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n352) );
  XNOR2_X1 U399 ( .A(G57GAT), .B(G64GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n348), .B(KEYINPUT13), .ZN(n370) );
  XOR2_X1 U401 ( .A(n370), .B(KEYINPUT12), .Z(n350) );
  NAND2_X1 U402 ( .A1(G231GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U404 ( .A(n352), .B(n351), .Z(n360) );
  XOR2_X1 U405 ( .A(KEYINPUT80), .B(KEYINPUT77), .Z(n354) );
  XNOR2_X1 U406 ( .A(G127GAT), .B(G71GAT), .ZN(n353) );
  XNOR2_X1 U407 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U408 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n356) );
  XNOR2_X1 U409 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U412 ( .A(n360), .B(n359), .Z(n474) );
  INV_X1 U413 ( .A(n474), .ZN(n571) );
  XOR2_X1 U414 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n391) );
  XOR2_X1 U415 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n362) );
  XNOR2_X1 U416 ( .A(KEYINPUT69), .B(KEYINPUT31), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n367) );
  XOR2_X1 U418 ( .A(n363), .B(G204GAT), .Z(n365) );
  XOR2_X1 U419 ( .A(G120GAT), .B(G71GAT), .Z(n430) );
  XNOR2_X1 U420 ( .A(G176GAT), .B(n430), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U422 ( .A(n367), .B(n366), .Z(n369) );
  NAND2_X1 U423 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n374) );
  XNOR2_X1 U425 ( .A(n370), .B(KEYINPUT70), .ZN(n372) );
  XNOR2_X1 U426 ( .A(n376), .B(n375), .ZN(n448) );
  XNOR2_X1 U427 ( .A(n448), .B(KEYINPUT41), .ZN(n542) );
  XNOR2_X1 U428 ( .A(G169GAT), .B(G15GAT), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n377), .B(G113GAT), .ZN(n438) );
  XOR2_X1 U430 ( .A(n438), .B(KEYINPUT67), .Z(n379) );
  NAND2_X1 U431 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U432 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U433 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n381) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U436 ( .A(n383), .B(n382), .Z(n387) );
  XNOR2_X1 U437 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U438 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U439 ( .A(n389), .B(n388), .Z(n493) );
  INV_X1 U440 ( .A(n493), .ZN(n564) );
  NAND2_X1 U441 ( .A1(n542), .A2(n564), .ZN(n390) );
  XOR2_X1 U442 ( .A(n391), .B(n390), .Z(n392) );
  NOR2_X1 U443 ( .A1(n571), .A2(n392), .ZN(n393) );
  NAND2_X1 U444 ( .A1(n552), .A2(n393), .ZN(n394) );
  XNOR2_X1 U445 ( .A(n394), .B(KEYINPUT47), .ZN(n400) );
  XNOR2_X1 U446 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n395) );
  XOR2_X1 U447 ( .A(KEYINPUT76), .B(n552), .Z(n558) );
  XOR2_X1 U448 ( .A(n395), .B(n558), .Z(n577) );
  NOR2_X1 U449 ( .A1(n577), .A2(n474), .ZN(n396) );
  XNOR2_X1 U450 ( .A(KEYINPUT45), .B(n396), .ZN(n397) );
  NAND2_X1 U451 ( .A1(n397), .A2(n448), .ZN(n398) );
  XOR2_X1 U452 ( .A(KEYINPUT68), .B(n493), .Z(n555) );
  NOR2_X1 U453 ( .A1(n398), .A2(n555), .ZN(n399) );
  NOR2_X1 U454 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U455 ( .A(KEYINPUT48), .B(n401), .ZN(n520) );
  NOR2_X1 U456 ( .A1(n511), .A2(n520), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n402), .B(KEYINPUT54), .ZN(n425) );
  XOR2_X1 U458 ( .A(KEYINPUT1), .B(G120GAT), .Z(n404) );
  XNOR2_X1 U459 ( .A(G141GAT), .B(G113GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U461 ( .A(KEYINPUT5), .B(G57GAT), .Z(n406) );
  XNOR2_X1 U462 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U464 ( .A(n408), .B(n407), .Z(n415) );
  XOR2_X1 U465 ( .A(G127GAT), .B(KEYINPUT81), .Z(n410) );
  XNOR2_X1 U466 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n437) );
  XOR2_X1 U468 ( .A(G85GAT), .B(G148GAT), .Z(n412) );
  XNOR2_X1 U469 ( .A(G29GAT), .B(G162GAT), .ZN(n411) );
  XNOR2_X1 U470 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n437), .B(n413), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n424) );
  XOR2_X1 U473 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n417) );
  XNOR2_X1 U474 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U476 ( .A(n418), .B(G1GAT), .Z(n420) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n508) );
  NAND2_X1 U481 ( .A1(n425), .A2(n508), .ZN(n563) );
  NOR2_X1 U482 ( .A1(n454), .A2(n563), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n426), .B(KEYINPUT55), .ZN(n443) );
  XOR2_X1 U484 ( .A(KEYINPUT84), .B(G99GAT), .Z(n428) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G190GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT64), .Z(n434) );
  XNOR2_X1 U491 ( .A(KEYINPUT82), .B(KEYINPUT85), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U494 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X2 U496 ( .A(n442), .B(n441), .Z(n522) );
  NOR2_X2 U497 ( .A1(n443), .A2(n522), .ZN(n559) );
  NAND2_X1 U498 ( .A1(n559), .A2(n542), .ZN(n447) );
  XOR2_X1 U499 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n445) );
  XNOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n444) );
  NAND2_X1 U501 ( .A1(n555), .A2(n448), .ZN(n480) );
  NOR2_X1 U502 ( .A1(n558), .A2(n474), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n449), .B(KEYINPUT16), .ZN(n463) );
  XNOR2_X1 U504 ( .A(n511), .B(KEYINPUT27), .ZN(n457) );
  NOR2_X1 U505 ( .A1(n508), .A2(n457), .ZN(n538) );
  XOR2_X1 U506 ( .A(KEYINPUT28), .B(n454), .Z(n516) );
  NAND2_X1 U507 ( .A1(n538), .A2(n516), .ZN(n521) );
  XNOR2_X1 U508 ( .A(n521), .B(KEYINPUT97), .ZN(n451) );
  XNOR2_X1 U509 ( .A(n522), .B(KEYINPUT86), .ZN(n450) );
  NAND2_X1 U510 ( .A1(n451), .A2(n450), .ZN(n462) );
  NOR2_X1 U511 ( .A1(n511), .A2(n522), .ZN(n452) );
  NOR2_X1 U512 ( .A1(n454), .A2(n452), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n453), .B(KEYINPUT25), .ZN(n459) );
  XOR2_X1 U514 ( .A(KEYINPUT98), .B(KEYINPUT26), .Z(n456) );
  NAND2_X1 U515 ( .A1(n454), .A2(n522), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(n455), .ZN(n537) );
  INV_X1 U517 ( .A(n537), .ZN(n562) );
  OR2_X1 U518 ( .A1(n562), .A2(n457), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n459), .A2(n458), .ZN(n460) );
  NAND2_X1 U520 ( .A1(n508), .A2(n460), .ZN(n461) );
  NAND2_X1 U521 ( .A1(n463), .A2(n475), .ZN(n494) );
  NOR2_X1 U522 ( .A1(n480), .A2(n494), .ZN(n464) );
  XNOR2_X1 U523 ( .A(KEYINPUT99), .B(n464), .ZN(n472) );
  NOR2_X1 U524 ( .A1(n508), .A2(n472), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT34), .B(KEYINPUT100), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U527 ( .A(G1GAT), .B(n467), .Z(G1324GAT) );
  NOR2_X1 U528 ( .A1(n511), .A2(n472), .ZN(n468) );
  XOR2_X1 U529 ( .A(G8GAT), .B(n468), .Z(G1325GAT) );
  NOR2_X1 U530 ( .A1(n522), .A2(n472), .ZN(n470) );
  XNOR2_X1 U531 ( .A(KEYINPUT101), .B(KEYINPUT35), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n470), .B(n469), .ZN(n471) );
  XOR2_X1 U533 ( .A(G15GAT), .B(n471), .Z(G1326GAT) );
  NOR2_X1 U534 ( .A1(n516), .A2(n472), .ZN(n473) );
  XOR2_X1 U535 ( .A(G22GAT), .B(n473), .Z(G1327GAT) );
  INV_X1 U536 ( .A(KEYINPUT38), .ZN(n482) );
  INV_X1 U537 ( .A(KEYINPUT103), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U540 ( .A(KEYINPUT37), .B(n479), .ZN(n505) );
  NOR2_X1 U541 ( .A1(n505), .A2(n480), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n508), .A2(n490), .ZN(n485) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  NOR2_X1 U546 ( .A1(n511), .A2(n490), .ZN(n486) );
  XOR2_X1 U547 ( .A(G36GAT), .B(n486), .Z(G1329GAT) );
  NOR2_X1 U548 ( .A1(n522), .A2(n490), .ZN(n488) );
  INV_X1 U549 ( .A(KEYINPUT40), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NOR2_X1 U552 ( .A1(n516), .A2(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(G1331GAT) );
  NAND2_X1 U555 ( .A1(n493), .A2(n542), .ZN(n506) );
  OR2_X1 U556 ( .A1(n506), .A2(n494), .ZN(n502) );
  NOR2_X1 U557 ( .A1(n508), .A2(n502), .ZN(n495) );
  XOR2_X1 U558 ( .A(n495), .B(KEYINPUT42), .Z(n496) );
  XNOR2_X1 U559 ( .A(G57GAT), .B(n496), .ZN(G1332GAT) );
  NOR2_X1 U560 ( .A1(n511), .A2(n502), .ZN(n497) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(n497), .Z(n498) );
  XNOR2_X1 U562 ( .A(G64GAT), .B(n498), .ZN(G1333GAT) );
  NOR2_X1 U563 ( .A1(n522), .A2(n502), .ZN(n500) );
  XNOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U566 ( .A(G71GAT), .B(n501), .ZN(G1334GAT) );
  NOR2_X1 U567 ( .A1(n516), .A2(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NOR2_X1 U570 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n507), .B(KEYINPUT109), .ZN(n515) );
  NOR2_X1 U572 ( .A1(n508), .A2(n515), .ZN(n509) );
  XOR2_X1 U573 ( .A(n509), .B(KEYINPUT110), .Z(n510) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NOR2_X1 U575 ( .A1(n511), .A2(n515), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(G1337GAT) );
  NOR2_X1 U578 ( .A1(n522), .A2(n515), .ZN(n514) );
  XOR2_X1 U579 ( .A(G99GAT), .B(n514), .Z(G1338GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U581 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U583 ( .A(G106GAT), .B(n519), .Z(G1339GAT) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n525) );
  OR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U586 ( .A1(n520), .A2(n523), .ZN(n534) );
  NAND2_X1 U587 ( .A1(n555), .A2(n534), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n527) );
  NAND2_X1 U590 ( .A1(n534), .A2(n542), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n529) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT115), .Z(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  XNOR2_X1 U594 ( .A(G127GAT), .B(KEYINPUT118), .ZN(n533) );
  XOR2_X1 U595 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n531) );
  NAND2_X1 U596 ( .A1(n534), .A2(n571), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(G134GAT), .B(KEYINPUT51), .Z(n536) );
  NAND2_X1 U600 ( .A1(n534), .A2(n558), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  XOR2_X1 U602 ( .A(G141GAT), .B(KEYINPUT119), .Z(n541) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n520), .A2(n539), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n550), .A2(n564), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(G1344GAT) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n544) );
  NAND2_X1 U609 ( .A1(n550), .A2(n542), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n548) );
  NAND2_X1 U613 ( .A1(n550), .A2(n571), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G155GAT), .B(n549), .ZN(G1346GAT) );
  INV_X1 U616 ( .A(n550), .ZN(n551) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U618 ( .A(G162GAT), .B(KEYINPUT123), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n559), .A2(n555), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U622 ( .A1(n559), .A2(n571), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n560), .B(KEYINPUT58), .ZN(n561) );
  XNOR2_X1 U626 ( .A(G190GAT), .B(n561), .ZN(G1351GAT) );
  XOR2_X1 U627 ( .A(G197GAT), .B(KEYINPUT60), .Z(n566) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n572), .A2(n564), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .Z(n570) );
  INV_X1 U634 ( .A(n572), .ZN(n576) );
  OR2_X1 U635 ( .A1(n576), .A2(n448), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n575) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n579) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(n579), .B(n578), .Z(G1355GAT) );
endmodule

