//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n204), .B1(KEYINPUT80), .B2(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(KEYINPUT80), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G57gat), .B(G64gat), .Z(new_n209));
  OR2_X1    g008(.A1(new_n209), .A2(KEYINPUT86), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(KEYINPUT86), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT9), .A3(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(G71gat), .A2(G78gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT85), .ZN(new_n214));
  INV_X1    g013(.A(G71gat), .ZN(new_n215));
  INV_X1    g014(.A(G78gat), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n212), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(KEYINPUT9), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n215), .B2(new_n216), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n209), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT87), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n208), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(KEYINPUT88), .ZN(new_n225));
  INV_X1    g024(.A(new_n222), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT21), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n225), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G183gat), .B(G211gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT89), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n228), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G155gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(G231gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n234), .B(new_n235), .Z(new_n236));
  OR2_X1    g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n236), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G190gat), .B(G218gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(G85gat), .A2(G92gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT7), .ZN(new_n243));
  INV_X1    g042(.A(G99gat), .ZN(new_n244));
  INV_X1    g043(.A(G106gat), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT8), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n243), .B(new_n246), .C1(G85gat), .C2(G92gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(G99gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT90), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G43gat), .B(G50gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(KEYINPUT15), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT79), .B(G29gat), .ZN(new_n254));
  INV_X1    g053(.A(G36gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(G29gat), .A2(G36gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT14), .ZN(new_n258));
  NOR3_X1   g057(.A1(new_n253), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(KEYINPUT15), .ZN(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n260), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT81), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT17), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n264), .A2(KEYINPUT17), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n263), .A2(new_n266), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n251), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n250), .A2(new_n263), .B1(KEYINPUT41), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n241), .B1(new_n272), .B2(KEYINPUT91), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(KEYINPUT91), .B2(new_n272), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n269), .A2(new_n275), .A3(new_n271), .A4(new_n241), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n270), .A2(KEYINPUT41), .ZN(new_n277));
  XNOR2_X1  g076(.A(G134gat), .B(G162gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT92), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n274), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n279), .A2(KEYINPUT92), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(new_n274), .B2(new_n276), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n240), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n222), .B(new_n249), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT10), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n250), .A2(KEYINPUT10), .A3(new_n226), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G230gat), .A2(G233gat), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(KEYINPUT93), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n290), .A2(KEYINPUT95), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT95), .B1(new_n290), .B2(new_n293), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n286), .A2(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT94), .B(G120gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n299), .B(G148gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(G176gat), .B(G204gat), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n300), .B(new_n301), .Z(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n290), .A2(new_n293), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n297), .A3(new_n302), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n285), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n263), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(new_n208), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT83), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n208), .B1(new_n267), .B2(new_n268), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT82), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(KEYINPUT82), .B(new_n208), .C1(new_n267), .C2(new_n268), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n311), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT84), .ZN(new_n317));
  NAND2_X1  g116(.A1(G229gat), .A2(G233gat), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n316), .A2(new_n317), .A3(KEYINPUT18), .A4(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n311), .A2(new_n314), .A3(new_n318), .A4(new_n315), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT18), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n309), .A2(new_n208), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n318), .B(KEYINPUT13), .Z(new_n324));
  AOI22_X1  g123(.A1(new_n320), .A2(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT84), .B1(new_n320), .B2(new_n321), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n319), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G113gat), .B(G141gat), .ZN(new_n328));
  INV_X1    g127(.A(G197gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT11), .B(G169gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n332), .B(KEYINPUT12), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n333), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n319), .A2(new_n325), .A3(new_n326), .A4(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT31), .B(G50gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  OR3_X1    g140(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(KEYINPUT73), .B(KEYINPUT2), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n348));
  INV_X1    g147(.A(G155gat), .ZN(new_n349));
  INV_X1    g148(.A(G162gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT72), .B1(G155gat), .B2(G162gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n341), .ZN(new_n353));
  NOR3_X1   g152(.A1(new_n346), .A2(new_n347), .A3(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n351), .A2(new_n352), .A3(new_n341), .ZN(new_n355));
  OR2_X1    g154(.A1(KEYINPUT73), .A2(KEYINPUT2), .ZN(new_n356));
  NAND2_X1  g155(.A1(KEYINPUT73), .A2(KEYINPUT2), .ZN(new_n357));
  INV_X1    g156(.A(G141gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G148gat), .ZN(new_n359));
  INV_X1    g158(.A(G148gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(G141gat), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n356), .B(new_n357), .C1(new_n359), .C2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT74), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n344), .B1(new_n354), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT71), .B(KEYINPUT29), .Z(new_n365));
  OR2_X1    g164(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n366));
  NAND2_X1  g165(.A1(G211gat), .A2(G218gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G211gat), .B(G218gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n369), .A2(new_n372), .A3(new_n370), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n365), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n376), .A2(KEYINPUT75), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n376), .B2(KEYINPUT75), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n364), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n374), .A2(new_n375), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n378), .B(new_n344), .C1(new_n354), .C2(new_n363), .ZN(new_n382));
  INV_X1    g181(.A(new_n365), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n380), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G22gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT3), .B1(new_n381), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n347), .B1(new_n346), .B2(new_n353), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n355), .A2(new_n362), .A3(KEYINPUT74), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n343), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(G228gat), .B(G233gat), .C1(new_n384), .C2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n387), .A2(new_n390), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n390), .B1(new_n387), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n339), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n338), .A3(new_n398), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G15gat), .B(G43gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G71gat), .B(G99gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n408), .B(KEYINPUT64), .Z(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g209(.A1(G169gat), .A2(G176gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT26), .ZN(new_n412));
  NAND2_X1  g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(G169gat), .A2(G176gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n412), .B(new_n413), .C1(new_n416), .C2(new_n411), .ZN(new_n417));
  INV_X1    g216(.A(G183gat), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT66), .B1(new_n418), .B2(KEYINPUT27), .ZN(new_n419));
  AOI21_X1  g218(.A(G190gat), .B1(new_n418), .B2(KEYINPUT27), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(G183gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n420), .A2(new_n419), .A3(new_n423), .A4(KEYINPUT67), .ZN(new_n427));
  XOR2_X1   g226(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n430), .B1(new_n422), .B2(G183gat), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT69), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n431), .A2(new_n432), .A3(new_n420), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n432), .B1(new_n431), .B2(new_n420), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n417), .B1(new_n429), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(G134gat), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(G127gat), .ZN(new_n438));
  INV_X1    g237(.A(G127gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(G134gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G113gat), .B(G120gat), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(KEYINPUT1), .ZN(new_n443));
  INV_X1    g242(.A(G120gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(G113gat), .ZN(new_n445));
  INV_X1    g244(.A(G113gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(G120gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G127gat), .B(G134gat), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT1), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n411), .A2(KEYINPUT23), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT23), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(G169gat), .B2(G176gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n414), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n459));
  INV_X1    g258(.A(G190gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n418), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(KEYINPUT24), .A3(new_n413), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT24), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n463), .A2(G183gat), .A3(G190gat), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n458), .A2(new_n459), .A3(new_n462), .A4(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT65), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n413), .A2(new_n466), .A3(new_n463), .ZN(new_n467));
  OAI211_X1 g266(.A(G183gat), .B(G190gat), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n467), .A2(new_n468), .A3(new_n461), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT25), .B1(new_n469), .B2(new_n457), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  OR3_X1    g270(.A1(new_n436), .A2(new_n453), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n453), .B1(new_n436), .B2(new_n471), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n410), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n407), .B1(new_n474), .B2(KEYINPUT33), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n410), .A3(new_n473), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT34), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n472), .A2(new_n479), .A3(new_n410), .A4(new_n473), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT32), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n478), .B(new_n480), .C1(new_n482), .C2(new_n474), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n476), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n383), .B1(new_n436), .B2(new_n471), .ZN(new_n488));
  NAND2_X1  g287(.A1(G226gat), .A2(G233gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n381), .ZN(new_n491));
  OAI211_X1 g290(.A(G226gat), .B(G233gat), .C1(new_n436), .C2(new_n471), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n391), .B1(new_n436), .B2(new_n471), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n489), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(new_n492), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT30), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n492), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n381), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G8gat), .B(G36gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(G64gat), .B(G92gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n497), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT30), .B(new_n505), .C1(new_n493), .C2(new_n496), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n484), .A2(new_n476), .A3(new_n485), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n404), .A2(new_n487), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G1gat), .B(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(G85gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT0), .B(G57gat), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n515), .B(new_n516), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT5), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n452), .B1(new_n395), .B2(new_n378), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n364), .A2(KEYINPUT3), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n344), .B(new_n452), .C1(new_n354), .C2(new_n363), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT4), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n395), .A2(new_n525), .A3(new_n452), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G225gat), .A2(G233gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n364), .A2(new_n453), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n528), .B1(new_n530), .B2(new_n523), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n519), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n521), .A2(new_n520), .B1(new_n524), .B2(new_n526), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT5), .B1(new_n534), .B2(new_n528), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n518), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n519), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n531), .B1(new_n534), .B2(new_n528), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n517), .B(new_n537), .C1(new_n538), .C2(new_n519), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n533), .A2(new_n535), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT6), .A3(new_n517), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n512), .A2(KEYINPUT35), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n487), .A2(KEYINPUT78), .A3(new_n510), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT78), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n484), .A2(new_n476), .A3(new_n485), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(new_n486), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n541), .A2(new_n543), .B1(new_n508), .B2(new_n507), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n546), .A2(new_n549), .A3(new_n550), .A4(new_n404), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT37), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n493), .A2(new_n496), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT37), .B1(new_n499), .B2(new_n501), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT38), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n541), .A2(new_n543), .A3(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT77), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n495), .A2(new_n491), .A3(new_n492), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(KEYINPUT37), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n490), .A2(new_n492), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n381), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n566), .A2(KEYINPUT77), .A3(KEYINPUT37), .A4(new_n561), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT38), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n555), .B1(new_n493), .B2(new_n496), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n564), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n505), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n493), .A2(new_n496), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n505), .A2(KEYINPUT38), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n401), .A2(new_n403), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n530), .A2(new_n578), .A3(new_n528), .A4(new_n523), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n579), .A2(KEYINPUT39), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n530), .A2(new_n528), .A3(new_n523), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n580), .B(new_n582), .C1(new_n528), .C2(new_n534), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n528), .B1(new_n522), .B2(new_n527), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n517), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(KEYINPUT40), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n539), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT40), .B1(new_n583), .B2(new_n586), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n509), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n577), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n487), .A2(KEYINPUT36), .A3(new_n510), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n548), .B2(new_n486), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n576), .A2(new_n592), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n550), .B2(new_n404), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n337), .B1(new_n554), .B2(new_n597), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n308), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n544), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n591), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT16), .B(G8gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n605), .B(KEYINPUT42), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(G8gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT96), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT97), .ZN(G1325gat));
  NAND2_X1  g409(.A1(new_n546), .A2(new_n549), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(G15gat), .B1(new_n599), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n593), .A2(new_n595), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n599), .A2(G15gat), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(G1326gat));
  NAND2_X1  g416(.A1(new_n599), .A2(new_n577), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT98), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT43), .B(G22gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(G1327gat));
  INV_X1    g420(.A(new_n254), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n554), .A2(new_n597), .ZN(new_n623));
  INV_X1    g422(.A(new_n284), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(KEYINPUT44), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n307), .B(KEYINPUT100), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n626), .A2(new_n240), .A3(new_n337), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n544), .A2(new_n509), .ZN(new_n628));
  AOI21_X1  g427(.A(KEYINPUT101), .B1(new_n628), .B2(new_n577), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n550), .A2(new_n630), .A3(new_n404), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n570), .A2(new_n505), .B1(new_n572), .B2(new_n573), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n541), .A2(new_n558), .A3(new_n543), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n583), .A2(new_n586), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n539), .A3(new_n587), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n404), .B1(new_n639), .B2(new_n509), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n614), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT102), .B1(new_n632), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n628), .A2(KEYINPUT101), .A3(new_n577), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n630), .B1(new_n550), .B2(new_n404), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n596), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n284), .B1(new_n648), .B2(new_n554), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n625), .B(new_n627), .C1(new_n649), .C2(KEYINPUT44), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n545), .A2(new_n553), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n654), .B1(new_n642), .B2(new_n647), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n653), .B1(new_n655), .B2(new_n284), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n656), .A2(KEYINPUT103), .A3(new_n625), .A4(new_n627), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n622), .B1(new_n659), .B2(new_n544), .ZN(new_n660));
  INV_X1    g459(.A(new_n307), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n239), .A2(new_n624), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n598), .A3(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n666), .A2(new_n544), .A3(new_n622), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n667), .B(KEYINPUT45), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n660), .A2(new_n668), .ZN(G1328gat));
  OAI21_X1  g468(.A(G36gat), .B1(new_n659), .B2(new_n509), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n666), .A2(G36gat), .A3(new_n509), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT46), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(G1329gat));
  OR3_X1    g472(.A1(new_n666), .A2(G43gat), .A3(new_n611), .ZN(new_n674));
  OAI21_X1  g473(.A(G43gat), .B1(new_n650), .B2(new_n614), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT47), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n653), .B(new_n284), .C1(new_n554), .C2(new_n597), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n596), .A2(new_n643), .A3(new_n646), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n643), .B1(new_n596), .B2(new_n646), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n554), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n624), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n681), .B2(new_n653), .ZN(new_n682));
  AOI21_X1  g481(.A(KEYINPUT103), .B1(new_n682), .B2(new_n627), .ZN(new_n683));
  INV_X1    g482(.A(new_n657), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n615), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT105), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(G43gat), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n614), .B1(new_n652), .B2(new_n657), .ZN(new_n688));
  INV_X1    g487(.A(G43gat), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT105), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n687), .A2(new_n690), .A3(new_n674), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n692));
  AND3_X1   g491(.A1(new_n691), .A2(KEYINPUT106), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(KEYINPUT106), .B1(new_n691), .B2(new_n692), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n676), .B1(new_n693), .B2(new_n694), .ZN(G1330gat));
  NOR3_X1   g494(.A1(new_n666), .A2(G50gat), .A3(new_n404), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G50gat), .B1(new_n650), .B2(new_n404), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(KEYINPUT48), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n658), .A2(new_n577), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n696), .B1(new_n700), .B2(G50gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n701), .B2(KEYINPUT48), .ZN(G1331gat));
  XOR2_X1   g501(.A(new_n307), .B(KEYINPUT100), .Z(new_n703));
  NAND2_X1  g502(.A1(new_n334), .A2(new_n336), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n285), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT107), .Z(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n655), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n544), .B(KEYINPUT108), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n591), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT109), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n707), .A2(new_n716), .A3(new_n591), .A4(new_n712), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n714), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(G1333gat));
  NAND3_X1  g519(.A1(new_n707), .A2(G71gat), .A3(new_n615), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n706), .A2(new_n611), .A3(new_n655), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n722), .B2(G71gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n577), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g525(.A1(new_n240), .A2(new_n704), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n649), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(new_n307), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n514), .A3(new_n600), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n656), .A2(new_n307), .A3(new_n625), .A4(new_n727), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n544), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT110), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n732), .B1(new_n735), .B2(new_n514), .ZN(G1336gat));
  INV_X1    g535(.A(G92gat), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n730), .A2(new_n737), .A3(new_n591), .A4(new_n626), .ZN(new_n738));
  OAI21_X1  g537(.A(G92gat), .B1(new_n733), .B2(new_n509), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT111), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n741), .B(G92gat), .C1(new_n733), .C2(new_n509), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n738), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT52), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n733), .A2(KEYINPUT112), .A3(new_n509), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT112), .B1(new_n733), .B2(new_n509), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(G92gat), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n748), .A3(new_n738), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n744), .A2(new_n749), .A3(KEYINPUT113), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1337gat));
  NAND3_X1  g553(.A1(new_n731), .A2(new_n244), .A3(new_n612), .ZN(new_n755));
  OAI21_X1  g554(.A(G99gat), .B1(new_n733), .B2(new_n614), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1338gat));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(KEYINPUT53), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n730), .A2(new_n245), .A3(new_n577), .A4(new_n626), .ZN(new_n760));
  OAI21_X1  g559(.A(G106gat), .B1(new_n733), .B2(new_n404), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n758), .A2(KEYINPUT53), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n762), .B(new_n763), .Z(G1339gat));
  INV_X1    g563(.A(KEYINPUT54), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(new_n294), .B2(new_n295), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n288), .A2(new_n292), .A3(new_n289), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n305), .A2(KEYINPUT54), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n303), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n766), .A2(KEYINPUT55), .A3(new_n768), .A4(new_n303), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n306), .A3(new_n772), .ZN(new_n773));
  OAI22_X1  g572(.A1(new_n316), .A2(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n332), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n336), .B(new_n775), .C1(new_n281), .C2(new_n283), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n307), .A2(new_n336), .A3(new_n775), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n337), .B2(new_n773), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(new_n284), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT115), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n704), .A2(new_n306), .A3(new_n771), .A4(new_n772), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n624), .B1(new_n783), .B2(new_n778), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n784), .B2(new_n777), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n781), .A2(new_n785), .A3(new_n239), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n308), .A2(new_n337), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n708), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n512), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n446), .A3(new_n704), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n239), .B1(new_n780), .B2(KEYINPUT115), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n784), .A2(new_n782), .A3(new_n777), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n544), .A2(new_n591), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n611), .A2(new_n577), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n796), .A2(KEYINPUT116), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(KEYINPUT116), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n799), .A2(new_n704), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n790), .B1(new_n800), .B2(new_n446), .ZN(G1340gat));
  NAND3_X1  g600(.A1(new_n789), .A2(new_n444), .A3(new_n307), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n797), .A2(new_n626), .A3(new_n798), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n803), .A2(KEYINPUT117), .A3(G120gat), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT117), .B1(new_n803), .B2(G120gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1341gat));
  AOI21_X1  g605(.A(G127gat), .B1(new_n789), .B2(new_n240), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n239), .A2(new_n439), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n799), .B2(new_n808), .ZN(G1342gat));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n437), .A3(new_n624), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT56), .Z(new_n811));
  NAND2_X1  g610(.A1(new_n799), .A2(new_n624), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G134gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(G1343gat));
  NAND2_X1  g613(.A1(new_n614), .A2(new_n794), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT118), .ZN(new_n816));
  XOR2_X1   g615(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n817));
  AOI21_X1  g616(.A(new_n817), .B1(new_n793), .B2(new_n577), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n769), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT55), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n769), .A2(new_n820), .A3(new_n770), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n822), .A2(new_n704), .A3(new_n306), .A4(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n624), .B1(new_n824), .B2(new_n778), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n239), .B1(new_n825), .B2(new_n777), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n819), .B(new_n404), .C1(new_n787), .C2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n704), .B(new_n816), .C1(new_n818), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(G141gat), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n788), .A2(KEYINPUT121), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n615), .A2(new_n404), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n788), .B2(KEYINPUT121), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n830), .A2(new_n833), .A3(new_n704), .A4(new_n509), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n829), .B1(new_n834), .B2(G141gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT58), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n829), .B(new_n837), .C1(new_n834), .C2(G141gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1344gat));
  OR2_X1    g638(.A1(new_n818), .A2(new_n827), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n816), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n307), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n787), .A2(new_n826), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n819), .B1(new_n844), .B2(new_n404), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n793), .A2(new_n577), .A3(new_n817), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n307), .A3(new_n816), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n830), .A2(new_n833), .A3(new_n509), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n842), .B1(new_n850), .B2(new_n307), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n843), .B(new_n849), .C1(new_n851), .C2(G148gat), .ZN(G1345gat));
  AOI21_X1  g651(.A(G155gat), .B1(new_n850), .B2(new_n240), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n239), .A2(new_n349), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n853), .B1(new_n841), .B2(new_n854), .ZN(G1346gat));
  OAI211_X1 g654(.A(new_n624), .B(new_n816), .C1(new_n818), .C2(new_n827), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT122), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(KEYINPUT122), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(G162gat), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n850), .A2(new_n350), .A3(new_n624), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1347gat));
  AND2_X1   g660(.A1(new_n793), .A2(new_n795), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n709), .A2(new_n509), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G169gat), .B1(new_n864), .B2(new_n337), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n600), .B1(new_n786), .B2(new_n787), .ZN(new_n866));
  NOR4_X1   g665(.A1(new_n577), .A2(new_n548), .A3(new_n509), .A4(new_n486), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT123), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n869), .A2(G169gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n865), .B1(new_n337), .B2(new_n870), .ZN(G1348gat));
  AND2_X1   g670(.A1(new_n862), .A2(new_n863), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(G176gat), .A3(new_n626), .ZN(new_n873));
  INV_X1    g672(.A(new_n869), .ZN(new_n874));
  AOI21_X1  g673(.A(G176gat), .B1(new_n874), .B2(new_n307), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n873), .A2(new_n875), .ZN(G1349gat));
  OAI21_X1  g675(.A(G183gat), .B1(new_n864), .B2(new_n239), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n418), .A2(KEYINPUT27), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n422), .A2(G183gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n874), .A2(new_n878), .A3(new_n879), .A4(new_n240), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n874), .A2(new_n460), .A3(new_n624), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n460), .B1(new_n872), .B2(new_n624), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(G1351gat));
  NAND3_X1  g687(.A1(new_n866), .A2(new_n591), .A3(new_n831), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n889), .A2(G197gat), .A3(new_n337), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n709), .A2(new_n509), .A3(new_n615), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT124), .Z(new_n892));
  AOI211_X1 g691(.A(new_n337), .B(new_n892), .C1(new_n845), .C2(new_n846), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n890), .B1(new_n893), .B2(new_n329), .ZN(G1352gat));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n896));
  INV_X1    g695(.A(G204gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n307), .A2(new_n897), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n889), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n895), .A2(KEYINPUT125), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n889), .A2(new_n898), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n703), .B(new_n892), .C1(new_n845), .C2(new_n846), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n899), .B(new_n901), .C1(new_n897), .C2(new_n902), .ZN(G1353gat));
  OR3_X1    g702(.A1(new_n889), .A2(G211gat), .A3(new_n239), .ZN(new_n904));
  INV_X1    g703(.A(new_n892), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n847), .A2(new_n240), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT63), .B1(new_n906), .B2(G211gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(G1354gat));
  OR2_X1    g708(.A1(new_n889), .A2(new_n284), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT126), .ZN(new_n911));
  INV_X1    g710(.A(G218gat), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n911), .B1(new_n910), .B2(new_n912), .ZN(new_n914));
  AND4_X1   g713(.A1(G218gat), .A2(new_n847), .A3(new_n624), .A4(new_n905), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(G1355gat));
endmodule


