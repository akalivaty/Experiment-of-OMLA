

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578;

  NAND2_X1 U322 ( .A1(n548), .A2(n557), .ZN(n365) );
  INV_X1 U323 ( .A(n559), .ZN(n573) );
  INV_X1 U324 ( .A(n569), .ZN(n404) );
  XOR2_X1 U325 ( .A(G8GAT), .B(G183GAT), .Z(n412) );
  NAND2_X1 U326 ( .A1(n519), .A2(n516), .ZN(n456) );
  NOR2_X1 U327 ( .A1(n573), .A2(n576), .ZN(n403) );
  NOR2_X1 U328 ( .A1(n522), .A2(n541), .ZN(n527) );
  NOR2_X1 U329 ( .A1(n513), .A2(n487), .ZN(n489) );
  XNOR2_X1 U330 ( .A(n552), .B(n402), .ZN(n576) );
  AND2_X1 U331 ( .A1(n448), .A2(n519), .ZN(n449) );
  XNOR2_X1 U332 ( .A(KEYINPUT122), .B(n449), .ZN(n556) );
  XOR2_X2 U333 ( .A(n381), .B(n380), .Z(n552) );
  XOR2_X2 U334 ( .A(n447), .B(n446), .Z(n519) );
  NOR2_X1 U335 ( .A1(n514), .A2(n427), .ZN(n562) );
  AND2_X1 U336 ( .A1(n464), .A2(n562), .ZN(n428) );
  XOR2_X1 U337 ( .A(KEYINPUT41), .B(n404), .Z(n548) );
  XOR2_X1 U338 ( .A(KEYINPUT45), .B(n403), .Z(n290) );
  XOR2_X1 U339 ( .A(n378), .B(n377), .Z(n291) );
  XOR2_X1 U340 ( .A(G57GAT), .B(KEYINPUT13), .Z(n384) );
  XNOR2_X1 U341 ( .A(n338), .B(KEYINPUT69), .ZN(n339) );
  XNOR2_X1 U342 ( .A(n340), .B(n339), .ZN(n343) );
  XNOR2_X1 U343 ( .A(n345), .B(n420), .ZN(n346) );
  XNOR2_X1 U344 ( .A(n347), .B(n346), .ZN(n569) );
  XNOR2_X1 U345 ( .A(n453), .B(G190GAT), .ZN(n454) );
  XNOR2_X1 U346 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  INV_X1 U347 ( .A(KEYINPUT55), .ZN(n429) );
  XNOR2_X1 U348 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n292) );
  XNOR2_X1 U349 ( .A(n292), .B(KEYINPUT82), .ZN(n293) );
  XOR2_X1 U350 ( .A(n293), .B(KEYINPUT83), .Z(n295) );
  XNOR2_X1 U351 ( .A(G197GAT), .B(G218GAT), .ZN(n294) );
  XOR2_X1 U352 ( .A(n295), .B(n294), .Z(n423) );
  XOR2_X1 U353 ( .A(G155GAT), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U354 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n317) );
  XOR2_X1 U356 ( .A(n317), .B(KEYINPUT23), .Z(n299) );
  XOR2_X1 U357 ( .A(G141GAT), .B(G22GAT), .Z(n352) );
  XNOR2_X1 U358 ( .A(n352), .B(KEYINPUT85), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U360 ( .A(n423), .B(n300), .Z(n310) );
  XOR2_X1 U361 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n302) );
  NAND2_X1 U362 ( .A1(G228GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U364 ( .A(n303), .B(KEYINPUT24), .Z(n308) );
  XNOR2_X1 U365 ( .A(G50GAT), .B(KEYINPUT70), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n304), .B(G162GAT), .ZN(n371) );
  XOR2_X1 U367 ( .A(G78GAT), .B(G148GAT), .Z(n306) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(G204GAT), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n345) );
  XNOR2_X1 U370 ( .A(n371), .B(n345), .ZN(n307) );
  XNOR2_X1 U371 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U372 ( .A(n310), .B(n309), .ZN(n464) );
  XOR2_X1 U373 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n312) );
  XNOR2_X1 U374 ( .A(KEYINPUT89), .B(KEYINPUT88), .ZN(n311) );
  XNOR2_X1 U375 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U376 ( .A(G1GAT), .B(n313), .Z(n315) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U378 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U379 ( .A(n316), .B(KEYINPUT87), .Z(n322) );
  XOR2_X1 U380 ( .A(G134GAT), .B(KEYINPUT71), .Z(n374) );
  XOR2_X1 U381 ( .A(G85GAT), .B(n374), .Z(n319) );
  XNOR2_X1 U382 ( .A(G162GAT), .B(n317), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U384 ( .A(n320), .B(KEYINPUT91), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U386 ( .A(G148GAT), .B(G120GAT), .Z(n324) );
  XNOR2_X1 U387 ( .A(G29GAT), .B(G141GAT), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U389 ( .A(n326), .B(n325), .Z(n334) );
  XOR2_X1 U390 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n328) );
  XNOR2_X1 U391 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U393 ( .A(G113GAT), .B(n329), .Z(n447) );
  XOR2_X1 U394 ( .A(KEYINPUT4), .B(G57GAT), .Z(n331) );
  XNOR2_X1 U395 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n447), .B(n332), .ZN(n333) );
  XOR2_X1 U398 ( .A(n334), .B(n333), .Z(n462) );
  INV_X1 U399 ( .A(n462), .ZN(n514) );
  XNOR2_X1 U400 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n335) );
  XNOR2_X1 U401 ( .A(n335), .B(KEYINPUT54), .ZN(n426) );
  XOR2_X1 U402 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U403 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n336), .B(n384), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n439), .B(n337), .ZN(n340) );
  AND2_X1 U406 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(G99GAT), .B(G85GAT), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n341), .B(KEYINPUT68), .ZN(n370) );
  XOR2_X1 U409 ( .A(n370), .B(KEYINPUT31), .Z(n342) );
  XNOR2_X1 U410 ( .A(n343), .B(n342), .ZN(n347) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(G92GAT), .ZN(n344) );
  XOR2_X1 U412 ( .A(n344), .B(G64GAT), .Z(n420) );
  XOR2_X1 U413 ( .A(G8GAT), .B(G197GAT), .Z(n349) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(G113GAT), .ZN(n348) );
  XNOR2_X1 U415 ( .A(n349), .B(n348), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n351) );
  XNOR2_X1 U417 ( .A(KEYINPUT65), .B(KEYINPUT66), .ZN(n350) );
  XNOR2_X1 U418 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U419 ( .A(G36GAT), .B(G50GAT), .Z(n354) );
  XOR2_X1 U420 ( .A(G15GAT), .B(G1GAT), .Z(n394) );
  XNOR2_X1 U421 ( .A(n352), .B(n394), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U423 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U424 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U427 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n362) );
  XNOR2_X1 U428 ( .A(G43GAT), .B(G29GAT), .ZN(n361) );
  XNOR2_X1 U429 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U430 ( .A(KEYINPUT67), .B(n363), .Z(n366) );
  XOR2_X1 U431 ( .A(n364), .B(n366), .Z(n557) );
  XNOR2_X1 U432 ( .A(n365), .B(KEYINPUT46), .ZN(n400) );
  INV_X1 U433 ( .A(n366), .ZN(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n368) );
  NAND2_X1 U435 ( .A1(G232GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U436 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U437 ( .A(n369), .B(KEYINPUT9), .Z(n373) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U440 ( .A(G36GAT), .B(G190GAT), .Z(n413) );
  XOR2_X1 U441 ( .A(n413), .B(G92GAT), .Z(n376) );
  XNOR2_X1 U442 ( .A(G106GAT), .B(n374), .ZN(n375) );
  XNOR2_X1 U443 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U444 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n291), .B(n379), .ZN(n380) );
  XOR2_X1 U446 ( .A(G78GAT), .B(G211GAT), .Z(n383) );
  XNOR2_X1 U447 ( .A(G127GAT), .B(G71GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n398) );
  XOR2_X1 U449 ( .A(n384), .B(n412), .Z(n386) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U452 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n388) );
  XNOR2_X1 U453 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n387) );
  XNOR2_X1 U454 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U455 ( .A(n390), .B(n389), .Z(n396) );
  XOR2_X1 U456 ( .A(KEYINPUT12), .B(G64GAT), .Z(n392) );
  XNOR2_X1 U457 ( .A(G22GAT), .B(G155GAT), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n559) );
  NOR2_X1 U462 ( .A1(n552), .A2(n559), .ZN(n399) );
  AND2_X1 U463 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n401), .B(KEYINPUT47), .ZN(n407) );
  XNOR2_X1 U465 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n402) );
  NOR2_X1 U466 ( .A1(n404), .A2(n290), .ZN(n405) );
  INV_X1 U467 ( .A(n557), .ZN(n563) );
  NAND2_X1 U468 ( .A1(n405), .A2(n563), .ZN(n406) );
  NAND2_X1 U469 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n408), .B(KEYINPUT48), .ZN(n540) );
  XOR2_X1 U471 ( .A(KEYINPUT19), .B(KEYINPUT79), .Z(n410) );
  XNOR2_X1 U472 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n409) );
  XNOR2_X1 U473 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U474 ( .A(G169GAT), .B(n411), .Z(n443) );
  XOR2_X1 U475 ( .A(KEYINPUT94), .B(n412), .Z(n415) );
  XNOR2_X1 U476 ( .A(G204GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U478 ( .A(n443), .B(n416), .Z(n418) );
  NAND2_X1 U479 ( .A1(G226GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U481 ( .A(n419), .B(KEYINPUT92), .Z(n422) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(n420), .Z(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n516) );
  NAND2_X1 U485 ( .A1(n540), .A2(n516), .ZN(n425) );
  XOR2_X1 U486 ( .A(n426), .B(n425), .Z(n427) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n448) );
  XOR2_X1 U488 ( .A(G176GAT), .B(G183GAT), .Z(n431) );
  XNOR2_X1 U489 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U491 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n433) );
  XNOR2_X1 U492 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n445) );
  XOR2_X1 U495 ( .A(G99GAT), .B(G134GAT), .Z(n437) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G190GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U499 ( .A1(G227GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U500 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U503 ( .A1(n556), .A2(n548), .ZN(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n450) );
  XNOR2_X1 U505 ( .A(n450), .B(G176GAT), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  NAND2_X1 U507 ( .A1(n556), .A2(n552), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n453) );
  XOR2_X1 U509 ( .A(KEYINPUT95), .B(n456), .Z(n457) );
  NAND2_X1 U510 ( .A1(n464), .A2(n457), .ZN(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT25), .B(n458), .Z(n461) );
  NOR2_X1 U512 ( .A1(n464), .A2(n519), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT26), .ZN(n561) );
  XNOR2_X1 U514 ( .A(n516), .B(KEYINPUT27), .ZN(n465) );
  NAND2_X1 U515 ( .A1(n561), .A2(n465), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n461), .A2(n460), .ZN(n463) );
  NAND2_X1 U517 ( .A1(n463), .A2(n462), .ZN(n467) );
  XOR2_X1 U518 ( .A(n464), .B(KEYINPUT28), .Z(n522) );
  NAND2_X1 U519 ( .A1(n514), .A2(n465), .ZN(n541) );
  INV_X1 U520 ( .A(n519), .ZN(n529) );
  NAND2_X1 U521 ( .A1(n527), .A2(n529), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n483) );
  XOR2_X1 U523 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n469) );
  OR2_X1 U524 ( .A1(n552), .A2(n573), .ZN(n468) );
  XNOR2_X1 U525 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U526 ( .A1(n483), .A2(n470), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n471), .B(KEYINPUT96), .ZN(n500) );
  NAND2_X1 U528 ( .A1(n557), .A2(n569), .ZN(n487) );
  NOR2_X1 U529 ( .A1(n500), .A2(n487), .ZN(n480) );
  NAND2_X1 U530 ( .A1(n480), .A2(n514), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT34), .ZN(n473) );
  XOR2_X1 U532 ( .A(n473), .B(KEYINPUT98), .Z(n475) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n480), .A2(n516), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n478) );
  NAND2_X1 U538 ( .A1(n480), .A2(n519), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U540 ( .A(G15GAT), .B(n479), .Z(G1326GAT) );
  NAND2_X1 U541 ( .A1(n480), .A2(n522), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(KEYINPUT100), .ZN(n482) );
  XNOR2_X1 U543 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  XNOR2_X1 U544 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n493) );
  NAND2_X1 U545 ( .A1(n573), .A2(n483), .ZN(n484) );
  NOR2_X1 U546 ( .A1(n576), .A2(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n513) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U551 ( .A(KEYINPUT104), .B(n490), .Z(n497) );
  NAND2_X1 U552 ( .A1(n497), .A2(n514), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n497), .A2(n516), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n497), .A2(n519), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(KEYINPUT40), .ZN(n496) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n497), .A2(n522), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(KEYINPUT106), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n502) );
  NAND2_X1 U564 ( .A1(n563), .A2(n548), .ZN(n512) );
  NOR2_X1 U565 ( .A1(n500), .A2(n512), .ZN(n507) );
  NAND2_X1 U566 ( .A1(n507), .A2(n514), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n507), .A2(n516), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(KEYINPUT108), .ZN(n505) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n507), .A2(n519), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n506), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U575 ( .A1(n507), .A2(n522), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT110), .Z(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n514), .A2(n523), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  XOR2_X1 U582 ( .A(G92GAT), .B(KEYINPUT111), .Z(n518) );
  NAND2_X1 U583 ( .A1(n523), .A2(n516), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n519), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(KEYINPUT112), .ZN(n521) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n525) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NAND2_X1 U592 ( .A1(n540), .A2(n527), .ZN(n528) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n557), .A2(n536), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U597 ( .A1(n536), .A2(n548), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U600 ( .A1(n559), .A2(n536), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U604 ( .A1(n536), .A2(n552), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U606 ( .A(G134GAT), .B(n539), .Z(G1343GAT) );
  NAND2_X1 U607 ( .A1(n540), .A2(n561), .ZN(n542) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n543), .B(KEYINPUT116), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n553), .A2(n557), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n544), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U615 ( .A(KEYINPUT117), .B(n547), .Z(n550) );
  NAND2_X1 U616 ( .A1(n548), .A2(n553), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n559), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U620 ( .A(G162GAT), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n556), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n575) );
  NOR2_X1 U628 ( .A1(n563), .A2(n575), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n565) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT124), .B(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n575), .ZN(n571) );
  XNOR2_X1 U635 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

