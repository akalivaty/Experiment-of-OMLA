//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(KEYINPUT65), .A3(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT2), .B(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  XOR2_X1   g010(.A(KEYINPUT2), .B(G113), .Z(new_n197));
  OAI211_X1 g011(.A(new_n197), .B(new_n189), .C1(new_n193), .C2(new_n192), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G137), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n201), .A2(G137), .ZN(new_n204));
  OAI21_X1  g018(.A(G131), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n201), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n207), .A2(new_n209), .A3(new_n210), .A4(new_n202), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n205), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  INV_X1    g029(.A(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n215), .A2(new_n217), .A3(new_n219), .A4(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI22_X1  g038(.A1(new_n215), .A2(new_n217), .B1(new_n219), .B2(G128), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT67), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n228));
  AOI211_X1 g042(.A(new_n228), .B(new_n225), .C1(new_n221), .C2(new_n223), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n200), .B(new_n213), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n207), .A2(new_n209), .A3(new_n202), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n211), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  OR2_X1    g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n218), .A2(G143), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n216), .A2(G146), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n236), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT0), .A4(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n232), .A2(KEYINPUT66), .A3(new_n211), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n235), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n230), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G143), .B(G146), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n222), .B1(new_n247), .B2(new_n215), .ZN(new_n248));
  AND4_X1   g062(.A1(new_n222), .A2(new_n215), .A3(new_n217), .A4(new_n219), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n226), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n228), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n225), .B1(new_n221), .B2(new_n223), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n200), .B1(new_n254), .B2(new_n213), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT30), .B1(new_n246), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n243), .A2(new_n233), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n212), .B2(new_n252), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT30), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n199), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n213), .B1(new_n227), .B2(new_n229), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT68), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n199), .B(KEYINPUT69), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n230), .A4(new_n245), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT26), .B(G101), .ZN(new_n266));
  INV_X1    g080(.A(G237), .ZN(new_n267));
  INV_X1    g081(.A(G953), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(G210), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n266), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n265), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT31), .B1(new_n261), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n272), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n246), .A2(new_n255), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n275), .B1(new_n276), .B2(new_n264), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n263), .A2(new_n230), .A3(new_n245), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n259), .B1(new_n279), .B2(KEYINPUT30), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n277), .B(new_n278), .C1(new_n280), .C2(new_n199), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n196), .A2(new_n198), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n258), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n265), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(KEYINPUT69), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n286), .B1(new_n213), .B2(new_n254), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT28), .B1(new_n287), .B2(new_n245), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n275), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n274), .A2(new_n281), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  XOR2_X1   g106(.A(new_n292), .B(KEYINPUT71), .Z(new_n293));
  AND3_X1   g107(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n290), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n187), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n290), .A2(KEYINPUT32), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n290), .A2(new_n299), .A3(KEYINPUT32), .A4(new_n293), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n265), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n275), .B1(new_n261), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n285), .A2(new_n288), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n275), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n279), .A2(new_n286), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n265), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n288), .B1(new_n308), .B2(KEYINPUT28), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n275), .A2(new_n304), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G472), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n301), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n315));
  INV_X1    g129(.A(G221), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT9), .B(G234), .Z(new_n317));
  INV_X1    g131(.A(G902), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n268), .A2(G227), .ZN(new_n322));
  XOR2_X1   g136(.A(new_n321), .B(new_n322), .Z(new_n323));
  NAND2_X1  g137(.A1(new_n235), .A2(new_n244), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  INV_X1    g140(.A(G104), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G107), .ZN(new_n328));
  INV_X1    g142(.A(G107), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT3), .A3(G104), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n328), .A2(new_n330), .B1(new_n327), .B2(G107), .ZN(new_n331));
  INV_X1    g145(.A(G101), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT78), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G101), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n327), .A2(G107), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n329), .A2(G104), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n331), .A2(new_n336), .B1(G101), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT10), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n251), .B2(new_n253), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n328), .A2(new_n330), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n337), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n343), .A2(new_n336), .A3(new_n337), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n331), .A2(new_n332), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n243), .B(new_n346), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n339), .A2(G101), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n351), .B1(new_n252), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n325), .B1(new_n342), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(KEYINPUT79), .B(new_n325), .C1(new_n342), .C2(new_n355), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(KEYINPUT10), .B(new_n340), .C1(new_n227), .C2(new_n229), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n361), .A2(new_n324), .A3(new_n350), .A4(new_n354), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n323), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n252), .B(new_n353), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n364), .A2(KEYINPUT12), .A3(new_n233), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT12), .B1(new_n364), .B2(new_n325), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n323), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n320), .B(new_n318), .C1(new_n363), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n368), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n372));
  INV_X1    g186(.A(new_n323), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n360), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(G469), .B1(new_n374), .B2(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n319), .B1(new_n370), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n380), .B(new_n226), .C1(new_n248), .C2(new_n249), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n242), .A2(G125), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT81), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n240), .B2(new_n241), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT82), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT82), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n382), .A2(KEYINPUT81), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n384), .B1(new_n252), .B2(new_n380), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(KEYINPUT81), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G224), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(new_n391), .A3(new_n394), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n283), .B(new_n346), .C1(new_n349), .C2(new_n348), .ZN(new_n399));
  XNOR2_X1  g213(.A(G110), .B(G122), .ZN(new_n400));
  OAI211_X1 g214(.A(KEYINPUT5), .B(new_n189), .C1(new_n192), .C2(new_n193), .ZN(new_n401));
  INV_X1    g215(.A(G113), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n193), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n340), .A2(new_n405), .A3(new_n198), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n399), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n400), .A2(KEYINPUT80), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n399), .B2(new_n406), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n407), .B1(new_n410), .B2(KEYINPUT6), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n412), .B(new_n409), .C1(new_n399), .C2(new_n406), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n379), .B1(new_n398), .B2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n387), .A2(new_n394), .A3(new_n391), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n394), .B1(new_n387), .B2(new_n391), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n399), .A2(new_n406), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n412), .B1(new_n419), .B2(new_n409), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n410), .A2(KEYINPUT6), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(new_n407), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n418), .A2(new_n422), .A3(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n395), .A2(KEYINPUT7), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(new_n389), .C1(new_n390), .C2(KEYINPUT81), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT84), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n405), .A2(new_n198), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n353), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n406), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n400), .B(KEYINPUT8), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n381), .A2(new_n382), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n432), .A2(new_n433), .B1(new_n425), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n385), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT84), .A3(new_n426), .A4(new_n389), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n429), .A2(new_n435), .A3(new_n437), .A4(new_n407), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n318), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(KEYINPUT85), .A3(new_n318), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n378), .B1(new_n424), .B2(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n424), .A2(new_n443), .A3(new_n378), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n376), .B(new_n377), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT89), .B(G104), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G125), .B(G140), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(G146), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT86), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n267), .A2(new_n268), .A3(G214), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n216), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT18), .A2(G131), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n461), .B1(new_n456), .B2(G131), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n455), .B(G143), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(KEYINPUT87), .A3(new_n210), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n456), .A2(G131), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n452), .A2(KEYINPUT16), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n380), .A2(KEYINPUT16), .A3(G140), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(G146), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT19), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(KEYINPUT88), .ZN(new_n472));
  MUX2_X1   g286(.A(new_n470), .B(new_n472), .S(new_n452), .Z(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n218), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n466), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n451), .B1(new_n460), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n467), .A2(new_n468), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n218), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n469), .ZN(new_n479));
  INV_X1    g293(.A(new_n465), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(KEYINPUT17), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(KEYINPUT17), .B2(new_n466), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n450), .A3(new_n459), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n447), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n447), .A3(new_n485), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n483), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n450), .B1(new_n482), .B2(new_n459), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n318), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G475), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n268), .A2(G952), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(G234), .B2(G237), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT21), .B(G898), .Z(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n318), .B(new_n268), .C1(G234), .C2(G237), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n191), .A2(G122), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n329), .B1(new_n502), .B2(KEYINPUT14), .ZN(new_n503));
  XNOR2_X1  g317(.A(G116), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G128), .B(G143), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT90), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n201), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n507), .A2(new_n201), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n504), .B(new_n329), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n214), .A2(G143), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n214), .A2(G143), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(KEYINPUT13), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(KEYINPUT13), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n508), .B(new_n512), .C1(new_n516), .C2(new_n201), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n317), .A2(G217), .A3(new_n268), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n519), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(G902), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G478), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n523), .A2(KEYINPUT91), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n525), .ZN(new_n527));
  INV_X1    g341(.A(new_n523), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT91), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n523), .A2(KEYINPUT91), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n526), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n494), .A2(new_n501), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n315), .B1(new_n446), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G234), .ZN(new_n536));
  OAI21_X1  g350(.A(G217), .B1(new_n536), .B2(G902), .ZN(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  OR3_X1    g352(.A1(new_n188), .A2(KEYINPUT23), .A3(G128), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT23), .B1(new_n188), .B2(G128), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n214), .A2(G119), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT74), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n214), .B2(G119), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n188), .A2(KEYINPUT74), .A3(G128), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n544), .A2(new_n545), .B1(G119), .B2(new_n214), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT24), .B(G110), .Z(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  OAI221_X1 g363(.A(new_n479), .B1(new_n538), .B2(new_n542), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(KEYINPUT75), .A3(new_n549), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n542), .A2(new_n538), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT75), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n546), .B2(new_n548), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n452), .A2(new_n218), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n469), .A3(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT76), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n550), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT22), .B(G137), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n316), .A2(new_n536), .A3(G953), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n550), .B(new_n564), .C1(new_n559), .C2(new_n560), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n318), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n537), .B1(new_n568), .B2(KEYINPUT25), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(KEYINPUT25), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n536), .B2(G217), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT77), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(KEYINPUT77), .A3(new_n573), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n489), .A2(new_n493), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n580), .A2(new_n532), .A3(new_n500), .ZN(new_n581));
  INV_X1    g395(.A(new_n377), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n398), .A2(new_n414), .A3(new_n379), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT83), .B1(new_n418), .B2(new_n422), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT85), .B1(new_n438), .B2(new_n318), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n438), .A2(KEYINPUT85), .A3(new_n318), .ZN(new_n586));
  OAI22_X1  g400(.A1(new_n583), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n378), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n424), .A2(new_n443), .A3(new_n378), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n582), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n581), .A2(new_n591), .A3(KEYINPUT92), .A4(new_n376), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n314), .A2(new_n535), .A3(new_n579), .A4(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(new_n336), .Z(G3));
  NOR2_X1   g408(.A1(new_n294), .A2(new_n295), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n290), .A2(new_n318), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n377), .B(new_n501), .C1(new_n445), .C2(new_n444), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(KEYINPUT93), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n520), .B2(new_n522), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n601), .A2(KEYINPUT93), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n603), .A2(new_n605), .ZN(new_n607));
  OAI211_X1 g421(.A(G478), .B(new_n318), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n528), .A2(new_n524), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n580), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n600), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n376), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n578), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n599), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT34), .B(G104), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(KEYINPUT95), .ZN(new_n618));
  INV_X1    g432(.A(new_n488), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n619), .A2(new_n620), .B1(new_n492), .B2(G475), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n487), .A2(KEYINPUT94), .A3(new_n488), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n532), .A3(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n618), .B1(new_n600), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n623), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n591), .A2(new_n625), .A3(KEYINPUT95), .A4(new_n501), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n599), .A3(new_n614), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(new_n329), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G9));
  NOR2_X1   g445(.A1(new_n565), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n561), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n573), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n570), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n535), .A2(new_n592), .A3(new_n599), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT37), .B(G110), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n636), .B(new_n638), .ZN(G12));
  INV_X1    g453(.A(G900), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n496), .B1(new_n499), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n621), .A2(new_n532), .A3(new_n622), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n446), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n314), .A2(new_n635), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(KEYINPUT98), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n314), .A2(new_n644), .A3(new_n647), .A4(new_n635), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  NOR2_X1   g464(.A1(new_n261), .A2(new_n273), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n275), .B2(new_n308), .ZN(new_n652));
  OAI21_X1  g466(.A(G472), .B1(new_n652), .B2(G902), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n296), .A2(new_n301), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT99), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n494), .A2(new_n533), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n377), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n635), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT100), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n641), .B(KEYINPUT39), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n613), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT40), .Z(new_n663));
  NOR2_X1   g477(.A1(new_n445), .A2(new_n444), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT38), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n656), .A2(new_n660), .A3(new_n663), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n216), .ZN(G45));
  NAND3_X1  g481(.A1(new_n580), .A2(new_n610), .A3(new_n642), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n446), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n314), .A2(new_n635), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G146), .ZN(G48));
  NOR2_X1   g485(.A1(new_n363), .A2(new_n369), .ZN(new_n672));
  OAI21_X1  g486(.A(G469), .B1(new_n672), .B2(G902), .ZN(new_n673));
  INV_X1    g487(.A(new_n319), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n370), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n314), .A2(new_n676), .A3(new_n612), .A4(new_n579), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G15));
  NAND4_X1  g493(.A1(new_n627), .A2(new_n314), .A3(new_n579), .A4(new_n676), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  OAI21_X1  g495(.A(new_n377), .B1(new_n445), .B2(new_n444), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n675), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n314), .A2(new_n581), .A3(new_n635), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  OAI211_X1 g499(.A(new_n274), .B(new_n281), .C1(new_n309), .C2(new_n272), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n293), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n597), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n578), .ZN(new_n689));
  INV_X1    g503(.A(new_n600), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n657), .A4(new_n676), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  AND3_X1   g506(.A1(new_n635), .A2(new_n597), .A3(new_n687), .ZN(new_n693));
  INV_X1    g507(.A(new_n668), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n683), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT101), .B(G125), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G27));
  NAND2_X1  g511(.A1(new_n290), .A2(new_n293), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n187), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n297), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n313), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n579), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n589), .A2(new_n377), .A3(new_n590), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT102), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n589), .A2(new_n708), .A3(new_n377), .A4(new_n590), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n707), .A2(new_n376), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n694), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT42), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n668), .A2(KEYINPUT42), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n710), .A2(new_n314), .A3(new_n579), .A4(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n210), .ZN(G33));
  XNOR2_X1  g530(.A(new_n643), .B(KEYINPUT104), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n710), .A2(new_n314), .A3(new_n579), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G134), .ZN(G36));
  INV_X1    g533(.A(new_n610), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n580), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT43), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n722), .A2(new_n635), .ZN(new_n723));
  INV_X1    g537(.A(new_n599), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n725), .A2(KEYINPUT44), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n707), .A2(new_n709), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n725), .A2(KEYINPUT44), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  OR2_X1    g543(.A1(new_n374), .A2(KEYINPUT45), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n374), .A2(KEYINPUT45), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(G469), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(G469), .A2(G902), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n735), .A2(KEYINPUT46), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n370), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n735), .B2(KEYINPUT46), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n736), .A2(new_n737), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n674), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g557(.A1(new_n743), .A2(new_n661), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n729), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n208), .ZN(G39));
  INV_X1    g560(.A(new_n727), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n579), .A3(new_n668), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n314), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G140), .ZN(G42));
  INV_X1    g571(.A(new_n673), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n739), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(KEYINPUT49), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(KEYINPUT49), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n579), .A2(new_n721), .A3(new_n377), .A4(new_n674), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n656), .A2(new_n665), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n680), .A2(new_n677), .A3(new_n684), .A4(new_n691), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n611), .B1(new_n580), .B2(new_n533), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n599), .A2(new_n690), .A3(new_n614), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n593), .A2(new_n636), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n593), .A2(new_n636), .A3(new_n772), .A4(new_n769), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n767), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n710), .A2(new_n694), .A3(new_n693), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n532), .A2(new_n641), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n622), .A2(new_n635), .A3(new_n621), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n710), .A2(new_n314), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n718), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n718), .A2(new_n775), .A3(new_n778), .A4(KEYINPUT108), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n715), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n774), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT109), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n715), .B1(new_n781), .B2(new_n782), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n774), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n766), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n785), .A2(KEYINPUT109), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n787), .A3(new_n774), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(KEYINPUT110), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n670), .A2(new_n695), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n664), .A2(new_n641), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n659), .A2(new_n376), .A3(new_n654), .A4(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n649), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n794), .B1(new_n648), .B2(new_n646), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(KEYINPUT112), .A3(new_n797), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n798), .B2(new_n804), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n801), .A2(KEYINPUT111), .A3(KEYINPUT52), .A4(new_n797), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT53), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n790), .A2(new_n793), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(new_n800), .B2(new_n802), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n800), .A2(KEYINPUT52), .A3(new_n802), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n791), .B(new_n792), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(KEYINPUT54), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n791), .A2(new_n792), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n813), .A2(new_n812), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n805), .A2(new_n809), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n767), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n767), .A2(new_n823), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n817), .B1(new_n771), .B2(new_n773), .ZN(new_n826));
  AND4_X1   g640(.A1(new_n788), .A2(new_n824), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n820), .A2(new_n821), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n816), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n727), .A2(new_n676), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n579), .A2(new_n656), .A3(new_n496), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n494), .A3(new_n720), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n722), .A2(new_n496), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n722), .A2(KEYINPUT115), .A3(new_n496), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n689), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n665), .A2(new_n582), .A3(new_n676), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT116), .Z(new_n842));
  OAI21_X1  g656(.A(KEYINPUT50), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(new_n693), .A3(new_n832), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n834), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n753), .A2(new_n754), .B1(new_n319), .B2(new_n759), .ZN(new_n846));
  OAI22_X1  g660(.A1(new_n846), .A2(new_n747), .B1(KEYINPUT50), .B2(new_n842), .ZN(new_n847));
  INV_X1    g661(.A(new_n840), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n849), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n495), .B1(new_n848), .B2(new_n683), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n705), .B(new_n831), .C1(new_n837), .C2(new_n838), .ZN(new_n855));
  XOR2_X1   g669(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n856));
  OR2_X1    g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n833), .A2(new_n580), .A3(new_n610), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n854), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT118), .Z(new_n861));
  NOR4_X1   g675(.A1(new_n830), .A2(new_n852), .A3(new_n853), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(G952), .A2(G953), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n765), .B1(new_n862), .B2(new_n863), .ZN(G75));
  XNOR2_X1  g678(.A(new_n418), .B(new_n414), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT55), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n820), .A2(new_n828), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(G902), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(G210), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n866), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(G210), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n871), .B(new_n866), .C1(new_n868), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n268), .A2(G952), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n872), .A2(new_n877), .ZN(G51));
  XNOR2_X1  g692(.A(new_n732), .B(KEYINPUT120), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n868), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n733), .B(KEYINPUT57), .Z(new_n881));
  AOI221_X4 g695(.A(KEYINPUT54), .B1(new_n822), .B2(new_n827), .C1(new_n814), .C2(new_n817), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n821), .B1(new_n820), .B2(new_n828), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n672), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT119), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n880), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(KEYINPUT119), .A3(new_n885), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n875), .B1(new_n888), .B2(new_n889), .ZN(G54));
  NAND4_X1  g704(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .A4(new_n484), .ZN(new_n891));
  NAND2_X1  g705(.A1(KEYINPUT58), .A2(G475), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n483), .B(new_n476), .C1(new_n868), .C2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n891), .A2(new_n876), .A3(new_n893), .ZN(G60));
  XNOR2_X1  g708(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n524), .A2(new_n318), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n830), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n606), .A2(new_n607), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n900), .B(new_n898), .C1(new_n882), .C2(new_n883), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n902), .A2(KEYINPUT122), .A3(new_n876), .A4(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n876), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n900), .B1(new_n830), .B2(new_n898), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n908), .ZN(G63));
  XOR2_X1   g723(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n910));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n910), .B(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n867), .A2(new_n633), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n876), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n572), .B1(new_n867), .B2(new_n912), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT61), .ZN(G66));
  OAI21_X1  g731(.A(G953), .B1(new_n498), .B2(new_n393), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n774), .B2(G953), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n414), .B1(G898), .B2(new_n268), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT124), .Z(new_n921));
  XNOR2_X1  g735(.A(new_n919), .B(new_n921), .ZN(G69));
  INV_X1    g736(.A(new_n745), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n662), .A2(new_n768), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n924), .A2(new_n727), .A3(new_n314), .A4(new_n579), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n923), .A2(new_n756), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n801), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n666), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n268), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n280), .B(new_n473), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n934), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n745), .B1(new_n755), .B2(new_n752), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n705), .A2(new_n664), .A3(new_n658), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n784), .B(new_n718), .C1(new_n744), .C2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n939), .A2(new_n927), .ZN(new_n940));
  AOI21_X1  g754(.A(G953), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n268), .A2(G900), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT125), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n936), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n935), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n268), .B1(G227), .B2(G900), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n935), .A2(new_n949), .A3(new_n945), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(G72));
  NOR2_X1   g765(.A1(new_n261), .A2(new_n302), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT127), .Z(new_n953));
  OAI211_X1 g767(.A(new_n926), .B(new_n774), .C1(new_n930), .C2(new_n931), .ZN(new_n954));
  NAND2_X1  g768(.A1(G472), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT63), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT126), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n275), .B(new_n953), .C1(new_n954), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n953), .A2(new_n275), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n937), .A2(new_n774), .A3(new_n940), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n957), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n811), .A2(new_n815), .ZN(new_n962));
  INV_X1    g776(.A(new_n303), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n963), .A2(new_n651), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n962), .A2(new_n956), .A3(new_n964), .ZN(new_n965));
  NOR4_X1   g779(.A1(new_n958), .A2(new_n961), .A3(new_n875), .A4(new_n965), .ZN(G57));
endmodule


