//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AND2_X1   g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G20), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n213), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n216), .B1(new_n218), .B2(new_n219), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT65), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n233), .B(new_n237), .Z(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(G41), .ZN(new_n246));
  INV_X1    g0046(.A(G45), .ZN(new_n247));
  AOI21_X1  g0047(.A(G1), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(G33), .A2(G41), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G1), .A3(G13), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(new_n250), .A3(G274), .ZN(new_n251));
  INV_X1    g0051(.A(G226), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n259), .A2(G223), .B1(new_n262), .B2(G77), .ZN(new_n263));
  INV_X1    g0063(.A(G222), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n258), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n256), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n263), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n250), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n255), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G1), .A2(G13), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n211), .A2(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(G150), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n204), .A2(G20), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n272), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n210), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G50), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(G50), .B2(new_n281), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n269), .A2(G169), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n269), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n280), .A2(new_n286), .ZN(new_n291));
  XOR2_X1   g0091(.A(new_n291), .B(KEYINPUT9), .Z(new_n292));
  NAND2_X1  g0092(.A1(new_n269), .A2(G190), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n269), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n282), .A2(new_n203), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n277), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n302));
  INV_X1    g0102(.A(G77), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n302), .B1(new_n303), .B2(new_n275), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(KEYINPUT11), .A3(new_n272), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n283), .A2(G68), .A3(new_n284), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(KEYINPUT11), .B1(new_n304), .B2(new_n272), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n252), .A2(new_n256), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n230), .A2(G1698), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n260), .C2(new_n261), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G97), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT67), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT67), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(new_n318), .A3(new_n315), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n268), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT13), .ZN(new_n321));
  INV_X1    g0121(.A(G238), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n251), .B1(new_n322), .B2(new_n254), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n320), .B2(new_n324), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n311), .B(G169), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n320), .A2(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n320), .A2(new_n321), .A3(new_n324), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(G179), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n330), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n311), .B1(new_n333), .B2(G169), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n310), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G200), .B1(new_n325), .B2(new_n326), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n329), .A2(G190), .A3(new_n330), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n336), .A2(new_n337), .A3(new_n309), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n274), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT66), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT15), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(G87), .ZN(new_n346));
  INV_X1    g0146(.A(G87), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(KEYINPUT15), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT66), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n344), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n341), .B1(new_n350), .B2(new_n275), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n272), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n303), .B1(new_n210), .B2(G20), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n283), .A2(new_n353), .B1(new_n303), .B2(new_n282), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n259), .A2(G238), .B1(new_n262), .B2(G107), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n230), .B2(new_n266), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n268), .ZN(new_n359));
  INV_X1    g0159(.A(new_n254), .ZN(new_n360));
  INV_X1    g0160(.A(G274), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n217), .B2(new_n249), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n360), .A2(G244), .B1(new_n362), .B2(new_n248), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n355), .B1(new_n356), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(new_n288), .A3(new_n363), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n355), .C1(new_n369), .C2(new_n364), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n299), .A2(new_n335), .A3(new_n339), .A4(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n283), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n340), .A2(new_n284), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(new_n281), .B2(new_n340), .ZN(new_n375));
  XNOR2_X1  g0175(.A(G58), .B(G68), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n377));
  NOR3_X1   g0177(.A1(new_n260), .A2(new_n261), .A3(G20), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT68), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT7), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT69), .B1(new_n378), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n257), .A2(new_n211), .A3(new_n258), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT69), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT68), .B(KEYINPUT7), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n257), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n258), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT70), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT70), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n262), .A2(new_n391), .A3(KEYINPUT7), .A4(new_n211), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n384), .A2(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n377), .B1(new_n393), .B2(new_n203), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G68), .B1(new_n378), .B2(new_n379), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n385), .A2(new_n383), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT16), .B(new_n377), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n272), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n375), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT71), .ZN(new_n403));
  OR2_X1    g0203(.A1(G223), .A2(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n252), .A2(G1698), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n404), .B(new_n405), .C1(new_n260), .C2(new_n261), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n268), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n250), .A2(G232), .A3(new_n253), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n251), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n411), .A3(new_n288), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n250), .B1(new_n406), .B2(new_n407), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n251), .A2(new_n410), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n356), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n403), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n412), .A2(new_n403), .A3(new_n415), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT18), .B1(new_n402), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n375), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n413), .A2(new_n414), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n369), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G200), .B2(new_n422), .ZN(new_n424));
  AND3_X1   g0224(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n390), .A2(new_n392), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT16), .B1(new_n429), .B2(new_n377), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n421), .B(new_n424), .C1(new_n430), .C2(new_n400), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g0233(.A1(new_n412), .A2(new_n403), .A3(new_n415), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n416), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n400), .B1(new_n394), .B2(new_n395), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n435), .B(new_n436), .C1(new_n437), .C2(new_n375), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n396), .A2(new_n401), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(KEYINPUT17), .A3(new_n421), .A4(new_n424), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n420), .A2(new_n433), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n372), .A2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(G257), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n257), .A2(G303), .A3(new_n258), .ZN(new_n444));
  OAI211_X1 g0244(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT75), .B1(new_n259), .B2(G264), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n268), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n210), .B(G45), .C1(new_n246), .C2(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT74), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT5), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G41), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT74), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n210), .A4(G45), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n452), .A2(G41), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n451), .A2(new_n455), .A3(new_n362), .A4(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G270), .B(new_n250), .C1(new_n450), .C2(new_n456), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n449), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G20), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n272), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n463), .A2(KEYINPUT20), .A3(new_n272), .A4(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n210), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n281), .A2(new_n471), .A3(new_n271), .A4(new_n270), .ZN(new_n472));
  MUX2_X1   g0272(.A(new_n281), .B(new_n472), .S(G116), .Z(new_n473));
  AOI21_X1  g0273(.A(new_n356), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n461), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT21), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT76), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT76), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n461), .A2(new_n474), .A3(new_n478), .A4(KEYINPUT21), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n461), .A2(G200), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n470), .A2(new_n473), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(new_n482), .C1(new_n369), .C2(new_n461), .ZN(new_n483));
  INV_X1    g0283(.A(new_n461), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n288), .B1(new_n470), .B2(new_n473), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n475), .A2(new_n476), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n480), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G257), .B(new_n250), .C1(new_n450), .C2(new_n456), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n458), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n462), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G250), .A2(G1698), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT4), .A2(G244), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n494), .B1(new_n495), .B2(G1698), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n265), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n250), .B1(new_n498), .B2(KEYINPUT73), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT73), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n492), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n288), .B(new_n489), .C1(new_n499), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n498), .A2(KEYINPUT73), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n268), .A3(new_n501), .ZN(new_n504));
  INV_X1    g0304(.A(new_n489), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n356), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(G107), .B1(new_n427), .B2(new_n428), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n508));
  XOR2_X1   g0308(.A(G97), .B(G107), .Z(new_n509));
  OAI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(G20), .B1(G77), .B2(new_n277), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n273), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n472), .A2(KEYINPUT72), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n472), .A2(KEYINPUT72), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(G97), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G97), .B2(new_n281), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n502), .A2(new_n506), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n511), .B1(new_n393), .B2(new_n207), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(new_n272), .ZN(new_n519));
  AOI211_X1 g0319(.A(G190), .B(new_n489), .C1(new_n499), .C2(new_n501), .ZN(new_n520));
  AOI21_X1  g0320(.A(G200), .B1(new_n504), .B2(new_n505), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G264), .B(new_n250), .C1(new_n450), .C2(new_n456), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n526));
  OAI211_X1 g0326(.A(G250), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n527));
  INV_X1    g0327(.A(G33), .ZN(new_n528));
  AND2_X1   g0328(.A1(KEYINPUT77), .A2(G294), .ZN(new_n529));
  NOR2_X1   g0329(.A1(KEYINPUT77), .A2(G294), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n525), .B1(new_n532), .B2(new_n268), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n288), .A3(new_n458), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n458), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n356), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n211), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT22), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT22), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n265), .A2(new_n539), .A3(new_n211), .A4(G87), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n528), .A2(new_n464), .A3(G20), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT23), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n211), .B2(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT24), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT24), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n541), .A2(new_n549), .A3(new_n546), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n273), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n513), .A2(G107), .A3(new_n514), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n281), .A2(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT25), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n534), .B(new_n536), .C1(new_n551), .C2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n211), .B1(new_n315), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G87), .B2(new_n208), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n211), .B(G68), .C1(new_n260), .C2(new_n261), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n275), .B2(new_n206), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n272), .B1(new_n350), .B2(new_n282), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n513), .A2(G87), .A3(new_n514), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G250), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n247), .B2(G1), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n210), .A2(new_n361), .A3(G45), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n250), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G244), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n571));
  OAI211_X1 g0371(.A(G238), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n528), .C2(new_n464), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n369), .B(new_n570), .C1(new_n573), .C2(new_n268), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n570), .B1(new_n573), .B2(new_n268), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  INV_X1    g0378(.A(new_n350), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(new_n513), .A3(new_n514), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n563), .A2(new_n580), .B1(new_n576), .B2(new_n288), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n577), .A2(new_n356), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n575), .A2(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n550), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n549), .B1(new_n541), .B2(new_n546), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n272), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n555), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n533), .A2(new_n369), .A3(new_n458), .ZN(new_n588));
  AOI21_X1  g0388(.A(G200), .B1(new_n533), .B2(new_n458), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n556), .A2(new_n583), .A3(new_n590), .ZN(new_n591));
  AND4_X1   g0391(.A1(new_n442), .A2(new_n487), .A3(new_n523), .A4(new_n591), .ZN(G372));
  INV_X1    g0392(.A(KEYINPUT78), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n573), .A2(new_n593), .A3(new_n268), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n573), .B2(new_n268), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n569), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n356), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(G200), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n581), .A2(new_n597), .B1(new_n598), .B2(new_n575), .ZN(new_n599));
  INV_X1    g0399(.A(new_n519), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n504), .A2(G179), .A3(new_n505), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n489), .B1(new_n499), .B2(new_n501), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(KEYINPUT79), .C1(new_n356), .C2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT79), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n502), .B2(new_n506), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n599), .A2(new_n600), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT26), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n601), .B1(new_n356), .B2(new_n602), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n583), .A2(KEYINPUT26), .A3(new_n609), .A4(new_n600), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n597), .A2(new_n581), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n598), .A2(new_n575), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n517), .A2(new_n522), .A3(new_n590), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n480), .A2(new_n556), .A3(new_n486), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n442), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n335), .A2(new_n367), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n339), .A2(new_n433), .A3(new_n440), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n420), .B(new_n438), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n297), .A2(new_n298), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n290), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n619), .A2(new_n624), .ZN(G369));
  NAND3_X1  g0425(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT80), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT27), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(G213), .ZN(new_n631));
  INV_X1    g0431(.A(G343), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n482), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n487), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n480), .A2(new_n486), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(new_n636), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(G330), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n556), .A2(new_n590), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n586), .A2(new_n587), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n644), .B2(new_n634), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n556), .B2(new_n634), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n556), .A2(new_n633), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n638), .A2(new_n633), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n642), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(G399));
  INV_X1    g0451(.A(new_n214), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(G41), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n210), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n347), .A2(new_n206), .A3(new_n207), .A4(new_n464), .ZN(new_n656));
  INV_X1    g0456(.A(new_n653), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n655), .A2(new_n656), .B1(new_n219), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT28), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT29), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n519), .B1(new_n609), .B2(new_n604), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(KEYINPUT26), .A3(new_n599), .A4(new_n603), .ZN(new_n662));
  INV_X1    g0462(.A(new_n583), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n607), .B1(new_n663), .B2(new_n517), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n616), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n517), .A2(new_n522), .A3(new_n590), .A4(new_n614), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n612), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n634), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT82), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n662), .A2(new_n664), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n617), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT82), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(new_n673), .A3(new_n634), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n660), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n633), .B1(new_n611), .B2(new_n617), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT83), .B1(new_n676), .B2(KEYINPUT29), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n487), .A2(new_n523), .A3(new_n591), .A4(new_n634), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT30), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n533), .A2(new_n449), .A3(new_n576), .A4(new_n460), .ZN(new_n681));
  OAI211_X1 g0481(.A(KEYINPUT81), .B(new_n680), .C1(new_n601), .C2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n504), .A2(new_n505), .ZN(new_n683));
  AOI21_X1  g0483(.A(G179), .B1(new_n449), .B2(new_n460), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n683), .A2(new_n535), .A3(new_n596), .A4(new_n684), .ZN(new_n685));
  AND4_X1   g0485(.A1(new_n449), .A2(new_n533), .A3(new_n576), .A4(new_n460), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n680), .A2(KEYINPUT81), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(G179), .A3(new_n602), .A4(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n633), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n633), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n679), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT83), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n673), .B1(new_n672), .B2(new_n634), .ZN(new_n697));
  AOI211_X1 g0497(.A(KEYINPUT82), .B(new_n633), .C1(new_n617), .C2(new_n671), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n696), .B(KEYINPUT29), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n678), .A2(new_n695), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n659), .B1(new_n701), .B2(G1), .ZN(G364));
  NAND2_X1  g0502(.A1(new_n211), .A2(G13), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT84), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G45), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n654), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n641), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(G330), .B2(new_n639), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n652), .A2(new_n262), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G355), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G116), .B2(new_n214), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n652), .A2(new_n265), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n219), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n247), .B2(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n241), .A2(new_n247), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(G13), .A2(G33), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n271), .B1(G20), .B2(new_n356), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n707), .B1(new_n718), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n211), .A2(new_n288), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G200), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT86), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(new_n369), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(G190), .ZN(new_n730));
  XNOR2_X1  g0530(.A(KEYINPUT33), .B(G317), .ZN(new_n731));
  AOI22_X1  g0531(.A1(G326), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n211), .A2(G179), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G190), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G329), .ZN(new_n737));
  INV_X1    g0537(.A(new_n726), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n369), .A3(G200), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G322), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n262), .B(new_n737), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n726), .A2(KEYINPUT85), .A3(new_n734), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT85), .B1(new_n726), .B2(new_n734), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n742), .B1(new_n746), .B2(G311), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n369), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n211), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n733), .A2(new_n369), .A3(G200), .ZN(new_n750));
  INV_X1    g0550(.A(G283), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n749), .A2(new_n531), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n733), .A2(G190), .A3(G200), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n752), .B1(G303), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n732), .A2(new_n747), .A3(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n749), .A2(new_n206), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n262), .B(new_n757), .C1(G58), .C2(new_n739), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n754), .A2(G87), .ZN(new_n759));
  INV_X1    g0559(.A(G159), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT32), .B1(new_n735), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n735), .A2(KEYINPUT32), .A3(new_n760), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n750), .A2(new_n207), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n746), .A2(G77), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n758), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n729), .ZN(new_n768));
  INV_X1    g0568(.A(new_n730), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n201), .A2(new_n768), .B1(new_n769), .B2(new_n203), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n756), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n725), .B1(new_n771), .B2(new_n722), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n721), .B(KEYINPUT87), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n639), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n709), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(G396));
  INV_X1    g0576(.A(new_n355), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n633), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n370), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n367), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n365), .A2(new_n366), .A3(new_n634), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT89), .Z(new_n783));
  INV_X1    g0583(.A(new_n782), .ZN(new_n784));
  MUX2_X1   g0584(.A(new_n783), .B(new_n784), .S(new_n676), .Z(new_n785));
  AOI21_X1  g0585(.A(new_n707), .B1(new_n785), .B2(new_n695), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n695), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n722), .A2(new_n719), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n706), .B1(new_n303), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  INV_X1    g0590(.A(G294), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n262), .B1(new_n735), .B2(new_n790), .C1(new_n740), .C2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n746), .B2(G116), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G283), .A2(new_n730), .B1(new_n729), .B2(G303), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n750), .A2(new_n347), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n795), .B(new_n757), .C1(G107), .C2(new_n754), .ZN(new_n796));
  AND3_X1   g0596(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n746), .A2(G159), .B1(G143), .B2(new_n739), .ZN(new_n798));
  INV_X1    g0598(.A(G150), .ZN(new_n799));
  INV_X1    g0599(.A(G137), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n798), .B1(new_n769), .B2(new_n799), .C1(new_n800), .C2(new_n768), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n265), .B1(new_n735), .B2(new_n803), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n201), .A2(new_n753), .B1(new_n750), .B2(new_n203), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT88), .Z(new_n806));
  INV_X1    g0606(.A(new_n749), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n804), .B(new_n806), .C1(G58), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n797), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n722), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n789), .B1(new_n809), .B2(new_n810), .C1(new_n720), .C2(new_n784), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n787), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(G384));
  NOR2_X1   g0613(.A1(new_n704), .A2(new_n210), .ZN(new_n814));
  INV_X1    g0614(.A(G330), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n690), .A2(KEYINPUT93), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT93), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n689), .A2(new_n817), .A3(KEYINPUT31), .A4(new_n633), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n679), .A2(new_n816), .A3(new_n693), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n310), .A2(new_n633), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n335), .A2(new_n339), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(G169), .B1(new_n325), .B2(new_n326), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT14), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n823), .A2(new_n331), .A3(new_n327), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n310), .B(new_n633), .C1(new_n824), .C2(new_n338), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n782), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n377), .B1(new_n397), .B2(new_n398), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n395), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n375), .B1(new_n401), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n830), .A2(new_n631), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT37), .ZN(new_n832));
  INV_X1    g0632(.A(new_n631), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n400), .B1(new_n395), .B2(new_n828), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n435), .A2(new_n833), .B1(new_n834), .B2(new_n375), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n832), .B1(new_n835), .B2(new_n431), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT91), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n441), .A2(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n830), .B1(new_n419), .B2(new_n631), .ZN(new_n839));
  INV_X1    g0639(.A(new_n424), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n437), .A2(new_n840), .A3(new_n375), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT37), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n435), .B1(new_n437), .B2(new_n375), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n833), .B1(new_n437), .B2(new_n375), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n844), .A3(new_n431), .A4(new_n832), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n842), .A2(KEYINPUT91), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n838), .A2(KEYINPUT38), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n441), .A2(new_n831), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n836), .A2(new_n837), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n827), .B1(new_n847), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT94), .B1(new_n853), .B2(KEYINPUT40), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n843), .A2(new_n844), .A3(new_n431), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT92), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n856), .A2(new_n857), .A3(new_n845), .ZN(new_n858));
  INV_X1    g0658(.A(new_n844), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n441), .A2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n858), .B(new_n860), .C1(new_n857), .C2(new_n856), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n851), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(new_n847), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n827), .A2(KEYINPUT95), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT95), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n819), .A2(new_n826), .A3(new_n865), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT40), .A4(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n854), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT94), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT40), .ZN(new_n870));
  AND4_X1   g0670(.A1(KEYINPUT38), .A2(new_n848), .A3(new_n846), .A4(new_n849), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n838), .B2(new_n846), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n869), .B(new_n870), .C1(new_n873), .C2(new_n827), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT96), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n442), .A2(new_n819), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n815), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n699), .B1(new_n675), .B2(new_n677), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n442), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n624), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n833), .B1(new_n420), .B2(new_n438), .ZN(new_n883));
  INV_X1    g0683(.A(new_n873), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n821), .A2(new_n825), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n618), .A2(new_n634), .A3(new_n784), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n781), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n883), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n891), .A2(KEYINPUT92), .B1(new_n441), .B2(new_n859), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n892), .B2(new_n858), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n890), .B1(new_n893), .B2(new_n871), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n824), .A2(new_n310), .A3(new_n634), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n852), .A2(KEYINPUT39), .A3(new_n847), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n889), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n882), .B(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n814), .B1(new_n879), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n900), .B2(new_n879), .ZN(new_n902));
  OAI21_X1  g0702(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n903), .A2(new_n219), .B1(G50), .B2(new_n203), .ZN(new_n904));
  INV_X1    g0704(.A(G13), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n904), .A2(G1), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT90), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n464), .B(new_n218), .C1(new_n510), .C2(KEYINPUT35), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(KEYINPUT35), .B2(new_n510), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT36), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n910), .B2(new_n909), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n902), .A2(new_n912), .ZN(G367));
  INV_X1    g0713(.A(new_n647), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n523), .B1(new_n519), .B2(new_n634), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n661), .A2(new_n603), .A3(new_n633), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT99), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n917), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n517), .B1(new_n922), .B2(new_n556), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n634), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n642), .A3(new_n649), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(KEYINPUT97), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n633), .A2(new_n565), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n599), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n612), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n927), .A2(KEYINPUT97), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT98), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n930), .A2(new_n935), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n933), .B(KEYINPUT43), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n914), .A2(KEYINPUT99), .A3(new_n917), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n921), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n653), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n650), .A2(new_n917), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT45), .Z(new_n949));
  NOR2_X1   g0749(.A1(new_n650), .A2(new_n917), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n647), .A2(KEYINPUT100), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n952), .B(new_n953), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n649), .A2(new_n642), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n646), .B2(new_n649), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n641), .B1(KEYINPUT101), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(KEYINPUT101), .B2(new_n956), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT102), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT102), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n956), .A2(new_n640), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n954), .A2(new_n700), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n947), .B1(new_n963), .B2(new_n700), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n705), .A2(G1), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT103), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n942), .A2(new_n919), .A3(new_n918), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n945), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(KEYINPUT104), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT104), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n945), .A2(new_n972), .A3(new_n968), .A4(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n237), .A2(new_n713), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n723), .B1(new_n350), .B2(new_n214), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n707), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G143), .A2(new_n729), .B1(new_n730), .B2(G159), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n202), .A2(new_n753), .B1(new_n750), .B2(new_n303), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G68), .B2(new_n807), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n746), .A2(G50), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n265), .B1(new_n735), .B2(new_n800), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n739), .B2(G150), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n749), .A2(new_n207), .B1(new_n750), .B2(new_n206), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n265), .B1(new_n739), .B2(G303), .ZN(new_n986));
  XNOR2_X1  g0786(.A(KEYINPUT106), .B(G317), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n986), .B1(new_n735), .B2(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n985), .B(new_n988), .C1(G283), .C2(new_n746), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n754), .A2(KEYINPUT46), .A3(G116), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n753), .B2(new_n464), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(new_n769), .C2(new_n531), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n989), .B1(KEYINPUT105), .B2(new_n993), .C1(new_n790), .C2(new_n768), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n993), .A2(KEYINPUT105), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n984), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n977), .B1(new_n997), .B2(new_n722), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n933), .A2(new_n773), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n974), .A2(new_n1000), .ZN(G387));
  INV_X1    g0801(.A(new_n962), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n701), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n962), .A2(new_n700), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1003), .A2(new_n653), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n646), .A2(new_n773), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n710), .A2(new_n656), .B1(new_n207), .B2(new_n652), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n233), .A2(new_n247), .ZN(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n656), .C1(G68), .C2(G77), .ZN(new_n1009));
  XOR2_X1   g0809(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n1010));
  OR3_X1    g0810(.A1(new_n1010), .A2(G50), .A3(new_n274), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(G50), .B2(new_n274), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n713), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1007), .B1(new_n1008), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n723), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n707), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n730), .A2(new_n340), .B1(G68), .B2(new_n746), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT108), .Z(new_n1019));
  OAI221_X1 g0819(.A(new_n265), .B1(new_n735), .B2(new_n799), .C1(new_n740), .C2(new_n201), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n750), .A2(new_n206), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n350), .A2(new_n749), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n753), .A2(new_n303), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1019), .B(new_n1024), .C1(new_n760), .C2(new_n768), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n265), .B1(new_n736), .B2(G326), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n749), .A2(new_n751), .B1(new_n753), .B2(new_n531), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n987), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n746), .A2(G303), .B1(new_n739), .B2(new_n1028), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n769), .B2(new_n790), .C1(new_n741), .C2(new_n768), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT48), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1026), .B1(new_n464), .B2(new_n750), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1025), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1006), .B(new_n1017), .C1(new_n1037), .C2(new_n722), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n1002), .B2(new_n966), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1005), .A2(new_n1039), .ZN(G393));
  NAND2_X1  g0840(.A1(new_n922), .A2(new_n721), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n729), .A2(G150), .B1(G159), .B2(new_n739), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT51), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n807), .A2(G77), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n203), .B2(new_n753), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n736), .A2(G143), .ZN(new_n1046));
  NOR4_X1   g0846(.A1(new_n1045), .A2(new_n262), .A3(new_n795), .A4(new_n1046), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n201), .B2(new_n769), .C1(new_n274), .C2(new_n745), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n729), .A2(G317), .B1(G311), .B2(new_n739), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT52), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n730), .A2(G303), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n746), .A2(G294), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n265), .B(new_n764), .C1(G322), .C2(new_n736), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n807), .A2(G116), .B1(new_n754), .B2(G283), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1043), .A2(new_n1048), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n722), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n723), .B1(new_n206), .B2(new_n214), .C1(new_n714), .C2(new_n244), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1041), .A2(new_n707), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n952), .B(new_n647), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n1060), .A2(KEYINPUT109), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n966), .B1(new_n1060), .B2(KEYINPUT109), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT110), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n963), .A2(new_n657), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1060), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1003), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G390));
  NAND2_X1  g0873(.A1(new_n894), .A2(new_n897), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n719), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n265), .B1(new_n739), .B2(G116), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n759), .A3(new_n1044), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n750), .A2(new_n203), .B1(new_n735), .B2(new_n791), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT117), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1079), .B1(new_n769), .B2(new_n207), .C1(new_n751), .C2(new_n768), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(G97), .C2(new_n746), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n749), .A2(new_n760), .B1(new_n750), .B2(new_n201), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n265), .B1(new_n740), .B2(new_n803), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1082), .B(new_n1083), .C1(G125), .C2(new_n736), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n729), .A2(G128), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n753), .A2(new_n799), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT53), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT54), .B(G143), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT115), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n730), .A2(G137), .B1(new_n746), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(KEYINPUT116), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(KEYINPUT116), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1081), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n810), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n706), .B(new_n1096), .C1(new_n274), .C2(new_n788), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1075), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n670), .A2(new_n674), .A3(new_n781), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n780), .A3(new_n885), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n896), .B1(new_n862), .B2(new_n847), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n781), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n676), .B2(new_n784), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n895), .B1(new_n1104), .B2(new_n886), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1074), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n819), .A2(new_n826), .A3(G330), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n694), .A2(G330), .A3(new_n784), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1111), .A2(new_n886), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1074), .B2(new_n1105), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT111), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n1102), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1113), .B2(new_n1102), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1110), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1098), .B1(new_n1117), .B2(new_n967), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(KEYINPUT118), .B(new_n1098), .C1(new_n1117), .C2(new_n967), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n819), .A2(G330), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n783), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1112), .B1(new_n1123), .B2(new_n886), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1099), .A2(new_n780), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT113), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1104), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1111), .A2(KEYINPUT112), .A3(new_n886), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1108), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT112), .B1(new_n1111), .B2(new_n886), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1127), .B(new_n1128), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1111), .A2(new_n886), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT112), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n1129), .A3(new_n1108), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1127), .B1(new_n1137), .B2(new_n1128), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1126), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n442), .A2(G330), .A3(new_n819), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n881), .A2(new_n624), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(KEYINPUT114), .B(new_n653), .C1(new_n1117), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1117), .A2(new_n1142), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1113), .A2(new_n1102), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT111), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1113), .A2(new_n1102), .A3(new_n1114), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1149), .A2(new_n1141), .A3(new_n1139), .A4(new_n1110), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT114), .B1(new_n1150), .B2(new_n653), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1120), .B(new_n1121), .C1(new_n1145), .C2(new_n1151), .ZN(G378));
  OAI21_X1  g0952(.A(new_n1128), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT113), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1154), .A2(new_n1132), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1141), .B1(new_n1117), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n854), .A2(new_n874), .A3(new_n867), .A4(G330), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n291), .A2(new_n631), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n299), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n299), .A2(new_n1161), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1162), .A3(new_n1158), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n899), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n868), .A2(G330), .A3(new_n874), .A4(new_n1168), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n899), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1157), .A2(new_n1169), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1156), .A2(new_n1177), .A3(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1156), .B2(new_n1177), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n653), .B(new_n1178), .C1(new_n1179), .C2(KEYINPUT120), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT120), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1181), .B(KEYINPUT57), .C1(new_n1156), .C2(new_n1177), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1169), .A2(new_n719), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n265), .A2(G41), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n751), .B2(new_n735), .C1(new_n740), .C2(new_n207), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n579), .B2(new_n746), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G97), .A2(new_n730), .B1(new_n729), .B2(G116), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n750), .A2(new_n202), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1023), .B(new_n1189), .C1(G68), .C2(new_n807), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1194));
  AOI211_X1 g0994(.A(G50), .B(new_n1185), .C1(new_n528), .C2(new_n246), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G128), .A2(new_n739), .B1(new_n807), .B2(G150), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1090), .A2(new_n754), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(new_n800), .C2(new_n745), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n769), .A2(new_n803), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(G125), .C2(new_n729), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT119), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n736), .C2(G124), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n760), .C2(new_n750), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1202), .A2(KEYINPUT119), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1193), .B(new_n1196), .C1(new_n1205), .C2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1207), .A2(new_n722), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n706), .B(new_n1208), .C1(new_n201), .C2(new_n788), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1177), .A2(new_n966), .B1(new_n1184), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1183), .A2(new_n1210), .ZN(G375));
  NAND3_X1  g1011(.A1(new_n881), .A2(new_n624), .A3(new_n1140), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1155), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1142), .A2(new_n1213), .A3(new_n947), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n886), .A2(new_n719), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1022), .B1(G283), .B2(new_n739), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT121), .Z(new_n1217));
  AOI21_X1  g1017(.A(new_n265), .B1(new_n736), .B2(G303), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n303), .B2(new_n750), .C1(new_n206), .C2(new_n753), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G107), .B2(new_n746), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G116), .A2(new_n730), .B1(new_n729), .B2(G294), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1217), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n262), .B1(new_n736), .B2(G128), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n740), .B2(new_n800), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n746), .B2(G150), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n729), .A2(G132), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n730), .A2(new_n1090), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n753), .A2(new_n760), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1189), .B(new_n1228), .C1(G50), .C2(new_n807), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n810), .B1(new_n1222), .B2(new_n1230), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n706), .B(new_n1231), .C1(new_n203), .C2(new_n788), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1139), .A2(new_n966), .B1(new_n1215), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1214), .A2(new_n1233), .ZN(G381));
  INV_X1    g1034(.A(KEYINPUT123), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1005), .A2(new_n775), .A3(new_n1039), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1072), .A2(new_n812), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(G387), .A2(G381), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(G375), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1118), .ZN(new_n1242));
  OAI211_X1 g1042(.A(KEYINPUT122), .B(new_n1242), .C1(new_n1145), .C2(new_n1151), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n653), .B1(new_n1117), .B2(new_n1142), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT114), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(new_n1144), .A3(new_n1143), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT122), .B1(new_n1248), .B2(new_n1242), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1235), .B1(new_n1241), .B2(new_n1251), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n1240), .A2(KEYINPUT123), .A3(new_n1250), .ZN(new_n1253));
  OR2_X1    g1053(.A1(new_n1252), .A2(new_n1253), .ZN(G407));
  INV_X1    g1054(.A(G213), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1239), .A2(new_n632), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1255), .B1(new_n1257), .B2(new_n1251), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1252), .B2(new_n1253), .ZN(G409));
  OAI21_X1  g1059(.A(KEYINPUT60), .B1(new_n1155), .B2(new_n1212), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1213), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1155), .A2(KEYINPUT60), .A3(new_n1212), .ZN(new_n1262));
  AND4_X1   g1062(.A1(KEYINPUT124), .A2(new_n1261), .A3(new_n653), .A4(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n657), .B1(new_n1260), .B2(new_n1213), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT124), .B1(new_n1264), .B2(new_n1262), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1233), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n812), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G384), .B(new_n1233), .C1(new_n1263), .C2(new_n1265), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1255), .A2(G343), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1270), .A2(KEYINPUT125), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1269), .A2(G2897), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1267), .A2(new_n1268), .A3(new_n1273), .A4(new_n1271), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(G378), .B(new_n1210), .C1(new_n1180), .C2(new_n1182), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1156), .A2(new_n1177), .A3(new_n947), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1210), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1242), .B1(new_n1145), .B2(new_n1151), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT122), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1285), .B2(new_n1243), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1270), .B1(new_n1279), .B2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1281), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1278), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(KEYINPUT126), .A3(new_n1270), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1277), .B1(new_n1289), .B2(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT127), .B1(new_n1293), .B2(KEYINPUT61), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT126), .B1(new_n1291), .B2(new_n1270), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n1288), .B(new_n1269), .C1(new_n1290), .C2(new_n1278), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1295), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1291), .A2(new_n1302), .A3(new_n1270), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1289), .A2(new_n1302), .A3(new_n1292), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1304), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1294), .A2(new_n1301), .A3(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G390), .B1(new_n974), .B2(new_n1000), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G393), .A2(G396), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1311), .A2(new_n1236), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n974), .A2(new_n1000), .A3(G390), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1312), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n974), .A2(new_n1000), .A3(G390), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1315), .B1(new_n1316), .B2(new_n1309), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1308), .A2(new_n1318), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(KEYINPUT61), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1289), .A2(new_n1292), .A3(KEYINPUT63), .A4(new_n1302), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1295), .A2(new_n1287), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1303), .A2(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .A4(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1319), .A2(new_n1325), .ZN(G405));
  NAND2_X1  g1126(.A1(new_n1251), .A2(G375), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1278), .ZN(new_n1328));
  XNOR2_X1  g1128(.A(new_n1328), .B(new_n1302), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(new_n1329), .B(new_n1318), .ZN(G402));
endmodule


