

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  NOR2_X1 U323 ( .A1(n388), .A2(n387), .ZN(n389) );
  INV_X1 U324 ( .A(n485), .ZN(n446) );
  XOR2_X1 U325 ( .A(KEYINPUT100), .B(n449), .Z(n498) );
  XOR2_X1 U326 ( .A(KEYINPUT28), .B(n471), .Z(n520) );
  XNOR2_X1 U327 ( .A(n362), .B(n361), .ZN(n514) );
  AND2_X1 U328 ( .A1(G230GAT), .A2(G233GAT), .ZN(n291) );
  INV_X1 U329 ( .A(KEYINPUT117), .ZN(n467) );
  INV_X1 U330 ( .A(KEYINPUT6), .ZN(n346) );
  XNOR2_X1 U331 ( .A(n467), .B(KEYINPUT54), .ZN(n468) );
  XNOR2_X1 U332 ( .A(n437), .B(n291), .ZN(n438) );
  XNOR2_X1 U333 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U334 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U335 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U336 ( .A(n349), .B(n348), .ZN(n352) );
  INV_X1 U337 ( .A(KEYINPUT37), .ZN(n412) );
  OR2_X1 U338 ( .A1(n513), .A2(n446), .ZN(n447) );
  XNOR2_X1 U339 ( .A(n413), .B(n412), .ZN(n513) );
  AND2_X1 U340 ( .A1(n475), .A2(n525), .ZN(n561) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n450) );
  XOR2_X1 U342 ( .A(n376), .B(n375), .Z(n525) );
  XNOR2_X1 U343 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U344 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U345 ( .A(n479), .B(n478), .ZN(G1351GAT) );
  XNOR2_X1 U346 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT101), .B(KEYINPUT38), .Z(n448) );
  XOR2_X1 U348 ( .A(G211GAT), .B(G155GAT), .Z(n293) );
  XNOR2_X1 U349 ( .A(G183GAT), .B(G71GAT), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U351 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n432) );
  XOR2_X1 U352 ( .A(n294), .B(n432), .Z(n296) );
  XNOR2_X1 U353 ( .A(G22GAT), .B(G78GAT), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n298) );
  NAND2_X1 U356 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U358 ( .A(n299), .B(KEYINPUT80), .Z(n307) );
  XOR2_X1 U359 ( .A(G64GAT), .B(G127GAT), .Z(n301) );
  XNOR2_X1 U360 ( .A(G15GAT), .B(G8GAT), .ZN(n300) );
  XNOR2_X1 U361 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U362 ( .A(KEYINPUT12), .B(KEYINPUT79), .Z(n303) );
  XNOR2_X1 U363 ( .A(G1GAT), .B(G57GAT), .ZN(n302) );
  XNOR2_X1 U364 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U366 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U367 ( .A(n309), .B(n308), .Z(n580) );
  INV_X1 U368 ( .A(n580), .ZN(n459) );
  XNOR2_X1 U369 ( .A(KEYINPUT88), .B(KEYINPUT87), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n310), .B(KEYINPUT3), .ZN(n311) );
  XOR2_X1 U371 ( .A(n311), .B(KEYINPUT2), .Z(n313) );
  XNOR2_X1 U372 ( .A(G155GAT), .B(G162GAT), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n360) );
  XOR2_X1 U374 ( .A(KEYINPUT89), .B(G204GAT), .Z(n315) );
  XNOR2_X1 U375 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n318) );
  XOR2_X1 U377 ( .A(G78GAT), .B(G148GAT), .Z(n317) );
  XNOR2_X1 U378 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n442) );
  XOR2_X1 U380 ( .A(n318), .B(n442), .Z(n327) );
  XOR2_X1 U381 ( .A(KEYINPUT21), .B(G218GAT), .Z(n320) );
  XNOR2_X1 U382 ( .A(KEYINPUT86), .B(G211GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U384 ( .A(G197GAT), .B(n321), .Z(n340) );
  XNOR2_X1 U385 ( .A(G50GAT), .B(G22GAT), .ZN(n322) );
  XNOR2_X1 U386 ( .A(n322), .B(G141GAT), .ZN(n424) );
  XOR2_X1 U387 ( .A(n424), .B(KEYINPUT24), .Z(n324) );
  NAND2_X1 U388 ( .A1(G228GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n340), .B(n325), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n360), .B(n328), .ZN(n471) );
  INV_X1 U393 ( .A(n520), .ZN(n364) );
  XOR2_X1 U394 ( .A(G36GAT), .B(G8GAT), .Z(n417) );
  XOR2_X1 U395 ( .A(KEYINPUT93), .B(n417), .Z(n330) );
  NAND2_X1 U396 ( .A1(G226GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U398 ( .A(KEYINPUT76), .B(G64GAT), .Z(n332) );
  XNOR2_X1 U399 ( .A(G204GAT), .B(G92GAT), .ZN(n331) );
  XNOR2_X1 U400 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U401 ( .A(G176GAT), .B(n333), .Z(n440) );
  XOR2_X1 U402 ( .A(n334), .B(n440), .Z(n342) );
  XOR2_X1 U403 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n336) );
  XNOR2_X1 U404 ( .A(G190GAT), .B(KEYINPUT82), .ZN(n335) );
  XNOR2_X1 U405 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U406 ( .A(n337), .B(KEYINPUT19), .Z(n339) );
  XNOR2_X1 U407 ( .A(G169GAT), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U408 ( .A(n339), .B(n338), .ZN(n374) );
  XNOR2_X1 U409 ( .A(n374), .B(n340), .ZN(n341) );
  XNOR2_X1 U410 ( .A(n342), .B(n341), .ZN(n517) );
  XNOR2_X1 U411 ( .A(n517), .B(KEYINPUT27), .ZN(n383) );
  XOR2_X1 U412 ( .A(G85GAT), .B(G57GAT), .Z(n431) );
  XOR2_X1 U413 ( .A(KEYINPUT78), .B(G148GAT), .Z(n344) );
  XNOR2_X1 U414 ( .A(G29GAT), .B(G141GAT), .ZN(n343) );
  XNOR2_X1 U415 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U416 ( .A(n431), .B(n345), .Z(n349) );
  NAND2_X1 U417 ( .A1(G225GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U418 ( .A(G134GAT), .B(G127GAT), .ZN(n350) );
  XNOR2_X1 U419 ( .A(n350), .B(KEYINPUT0), .ZN(n371) );
  XNOR2_X1 U420 ( .A(n371), .B(KEYINPUT4), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U422 ( .A(KEYINPUT92), .B(G120GAT), .Z(n354) );
  XNOR2_X1 U423 ( .A(G113GAT), .B(G1GAT), .ZN(n353) );
  XNOR2_X1 U424 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n362) );
  XOR2_X1 U426 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n358) );
  XNOR2_X1 U427 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n357) );
  XNOR2_X1 U428 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U429 ( .A(n360), .B(n359), .Z(n361) );
  NAND2_X1 U430 ( .A1(n383), .A2(n514), .ZN(n363) );
  XOR2_X1 U431 ( .A(KEYINPUT94), .B(n363), .Z(n539) );
  NAND2_X1 U432 ( .A1(n364), .A2(n539), .ZN(n527) );
  XOR2_X1 U433 ( .A(G176GAT), .B(KEYINPUT83), .Z(n370) );
  XOR2_X1 U434 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n366) );
  NAND2_X1 U435 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n366), .B(n365), .ZN(n368) );
  XNOR2_X1 U437 ( .A(G99GAT), .B(G71GAT), .ZN(n367) );
  XNOR2_X1 U438 ( .A(n367), .B(G120GAT), .ZN(n443) );
  XNOR2_X1 U439 ( .A(n368), .B(n443), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U441 ( .A(n372), .B(n371), .Z(n376) );
  XNOR2_X1 U442 ( .A(G43GAT), .B(G15GAT), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n373), .B(G113GAT), .ZN(n423) );
  XNOR2_X1 U444 ( .A(n423), .B(n374), .ZN(n375) );
  XOR2_X1 U445 ( .A(KEYINPUT85), .B(n525), .Z(n377) );
  NOR2_X1 U446 ( .A1(n527), .A2(n377), .ZN(n388) );
  NAND2_X1 U447 ( .A1(n517), .A2(n525), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n378), .B(KEYINPUT96), .ZN(n379) );
  NAND2_X1 U449 ( .A1(n379), .A2(n471), .ZN(n380) );
  XNOR2_X1 U450 ( .A(n380), .B(KEYINPUT25), .ZN(n385) );
  NOR2_X1 U451 ( .A1(n525), .A2(n471), .ZN(n382) );
  XNOR2_X1 U452 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n382), .B(n381), .ZN(n542) );
  INV_X1 U454 ( .A(n542), .ZN(n570) );
  AND2_X1 U455 ( .A1(n383), .A2(n570), .ZN(n384) );
  NOR2_X1 U456 ( .A1(n385), .A2(n384), .ZN(n386) );
  NOR2_X1 U457 ( .A1(n514), .A2(n386), .ZN(n387) );
  XOR2_X1 U458 ( .A(KEYINPUT97), .B(n389), .Z(n484) );
  XOR2_X1 U459 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n391) );
  XNOR2_X1 U460 ( .A(KEYINPUT8), .B(G29GAT), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U462 ( .A(KEYINPUT7), .B(n392), .Z(n429) );
  INV_X1 U463 ( .A(n429), .ZN(n410) );
  XOR2_X1 U464 ( .A(G106GAT), .B(G162GAT), .Z(n394) );
  XNOR2_X1 U465 ( .A(G134GAT), .B(G99GAT), .ZN(n393) );
  XNOR2_X1 U466 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U467 ( .A(G218GAT), .B(G36GAT), .Z(n396) );
  XNOR2_X1 U468 ( .A(G50GAT), .B(G43GAT), .ZN(n395) );
  XNOR2_X1 U469 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U470 ( .A(n398), .B(n397), .Z(n400) );
  NAND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n400), .B(n399), .ZN(n408) );
  XOR2_X1 U473 ( .A(G85GAT), .B(KEYINPUT78), .Z(n402) );
  XNOR2_X1 U474 ( .A(G190GAT), .B(KEYINPUT64), .ZN(n401) );
  XNOR2_X1 U475 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U476 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n404) );
  XNOR2_X1 U477 ( .A(G92GAT), .B(KEYINPUT11), .ZN(n403) );
  XNOR2_X1 U478 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U479 ( .A(n406), .B(n405), .Z(n407) );
  XNOR2_X1 U480 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U481 ( .A(n410), .B(n409), .Z(n480) );
  INV_X1 U482 ( .A(n480), .ZN(n552) );
  XOR2_X1 U483 ( .A(n552), .B(KEYINPUT36), .Z(n584) );
  NOR2_X1 U484 ( .A1(n484), .A2(n584), .ZN(n411) );
  NAND2_X1 U485 ( .A1(n459), .A2(n411), .ZN(n413) );
  XOR2_X1 U486 ( .A(KEYINPUT66), .B(KEYINPUT30), .Z(n415) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n414) );
  XNOR2_X1 U488 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U489 ( .A(n416), .B(G197GAT), .Z(n419) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U491 ( .A(n419), .B(n418), .ZN(n428) );
  XOR2_X1 U492 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n421) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U494 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U495 ( .A(n422), .B(KEYINPUT29), .Z(n426) );
  XNOR2_X1 U496 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U497 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U498 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U499 ( .A(n430), .B(n429), .Z(n571) );
  INV_X1 U500 ( .A(n571), .ZN(n501) );
  XOR2_X1 U501 ( .A(KEYINPUT71), .B(n501), .Z(n528) );
  XOR2_X1 U502 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n434) );
  XNOR2_X1 U503 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U504 ( .A(n434), .B(n433), .ZN(n439) );
  XOR2_X1 U505 ( .A(KEYINPUT73), .B(KEYINPUT33), .Z(n436) );
  XNOR2_X1 U506 ( .A(KEYINPUT77), .B(KEYINPUT32), .ZN(n435) );
  XNOR2_X1 U507 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U508 ( .A(n441), .B(n440), .Z(n445) );
  XNOR2_X1 U509 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U510 ( .A(n445), .B(n444), .ZN(n576) );
  NOR2_X1 U511 ( .A1(n528), .A2(n576), .ZN(n485) );
  XNOR2_X1 U512 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U513 ( .A1(n498), .A2(n525), .ZN(n453) );
  XOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT102), .Z(n451) );
  XNOR2_X1 U515 ( .A(KEYINPUT116), .B(n517), .ZN(n466) );
  NOR2_X1 U516 ( .A1(n459), .A2(n584), .ZN(n454) );
  XNOR2_X1 U517 ( .A(KEYINPUT45), .B(n454), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n455), .A2(n528), .ZN(n456) );
  NOR2_X1 U519 ( .A1(n576), .A2(n456), .ZN(n457) );
  XOR2_X1 U520 ( .A(KEYINPUT108), .B(n457), .Z(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT41), .B(n576), .Z(n548) );
  NAND2_X1 U522 ( .A1(n548), .A2(n571), .ZN(n458) );
  XNOR2_X1 U523 ( .A(n458), .B(KEYINPUT46), .ZN(n461) );
  AND2_X1 U524 ( .A1(n459), .A2(n480), .ZN(n460) );
  AND2_X1 U525 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U526 ( .A(n462), .B(KEYINPUT47), .ZN(n463) );
  NAND2_X1 U527 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U528 ( .A(n465), .B(KEYINPUT48), .ZN(n540) );
  NAND2_X1 U529 ( .A1(n466), .A2(n540), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n514), .A2(n470), .ZN(n569) );
  NAND2_X1 U531 ( .A1(n569), .A2(n471), .ZN(n473) );
  XOR2_X1 U532 ( .A(KEYINPUT119), .B(KEYINPUT55), .Z(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT118), .B(n474), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n561), .A2(n552), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n477) );
  INV_X1 U537 ( .A(G190GAT), .ZN(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n482) );
  NAND2_X1 U539 ( .A1(n580), .A2(n480), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n502) );
  AND2_X1 U542 ( .A1(n485), .A2(n502), .ZN(n493) );
  NAND2_X1 U543 ( .A1(n493), .A2(n514), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n486), .B(KEYINPUT34), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n493), .A2(n517), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT98), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G8GAT), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U550 ( .A1(n493), .A2(n525), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U552 ( .A(G15GAT), .B(n492), .Z(G1326GAT) );
  NAND2_X1 U553 ( .A1(n520), .A2(n493), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  NAND2_X1 U556 ( .A1(n498), .A2(n514), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n498), .A2(n517), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(G50GAT), .B(KEYINPUT103), .Z(n500) );
  NAND2_X1 U561 ( .A1(n498), .A2(n520), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U563 ( .A(n548), .B(KEYINPUT104), .ZN(n560) );
  NAND2_X1 U564 ( .A1(n501), .A2(n560), .ZN(n512) );
  INV_X1 U565 ( .A(n502), .ZN(n503) );
  NOR2_X1 U566 ( .A1(n512), .A2(n503), .ZN(n509) );
  NAND2_X1 U567 ( .A1(n514), .A2(n509), .ZN(n504) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(n504), .ZN(n505) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n509), .A2(n517), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U572 ( .A(G71GAT), .B(KEYINPUT105), .Z(n508) );
  NAND2_X1 U573 ( .A1(n509), .A2(n525), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U576 ( .A1(n509), .A2(n520), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(KEYINPUT106), .ZN(n516) );
  NOR2_X1 U579 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n514), .A2(n521), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n525), .A2(n521), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT107), .B(KEYINPUT44), .Z(n523) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT109), .Z(n530) );
  NAND2_X1 U591 ( .A1(n540), .A2(n525), .ZN(n526) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n535) );
  INV_X1 U593 ( .A(n528), .ZN(n557) );
  NAND2_X1 U594 ( .A1(n535), .A2(n557), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U597 ( .A1(n535), .A2(n560), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n535), .A2(n580), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT110), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U603 ( .A1(n535), .A2(n552), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  XOR2_X1 U606 ( .A(G141GAT), .B(KEYINPUT111), .Z(n544) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n553) );
  NAND2_X1 U609 ( .A1(n553), .A2(n571), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT113), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT112), .B(n547), .Z(n550) );
  NAND2_X1 U615 ( .A1(n553), .A2(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n580), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  XNOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n559) );
  NAND2_X1 U624 ( .A1(n561), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT57), .Z(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n561), .A2(n580), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n575) );
  XOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT123), .Z(n573) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n583) );
  INV_X1 U638 ( .A(n583), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n581), .A2(n571), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U641 ( .A(n575), .B(n574), .Z(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n578) );
  NAND2_X1 U643 ( .A1(n581), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

