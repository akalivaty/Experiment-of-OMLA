//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT95), .Z(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT13), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT92), .ZN(new_n205));
  INV_X1    g004(.A(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT91), .B(G36gat), .Z(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(G29gat), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(G43gat), .A2(G50gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218));
  NAND2_X1  g017(.A1(G43gat), .A2(G50gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT15), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(new_n214), .B2(KEYINPUT90), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n213), .A2(new_n216), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n220), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT91), .B(G36gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n210), .B(new_n208), .C1(new_n225), .C2(new_n206), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n205), .B1(new_n223), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n224), .B1(new_n215), .B2(new_n226), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n220), .A3(new_n222), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(KEYINPUT92), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT93), .ZN(new_n234));
  INV_X1    g033(.A(G8gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n233), .B2(new_n234), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  OAI22_X1  g039(.A1(new_n237), .A2(new_n238), .B1(new_n240), .B2(G1gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n238), .ZN(new_n242));
  AOI21_X1  g041(.A(G1gat), .B1(new_n233), .B2(new_n239), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n236), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n232), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n228), .A2(new_n231), .A3(new_n245), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n204), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n229), .A2(KEYINPUT92), .A3(new_n230), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT92), .B1(new_n229), .B2(new_n230), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n250), .B1(new_n229), .B2(new_n230), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n241), .A2(new_n244), .A3(KEYINPUT94), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT94), .B1(new_n241), .B2(new_n244), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n259), .A2(new_n203), .A3(new_n247), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT18), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n249), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n254), .B1(new_n232), .B2(new_n250), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n263), .A2(new_n258), .B1(new_n232), .B2(new_n246), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n264), .A2(KEYINPUT96), .A3(KEYINPUT18), .A4(new_n203), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n259), .A2(KEYINPUT18), .A3(new_n203), .A4(new_n247), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT96), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n262), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G141gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT89), .B(G197gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT11), .B(G169gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n274), .B(KEYINPUT12), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n262), .A2(new_n265), .A3(new_n268), .A4(new_n275), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G141gat), .B(G148gat), .Z(new_n281));
  INV_X1    g080(.A(G155gat), .ZN(new_n282));
  INV_X1    g081(.A(G162gat), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT2), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G155gat), .B(G162gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(KEYINPUT1), .ZN(new_n290));
  XNOR2_X1  g089(.A(G127gat), .B(G134gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n281), .A2(new_n286), .A3(new_n284), .ZN(new_n293));
  INV_X1    g092(.A(new_n291), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(KEYINPUT1), .B2(new_n289), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n288), .A2(new_n292), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(KEYINPUT4), .ZN(new_n297));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n288), .A2(new_n293), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT3), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT3), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n288), .A2(new_n301), .A3(new_n293), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n292), .A2(new_n295), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n298), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n303), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n306), .A2(new_n296), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT5), .B1(new_n307), .B2(new_n298), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G1gat), .B(G29gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT0), .ZN(new_n311));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n297), .A2(KEYINPUT5), .A3(new_n298), .A4(new_n304), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n309), .A2(KEYINPUT6), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n314), .A3(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT6), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n314), .B1(new_n309), .B2(new_n315), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G169gat), .ZN(new_n324));
  INV_X1    g123(.A(G176gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT68), .B1(new_n326), .B2(KEYINPUT26), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT69), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n332), .B2(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT69), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n329), .A4(new_n328), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n331), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  INV_X1    g139(.A(G183gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT27), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT27), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G183gat), .ZN(new_n344));
  INV_X1    g143(.A(G190gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT67), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT28), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n346), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT23), .B1(new_n332), .B2(KEYINPUT64), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT64), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354));
  OAI211_X1 g153(.A(new_n353), .B(new_n354), .C1(G169gat), .C2(G176gat), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n352), .A2(new_n355), .A3(new_n329), .ZN(new_n356));
  AND3_X1   g155(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359));
  NOR3_X1   g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT25), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n352), .A2(KEYINPUT25), .A3(new_n355), .A4(new_n329), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT66), .ZN(new_n364));
  NOR3_X1   g163(.A1(new_n364), .A2(G183gat), .A3(G190gat), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT66), .B1(new_n341), .B2(new_n345), .ZN(new_n366));
  NOR3_X1   g165(.A1(new_n365), .A2(new_n366), .A3(new_n357), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT65), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n358), .B(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n363), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n339), .A2(new_n351), .B1(new_n362), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT72), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G211gat), .A2(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(G211gat), .ZN(new_n376));
  INV_X1    g175(.A(G218gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g177(.A1(G197gat), .A2(G204gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(G197gat), .A2(G204gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT22), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n375), .B(new_n378), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n378), .A2(new_n375), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n375), .A2(new_n382), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n384), .B(new_n385), .C1(new_n380), .C2(new_n379), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n346), .A2(new_n347), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT28), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n331), .A2(new_n334), .A3(new_n338), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n340), .ZN(new_n393));
  INV_X1    g192(.A(new_n363), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n366), .A2(new_n357), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n359), .A2(KEYINPUT66), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT24), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n340), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n368), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n358), .A2(KEYINPUT65), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n395), .A2(new_n396), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT25), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n352), .A2(new_n355), .A3(new_n329), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n360), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n393), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n372), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n374), .B(new_n387), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT73), .ZN(new_n410));
  XOR2_X1   g209(.A(G8gat), .B(G36gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT75), .ZN(new_n412));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n387), .B(KEYINPUT71), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT29), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n373), .B1(new_n371), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n340), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n389), .B2(new_n390), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n419), .A2(new_n392), .B1(new_n402), .B2(new_n405), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(new_n372), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n415), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n372), .B1(new_n420), .B2(KEYINPUT29), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT73), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n387), .A4(new_n374), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n410), .A2(new_n414), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n316), .A2(KEYINPUT87), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n323), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n415), .ZN(new_n429));
  OAI221_X1 g228(.A(new_n429), .B1(new_n420), .B2(new_n372), .C1(new_n407), .C2(new_n373), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n387), .B1(new_n423), .B2(new_n374), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n373), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n393), .B2(new_n406), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n371), .A2(new_n416), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n436), .B2(new_n372), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n437), .A2(KEYINPUT83), .A3(new_n387), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT37), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n425), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n424), .B1(new_n437), .B2(new_n387), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n414), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT85), .B(KEYINPUT38), .Z(new_n447));
  OAI211_X1 g246(.A(KEYINPUT84), .B(KEYINPUT37), .C1(new_n433), .C2(new_n438), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n441), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT86), .ZN(new_n450));
  INV_X1    g249(.A(new_n447), .ZN(new_n451));
  AOI211_X1 g250(.A(new_n414), .B(new_n451), .C1(new_n444), .C2(new_n445), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n441), .A4(new_n448), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n428), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT88), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT74), .B1(new_n442), .B2(new_n443), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT74), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n410), .A2(new_n458), .A3(new_n422), .A4(new_n425), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(KEYINPUT37), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n446), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n456), .B1(new_n461), .B2(new_n451), .ZN(new_n462));
  AOI211_X1 g261(.A(KEYINPUT88), .B(new_n447), .C1(new_n460), .C2(new_n446), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n455), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT29), .B1(new_n383), .B2(new_n386), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n299), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT80), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n302), .A2(new_n416), .ZN(new_n469));
  INV_X1    g268(.A(new_n387), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n299), .B(new_n472), .C1(new_n466), .C2(KEYINPUT3), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n415), .B2(new_n469), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n466), .A2(KEYINPUT81), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n301), .B1(new_n466), .B2(KEYINPUT81), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n299), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT82), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G78gat), .B(G106gat), .Z(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT79), .B(G50gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(KEYINPUT78), .B(KEYINPUT31), .Z(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(G22gat), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n474), .A2(new_n475), .B1(new_n477), .B2(new_n480), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n490), .A2(KEYINPUT82), .ZN(new_n491));
  INV_X1    g290(.A(G22gat), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(new_n487), .C1(new_n490), .C2(KEYINPUT82), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n489), .B2(new_n493), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n497));
  NAND2_X1  g296(.A1(new_n426), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n422), .A2(new_n425), .ZN(new_n499));
  NOR2_X1   g298(.A1(KEYINPUT77), .A2(KEYINPUT30), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(new_n414), .A3(new_n410), .A4(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n414), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n457), .A2(new_n503), .A3(new_n459), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT76), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n457), .A2(new_n506), .A3(new_n503), .A4(new_n459), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n297), .A2(new_n304), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(G225gat), .A3(G233gat), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n510), .A2(KEYINPUT39), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n307), .A2(new_n298), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(KEYINPUT39), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(new_n313), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT40), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n511), .A2(KEYINPUT40), .A3(new_n313), .A4(new_n513), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n317), .A3(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n496), .B1(new_n508), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n465), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522));
  XOR2_X1   g321(.A(G15gat), .B(G43gat), .Z(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n371), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n420), .A2(KEYINPUT70), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n529), .A3(new_n303), .ZN(new_n530));
  INV_X1    g329(.A(G227gat), .ZN(new_n531));
  INV_X1    g330(.A(G233gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n371), .A2(new_n527), .A3(new_n292), .A4(new_n295), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT33), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT34), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n530), .A2(new_n534), .ZN(new_n539));
  INV_X1    g338(.A(new_n533), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI211_X1 g340(.A(KEYINPUT34), .B(new_n533), .C1(new_n530), .C2(new_n534), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n537), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n537), .A2(new_n541), .A3(new_n542), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n535), .A2(KEYINPUT32), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n546), .ZN(new_n548));
  INV_X1    g347(.A(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n539), .A2(new_n540), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT34), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n549), .B(new_n551), .C1(new_n552), .C2(new_n526), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n548), .B1(new_n553), .B2(new_n543), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n522), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n546), .B1(new_n544), .B2(new_n545), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n548), .A3(new_n543), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(KEYINPUT36), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n505), .A2(new_n507), .ZN(new_n560));
  INV_X1    g359(.A(new_n502), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n321), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n496), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n521), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n556), .A2(new_n496), .A3(new_n557), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT35), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n547), .A2(new_n554), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT35), .B1(new_n323), .B2(new_n427), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n496), .A3(new_n508), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n280), .B1(new_n566), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574));
  XOR2_X1   g373(.A(G57gat), .B(G64gat), .Z(new_n575));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g376(.A(G71gat), .ZN(new_n578));
  INV_X1    g377(.A(G78gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  XOR2_X1   g380(.A(G71gat), .B(G78gat), .Z(new_n582));
  AND2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n581), .A2(new_n582), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n574), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n581), .A2(new_n582), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(new_n582), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT98), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n246), .B1(new_n589), .B2(KEYINPUT21), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT99), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n282), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT99), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n590), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n593), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G183gat), .B(G211gat), .Z(new_n600));
  NAND2_X1  g399(.A1(new_n586), .A2(new_n587), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT21), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G127gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n605), .A2(new_n606), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n600), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  INV_X1    g410(.A(new_n600), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n595), .A2(new_n598), .A3(new_n610), .A4(new_n613), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n617), .B1(new_n618), .B2(KEYINPUT101), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(KEYINPUT7), .C1(new_n617), .C2(new_n618), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT7), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n617), .B(new_n621), .C1(new_n618), .C2(KEYINPUT101), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  INV_X1    g422(.A(G85gat), .ZN(new_n624));
  INV_X1    g423(.A(G92gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(KEYINPUT8), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G99gat), .B(G106gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n620), .A2(new_n628), .A3(new_n622), .A4(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n263), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n232), .A2(new_n634), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n640));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n638), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n633), .A2(new_n643), .A3(new_n636), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n644), .ZN(new_n646));
  INV_X1    g445(.A(new_n642), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n615), .A2(new_n616), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AND4_X1   g449(.A1(KEYINPUT10), .A2(new_n634), .A3(new_n588), .A4(new_n585), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT102), .B(KEYINPUT10), .Z(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n601), .A2(new_n631), .A3(new_n630), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n583), .A2(new_n584), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n632), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n653), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G230gat), .ZN(new_n658));
  OAI22_X1  g457(.A1(new_n651), .A2(new_n657), .B1(new_n658), .B2(new_n532), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n532), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n659), .A2(new_n661), .A3(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n650), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n573), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n321), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT103), .B(G1gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1324gat));
  INV_X1    g474(.A(new_n508), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT105), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(G8gat), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT16), .B(G8gat), .ZN(new_n681));
  OR3_X1    g480(.A1(new_n677), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n678), .A2(new_n681), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n684));
  OAI211_X1 g483(.A(new_n679), .B(new_n682), .C1(new_n683), .C2(new_n684), .ZN(G1325gat));
  INV_X1    g484(.A(new_n671), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n559), .B(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G15gat), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n569), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n690), .A2(G15gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n689), .B1(new_n686), .B2(new_n691), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n671), .A2(new_n563), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT107), .B(KEYINPUT108), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1327gat));
  AOI21_X1  g496(.A(new_n519), .B1(new_n455), .B2(new_n464), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n559), .A2(new_n564), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n572), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n648), .A2(new_n645), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n615), .A2(new_n616), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n669), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n279), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n707), .A2(new_n206), .A3(new_n672), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT45), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n703), .A2(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT109), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n703), .A2(new_n712), .A3(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n566), .A2(KEYINPUT110), .A3(new_n572), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n715), .A2(new_n717), .A3(new_n718), .A4(new_n702), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n706), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(new_n672), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n709), .B1(new_n721), .B2(new_n206), .ZN(G1328gat));
  NOR2_X1   g521(.A1(new_n701), .A2(new_n212), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n573), .A2(new_n676), .A3(new_n705), .A4(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(KEYINPUT111), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(KEYINPUT111), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n720), .A2(new_n676), .ZN(new_n729));
  OAI221_X1 g528(.A(new_n728), .B1(new_n726), .B2(new_n724), .C1(new_n729), .C2(new_n225), .ZN(G1329gat));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n712), .B1(new_n703), .B2(KEYINPUT44), .ZN(new_n732));
  AOI211_X1 g531(.A(KEYINPUT109), .B(new_n718), .C1(new_n700), .C2(new_n702), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n719), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n559), .ZN(new_n735));
  INV_X1    g534(.A(new_n706), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G43gat), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n690), .A2(G43gat), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n700), .A2(new_n702), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT112), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n731), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n731), .ZN(new_n744));
  INV_X1    g543(.A(new_n688), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n734), .A2(new_n745), .A3(new_n736), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n744), .B1(new_n746), .B2(G43gat), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT113), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(G43gat), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n741), .B1(new_n737), .B2(G43gat), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n751), .B(new_n752), .C1(new_n731), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n748), .A2(new_n754), .ZN(G1330gat));
  INV_X1    g554(.A(G50gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n720), .B2(new_n563), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n707), .A2(new_n756), .A3(new_n563), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT48), .B1(new_n758), .B2(KEYINPUT114), .ZN(new_n760));
  OR3_X1    g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n760), .B1(new_n757), .B2(new_n759), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1331gat));
  AND2_X1   g562(.A1(new_n715), .A2(new_n717), .ZN(new_n764));
  INV_X1    g563(.A(new_n669), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n279), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n650), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n672), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n508), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(G1333gat));
  OAI21_X1  g576(.A(G71gat), .B1(new_n769), .B2(new_n688), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n569), .A2(new_n578), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n769), .B2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1334gat));
  NOR2_X1   g581(.A1(new_n769), .A2(new_n496), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(new_n579), .ZN(G1335gat));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n704), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n734), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT116), .B1(new_n786), .B2(new_n321), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G85gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n786), .A2(KEYINPUT116), .A3(new_n321), .ZN(new_n789));
  INV_X1    g588(.A(new_n704), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n700), .A2(new_n280), .A3(new_n790), .A4(new_n702), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n669), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n672), .A2(new_n624), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n788), .A2(new_n789), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  OAI21_X1  g596(.A(G92gat), .B1(new_n786), .B2(new_n508), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n676), .A2(new_n625), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT52), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n798), .B(new_n802), .C1(new_n795), .C2(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1337gat));
  OAI21_X1  g603(.A(G99gat), .B1(new_n786), .B2(new_n688), .ZN(new_n805));
  OR2_X1    g604(.A1(new_n690), .A2(G99gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n795), .B2(new_n806), .ZN(G1338gat));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(KEYINPUT53), .ZN(new_n810));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  INV_X1    g610(.A(new_n785), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n714), .B2(new_n719), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n563), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n496), .A2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n795), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n809), .B(new_n810), .C1(new_n814), .C2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n786), .B2(new_n496), .ZN(new_n819));
  INV_X1    g618(.A(new_n817), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n820), .A3(new_n808), .A4(KEYINPUT53), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n818), .A2(new_n821), .ZN(G1339gat));
  NOR3_X1   g621(.A1(new_n650), .A2(new_n279), .A3(new_n669), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n264), .A2(new_n203), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n247), .A2(new_n248), .A3(new_n204), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n274), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n278), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n654), .A2(new_n656), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n652), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n589), .A2(KEYINPUT10), .A3(new_n634), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n660), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n665), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n829), .A2(new_n830), .A3(new_n660), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n659), .A2(new_n834), .A3(KEYINPUT54), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI221_X1 g637(.A(new_n832), .B1(new_n658), .B2(new_n532), .C1(new_n651), .C2(new_n657), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n835), .A2(KEYINPUT55), .A3(new_n666), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n668), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n702), .A2(new_n827), .A3(new_n838), .A4(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n278), .A2(new_n669), .A3(new_n826), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n841), .B1(new_n277), .B2(new_n278), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n838), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n843), .B1(new_n846), .B2(new_n702), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n823), .B1(new_n847), .B2(new_n790), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n321), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n496), .A3(new_n569), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT119), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n676), .B1(new_n850), .B2(KEYINPUT119), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853), .B2(new_n279), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n676), .A2(new_n321), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT118), .B1(new_n848), .B2(new_n563), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT55), .B1(new_n833), .B2(new_n835), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n859), .B(new_n841), .C1(new_n277), .C2(new_n278), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n701), .B1(new_n860), .B2(new_n844), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n704), .B1(new_n861), .B2(new_n843), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n858), .B(new_n496), .C1(new_n862), .C2(new_n823), .ZN(new_n863));
  AOI211_X1 g662(.A(new_n690), .B(new_n856), .C1(new_n857), .C2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n279), .A2(G113gat), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n854), .B1(new_n864), .B2(new_n865), .ZN(G1340gat));
  AOI21_X1  g665(.A(G120gat), .B1(new_n853), .B2(new_n669), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n669), .A2(G120gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(new_n864), .B2(new_n868), .ZN(G1341gat));
  AND4_X1   g668(.A1(new_n606), .A2(new_n851), .A3(new_n704), .A4(new_n852), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n606), .B1(new_n864), .B2(new_n704), .ZN(new_n871));
  OR3_X1    g670(.A1(new_n870), .A2(KEYINPUT120), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(KEYINPUT120), .B1(new_n870), .B2(new_n871), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1342gat));
  AND2_X1   g673(.A1(new_n864), .A2(new_n702), .ZN(new_n875));
  INV_X1    g674(.A(G134gat), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n853), .A2(new_n876), .A3(new_n702), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n879), .B1(KEYINPUT56), .B2(new_n878), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n745), .A2(new_n496), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT122), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n676), .B1(new_n881), .B2(KEYINPUT122), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(new_n849), .A3(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(G141gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n279), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n838), .B(KEYINPUT121), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n844), .B1(new_n887), .B2(new_n845), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n843), .B1(new_n888), .B2(new_n702), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n823), .B1(new_n889), .B2(new_n790), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT57), .B1(new_n890), .B2(new_n496), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n279), .A2(new_n838), .A3(new_n842), .ZN(new_n892));
  INV_X1    g691(.A(new_n844), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n702), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n843), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n790), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n823), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n899), .A3(new_n563), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n856), .A2(new_n735), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n891), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G141gat), .B1(new_n902), .B2(new_n280), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g704(.A(G148gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n906), .A3(new_n669), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n902), .A2(new_n765), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(KEYINPUT59), .A3(new_n906), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n899), .B1(new_n890), .B2(new_n496), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n848), .A2(new_n899), .A3(new_n496), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n669), .B(new_n901), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n910), .B1(new_n914), .B2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n907), .B1(new_n909), .B2(new_n915), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n884), .A2(new_n282), .A3(new_n704), .ZN(new_n917));
  OAI21_X1  g716(.A(G155gat), .B1(new_n902), .B2(new_n790), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n283), .A3(new_n701), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n884), .A2(new_n702), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n283), .ZN(G1347gat));
  NOR2_X1   g721(.A1(new_n848), .A2(new_n672), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n567), .A2(new_n508), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(G169gat), .B1(new_n926), .B2(new_n279), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n857), .A2(new_n863), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n508), .A2(new_n672), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n569), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n928), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g735(.A(KEYINPUT124), .B(new_n934), .C1(new_n857), .C2(new_n863), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n280), .A2(new_n324), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n927), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  NAND3_X1  g739(.A1(new_n926), .A2(new_n325), .A3(new_n669), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n936), .A2(new_n937), .A3(new_n765), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n325), .ZN(G1349gat));
  AND4_X1   g742(.A1(new_n342), .A2(new_n926), .A3(new_n344), .A4(new_n704), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n936), .A2(new_n937), .A3(new_n790), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n341), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT60), .ZN(new_n949));
  XOR2_X1   g748(.A(new_n947), .B(new_n949), .Z(G1350gat));
  NAND3_X1  g749(.A1(new_n926), .A2(new_n345), .A3(new_n702), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n858), .B1(new_n898), .B2(new_n496), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT118), .B(new_n563), .C1(new_n896), .C2(new_n897), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n935), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT124), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n929), .A2(new_n928), .A3(new_n935), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n702), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT126), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n957), .A2(new_n958), .A3(G190gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n957), .B2(G190gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(KEYINPUT61), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n936), .A2(new_n937), .A3(new_n701), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT126), .B1(new_n963), .B2(new_n345), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n957), .A2(new_n958), .A3(G190gat), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n951), .B1(new_n961), .B2(new_n966), .ZN(G1351gat));
  OAI211_X1 g766(.A(new_n688), .B(new_n930), .C1(new_n912), .C2(new_n913), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(G197gat), .A3(new_n279), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n881), .A2(new_n676), .A3(new_n923), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n279), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n970), .A2(new_n972), .ZN(G1352gat));
  AOI21_X1  g772(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n971), .A2(new_n669), .A3(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G204gat), .B1(new_n968), .B2(new_n765), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1353gat));
  NAND3_X1  g778(.A1(new_n971), .A2(new_n376), .A3(new_n704), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n376), .B1(new_n969), .B2(new_n704), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n981), .A2(KEYINPUT63), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(KEYINPUT63), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n968), .B2(new_n701), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n971), .A2(new_n377), .A3(new_n702), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


