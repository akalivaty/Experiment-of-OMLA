

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X2 U550 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n727) );
  XOR2_X2 U551 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X2 U552 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n786) );
  NOR2_X1 U553 ( .A1(n529), .A2(n527), .ZN(n523) );
  NOR2_X2 U554 ( .A1(G651), .A2(G543), .ZN(n649) );
  AND2_X1 U555 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X2 U556 ( .A1(n578), .A2(n577), .ZN(n988) );
  NOR2_X2 U557 ( .A1(n576), .A2(n575), .ZN(n578) );
  INV_X2 U558 ( .A(n724), .ZN(n726) );
  AND2_X2 U559 ( .A1(n726), .A2(n725), .ZN(n516) );
  NOR2_X4 U560 ( .A1(n543), .A2(G2105), .ZN(n891) );
  NOR2_X1 U561 ( .A1(n827), .A2(n826), .ZN(n829) );
  NOR2_X1 U562 ( .A1(n823), .A2(n822), .ZN(n825) );
  NOR2_X1 U563 ( .A1(n738), .A2(n1002), .ZN(n733) );
  INV_X2 U564 ( .A(G2104), .ZN(n543) );
  XNOR2_X1 U565 ( .A(n825), .B(n824), .ZN(n826) );
  OR2_X1 U566 ( .A1(n545), .A2(n544), .ZN(n707) );
  AND2_X1 U567 ( .A1(n561), .A2(n560), .ZN(n563) );
  AND2_X1 U568 ( .A1(n706), .A2(G137), .ZN(n519) );
  BUF_X1 U569 ( .A(n706), .Z(n539) );
  XNOR2_X1 U570 ( .A(n559), .B(n558), .ZN(n561) );
  BUF_X1 U571 ( .A(n517), .Z(n609) );
  XNOR2_X1 U572 ( .A(n538), .B(n537), .ZN(n706) );
  XNOR2_X1 U573 ( .A(n536), .B(KEYINPUT66), .ZN(n538) );
  XNOR2_X1 U574 ( .A(n540), .B(KEYINPUT65), .ZN(n517) );
  BUF_X1 U575 ( .A(n789), .Z(n518) );
  XNOR2_X1 U576 ( .A(n540), .B(KEYINPUT65), .ZN(n608) );
  XNOR2_X1 U577 ( .A(G543), .B(KEYINPUT0), .ZN(n522) );
  INV_X1 U578 ( .A(KEYINPUT96), .ZN(n750) );
  XNOR2_X1 U579 ( .A(n523), .B(KEYINPUT68), .ZN(n581) );
  NAND2_X1 U580 ( .A1(n557), .A2(G2104), .ZN(n559) );
  NOR2_X1 U581 ( .A1(n556), .A2(G2105), .ZN(n557) );
  XOR2_X1 U582 ( .A(KEYINPUT89), .B(n821), .Z(n822) );
  NOR2_X1 U583 ( .A1(G543), .A2(n527), .ZN(n528) );
  INV_X1 U584 ( .A(KEYINPUT17), .ZN(n536) );
  AND2_X1 U585 ( .A1(G66), .A2(n648), .ZN(n520) );
  INV_X1 U586 ( .A(KEYINPUT94), .ZN(n732) );
  XNOR2_X1 U587 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n768) );
  XNOR2_X1 U588 ( .A(n769), .B(n768), .ZN(n770) );
  BUF_X1 U589 ( .A(n764), .Z(n778) );
  INV_X1 U590 ( .A(G101), .ZN(n556) );
  INV_X1 U591 ( .A(KEYINPUT23), .ZN(n558) );
  INV_X1 U592 ( .A(KEYINPUT103), .ZN(n824) );
  AND2_X1 U593 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U594 ( .A(KEYINPUT13), .ZN(n573) );
  INV_X1 U595 ( .A(KEYINPUT104), .ZN(n828) );
  BUF_X1 U596 ( .A(n529), .Z(n628) );
  BUF_X1 U597 ( .A(n581), .Z(n653) );
  NAND2_X1 U598 ( .A1(n649), .A2(G89), .ZN(n521) );
  XNOR2_X1 U599 ( .A(n521), .B(KEYINPUT4), .ZN(n525) );
  INV_X1 U600 ( .A(n522), .ZN(n529) );
  INV_X1 U601 ( .A(G651), .ZN(n527) );
  NAND2_X1 U602 ( .A1(G76), .A2(n653), .ZN(n524) );
  NAND2_X1 U603 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U604 ( .A(n526), .B(KEYINPUT5), .ZN(n534) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n528), .Z(n568) );
  BUF_X2 U606 ( .A(n568), .Z(n648) );
  NAND2_X1 U607 ( .A1(G63), .A2(n648), .ZN(n531) );
  NOR2_X4 U608 ( .A1(n628), .A2(G651), .ZN(n650) );
  NAND2_X1 U609 ( .A1(G51), .A2(n650), .ZN(n530) );
  NAND2_X1 U610 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U611 ( .A(KEYINPUT6), .B(n532), .Z(n533) );
  NAND2_X1 U612 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U613 ( .A(n535), .B(KEYINPUT7), .ZN(G168) );
  NOR2_X1 U614 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  NAND2_X1 U615 ( .A1(G138), .A2(n539), .ZN(n547) );
  NAND2_X1 U616 ( .A1(G114), .A2(n888), .ZN(n542) );
  NAND2_X1 U617 ( .A1(n543), .A2(G2105), .ZN(n540) );
  NAND2_X1 U618 ( .A1(n608), .A2(G126), .ZN(n541) );
  NAND2_X1 U619 ( .A1(n542), .A2(n541), .ZN(n545) );
  AND2_X1 U620 ( .A1(G102), .A2(n891), .ZN(n544) );
  INV_X1 U621 ( .A(n707), .ZN(n546) );
  AND2_X1 U622 ( .A1(n547), .A2(n546), .ZN(G164) );
  NAND2_X1 U623 ( .A1(G64), .A2(n648), .ZN(n549) );
  NAND2_X1 U624 ( .A1(G52), .A2(n650), .ZN(n548) );
  NAND2_X1 U625 ( .A1(n549), .A2(n548), .ZN(n555) );
  NAND2_X1 U626 ( .A1(G77), .A2(n653), .ZN(n550) );
  XNOR2_X1 U627 ( .A(n550), .B(KEYINPUT70), .ZN(n552) );
  NAND2_X1 U628 ( .A1(G90), .A2(n649), .ZN(n551) );
  NAND2_X1 U629 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U630 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U631 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U632 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U633 ( .A(G57), .ZN(G237) );
  NAND2_X1 U634 ( .A1(n888), .A2(G113), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n517), .A2(G125), .ZN(n562) );
  NAND2_X1 U636 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X2 U637 ( .A1(n564), .A2(n519), .ZN(n710) );
  BUF_X1 U638 ( .A(n710), .Z(G160) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U640 ( .A(n566), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n846) );
  NAND2_X1 U642 ( .A1(n846), .A2(G567), .ZN(n567) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  NAND2_X1 U644 ( .A1(G56), .A2(n568), .ZN(n569) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n569), .Z(n576) );
  NAND2_X1 U646 ( .A1(n649), .A2(G81), .ZN(n570) );
  XNOR2_X1 U647 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n581), .A2(G68), .ZN(n571) );
  NAND2_X1 U649 ( .A1(n572), .A2(n571), .ZN(n574) );
  XNOR2_X1 U650 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n650), .A2(G43), .ZN(n577) );
  INV_X1 U652 ( .A(G860), .ZN(n600) );
  OR2_X1 U653 ( .A1(n988), .A2(n600), .ZN(G153) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(n649), .A2(G92), .ZN(n579) );
  XOR2_X1 U656 ( .A(KEYINPUT72), .B(n579), .Z(n580) );
  NOR2_X1 U657 ( .A1(n520), .A2(n580), .ZN(n586) );
  NAND2_X1 U658 ( .A1(G79), .A2(n581), .ZN(n583) );
  NAND2_X1 U659 ( .A1(n650), .A2(G54), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U661 ( .A(n584), .B(KEYINPUT73), .ZN(n585) );
  XNOR2_X2 U662 ( .A(KEYINPUT15), .B(n587), .ZN(n1002) );
  NOR2_X1 U663 ( .A1(G868), .A2(n1002), .ZN(n589) );
  INV_X1 U664 ( .A(G868), .ZN(n670) );
  NOR2_X1 U665 ( .A1(n670), .A2(G301), .ZN(n588) );
  NOR2_X1 U666 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U667 ( .A(KEYINPUT74), .B(n590), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n649), .A2(G91), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G78), .A2(n653), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G65), .A2(n648), .ZN(n593) );
  XNOR2_X1 U672 ( .A(KEYINPUT71), .B(n593), .ZN(n594) );
  NOR2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U674 ( .A1(n650), .A2(G53), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U676 ( .A1(G286), .A2(n670), .ZN(n599) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U678 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n600), .A2(G559), .ZN(n601) );
  INV_X1 U680 ( .A(n1002), .ZN(n913) );
  NAND2_X1 U681 ( .A1(n601), .A2(n913), .ZN(n602) );
  XNOR2_X1 U682 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n988), .ZN(n605) );
  NAND2_X1 U684 ( .A1(G868), .A2(n913), .ZN(n603) );
  NOR2_X1 U685 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U686 ( .A1(n605), .A2(n604), .ZN(G282) );
  XNOR2_X1 U687 ( .A(G2100), .B(KEYINPUT75), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G99), .A2(n891), .ZN(n607) );
  NAND2_X1 U689 ( .A1(G111), .A2(n888), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G123), .A2(n609), .ZN(n610) );
  XNOR2_X1 U692 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G135), .A2(n539), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n938) );
  XNOR2_X1 U696 ( .A(n938), .B(G2096), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U698 ( .A1(n913), .A2(G559), .ZN(n667) );
  XNOR2_X1 U699 ( .A(n988), .B(n667), .ZN(n617) );
  NOR2_X1 U700 ( .A1(n617), .A2(G860), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n649), .A2(G93), .ZN(n619) );
  NAND2_X1 U702 ( .A1(G80), .A2(n653), .ZN(n618) );
  NAND2_X1 U703 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U704 ( .A(KEYINPUT76), .B(n620), .Z(n622) );
  NAND2_X1 U705 ( .A1(n648), .A2(G67), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U707 ( .A1(G55), .A2(n650), .ZN(n623) );
  XNOR2_X1 U708 ( .A(KEYINPUT77), .B(n623), .ZN(n624) );
  OR2_X1 U709 ( .A1(n625), .A2(n624), .ZN(n669) );
  XOR2_X1 U710 ( .A(n626), .B(n669), .Z(G145) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n627) );
  XNOR2_X1 U712 ( .A(n627), .B(KEYINPUT78), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G49), .A2(n650), .ZN(n630) );
  NAND2_X1 U714 ( .A1(G87), .A2(n628), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U716 ( .A1(n648), .A2(n631), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(G288) );
  NAND2_X1 U718 ( .A1(n649), .A2(G88), .ZN(n635) );
  NAND2_X1 U719 ( .A1(G75), .A2(n653), .ZN(n634) );
  NAND2_X1 U720 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G62), .A2(n648), .ZN(n637) );
  NAND2_X1 U722 ( .A1(G50), .A2(n650), .ZN(n636) );
  NAND2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U724 ( .A1(n639), .A2(n638), .ZN(G166) );
  NAND2_X1 U725 ( .A1(G60), .A2(n648), .ZN(n641) );
  NAND2_X1 U726 ( .A1(G47), .A2(n650), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U728 ( .A1(G72), .A2(n653), .ZN(n642) );
  XNOR2_X1 U729 ( .A(KEYINPUT69), .B(n642), .ZN(n643) );
  NOR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n649), .A2(G85), .ZN(n645) );
  XOR2_X1 U732 ( .A(KEYINPUT67), .B(n645), .Z(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(G290) );
  NAND2_X1 U734 ( .A1(n648), .A2(G61), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G86), .A2(n649), .ZN(n652) );
  NAND2_X1 U736 ( .A1(G48), .A2(n650), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U739 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U740 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U742 ( .A(KEYINPUT79), .B(n659), .Z(G305) );
  XOR2_X1 U743 ( .A(KEYINPUT80), .B(KEYINPUT19), .Z(n660) );
  XNOR2_X1 U744 ( .A(G288), .B(n660), .ZN(n663) );
  XNOR2_X1 U745 ( .A(G166), .B(G299), .ZN(n661) );
  XNOR2_X1 U746 ( .A(n661), .B(n988), .ZN(n662) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n665) );
  XOR2_X1 U748 ( .A(G290), .B(n669), .Z(n664) );
  XNOR2_X1 U749 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n666), .B(G305), .ZN(n912) );
  XNOR2_X1 U751 ( .A(n667), .B(n912), .ZN(n668) );
  NAND2_X1 U752 ( .A1(n668), .A2(G868), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U755 ( .A(KEYINPUT81), .B(n673), .Z(G295) );
  NAND2_X1 U756 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(KEYINPUT82), .Z(n679) );
  NAND2_X1 U763 ( .A1(G132), .A2(G82), .ZN(n678) );
  XNOR2_X1 U764 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n680), .A2(G96), .ZN(n681) );
  NOR2_X1 U766 ( .A1(n681), .A2(G218), .ZN(n682) );
  XNOR2_X1 U767 ( .A(n682), .B(KEYINPUT83), .ZN(n850) );
  NAND2_X1 U768 ( .A1(n850), .A2(G2106), .ZN(n686) );
  NAND2_X1 U769 ( .A1(G120), .A2(G69), .ZN(n683) );
  NOR2_X1 U770 ( .A1(G237), .A2(n683), .ZN(n684) );
  NAND2_X1 U771 ( .A1(G108), .A2(n684), .ZN(n851) );
  NAND2_X1 U772 ( .A1(n851), .A2(G567), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n852) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n687) );
  NOR2_X1 U775 ( .A1(n852), .A2(n687), .ZN(n849) );
  NAND2_X1 U776 ( .A1(n849), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  XOR2_X1 U778 ( .A(G1986), .B(G290), .Z(n992) );
  NAND2_X1 U779 ( .A1(G95), .A2(n891), .ZN(n689) );
  NAND2_X1 U780 ( .A1(G107), .A2(n888), .ZN(n688) );
  NAND2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n609), .A2(G119), .ZN(n691) );
  NAND2_X1 U783 ( .A1(G131), .A2(n539), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n901) );
  NAND2_X1 U786 ( .A1(G1991), .A2(n901), .ZN(n694) );
  XOR2_X1 U787 ( .A(KEYINPUT86), .B(n694), .Z(n703) );
  NAND2_X1 U788 ( .A1(n891), .A2(G105), .ZN(n695) );
  XNOR2_X1 U789 ( .A(n695), .B(KEYINPUT38), .ZN(n697) );
  NAND2_X1 U790 ( .A1(G117), .A2(n888), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n609), .A2(G129), .ZN(n699) );
  NAND2_X1 U793 ( .A1(G141), .A2(n539), .ZN(n698) );
  NAND2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n902) );
  INV_X1 U796 ( .A(G1996), .ZN(n965) );
  NOR2_X1 U797 ( .A1(n902), .A2(n965), .ZN(n702) );
  NOR2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n830) );
  NAND2_X1 U799 ( .A1(n992), .A2(n830), .ZN(n711) );
  INV_X1 U800 ( .A(G1384), .ZN(n704) );
  AND2_X1 U801 ( .A1(G138), .A2(n704), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n704), .A2(n707), .ZN(n708) );
  NAND2_X1 U804 ( .A1(n709), .A2(n708), .ZN(n725) );
  NAND2_X1 U805 ( .A1(n710), .A2(G40), .ZN(n724) );
  NOR2_X1 U806 ( .A1(n725), .A2(n724), .ZN(n841) );
  NAND2_X1 U807 ( .A1(n711), .A2(n841), .ZN(n723) );
  NAND2_X1 U808 ( .A1(G104), .A2(n891), .ZN(n713) );
  NAND2_X1 U809 ( .A1(G140), .A2(n539), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U811 ( .A(KEYINPUT34), .B(n714), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n609), .A2(G128), .ZN(n715) );
  XNOR2_X1 U813 ( .A(n715), .B(KEYINPUT84), .ZN(n717) );
  NAND2_X1 U814 ( .A1(G116), .A2(n888), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U816 ( .A(n718), .B(KEYINPUT35), .Z(n719) );
  NOR2_X1 U817 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U818 ( .A(KEYINPUT36), .B(n721), .Z(n722) );
  XNOR2_X1 U819 ( .A(KEYINPUT85), .B(n722), .ZN(n909) );
  XNOR2_X1 U820 ( .A(KEYINPUT37), .B(G2067), .ZN(n838) );
  NOR2_X1 U821 ( .A1(n909), .A2(n838), .ZN(n945) );
  NAND2_X1 U822 ( .A1(n841), .A2(n945), .ZN(n836) );
  NAND2_X1 U823 ( .A1(n723), .A2(n836), .ZN(n827) );
  NAND2_X1 U824 ( .A1(n726), .A2(n725), .ZN(n764) );
  NAND2_X1 U825 ( .A1(n516), .A2(G1996), .ZN(n728) );
  XNOR2_X1 U826 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U827 ( .A1(n729), .A2(n988), .ZN(n731) );
  NAND2_X1 U828 ( .A1(G1341), .A2(n778), .ZN(n730) );
  NAND2_X1 U829 ( .A1(n731), .A2(n730), .ZN(n738) );
  XNOR2_X1 U830 ( .A(n733), .B(n732), .ZN(n737) );
  NAND2_X1 U831 ( .A1(G1348), .A2(n778), .ZN(n735) );
  INV_X1 U832 ( .A(n764), .ZN(n759) );
  XOR2_X1 U833 ( .A(n759), .B(KEYINPUT90), .Z(n758) );
  INV_X1 U834 ( .A(n758), .ZN(n742) );
  NAND2_X1 U835 ( .A1(G2067), .A2(n742), .ZN(n734) );
  NAND2_X1 U836 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U837 ( .A1(n737), .A2(n736), .ZN(n740) );
  NAND2_X1 U838 ( .A1(n738), .A2(n1002), .ZN(n739) );
  NAND2_X1 U839 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U840 ( .A(n741), .B(KEYINPUT95), .ZN(n749) );
  XOR2_X1 U841 ( .A(KEYINPUT27), .B(KEYINPUT92), .Z(n744) );
  NAND2_X1 U842 ( .A1(G2072), .A2(n742), .ZN(n743) );
  XNOR2_X1 U843 ( .A(n744), .B(n743), .ZN(n747) );
  NAND2_X1 U844 ( .A1(n758), .A2(G1956), .ZN(n745) );
  XOR2_X1 U845 ( .A(KEYINPUT93), .B(n745), .Z(n746) );
  NAND2_X1 U846 ( .A1(n747), .A2(n746), .ZN(n752) );
  NOR2_X1 U847 ( .A1(G299), .A2(n752), .ZN(n748) );
  NOR2_X1 U848 ( .A1(n749), .A2(n748), .ZN(n751) );
  XNOR2_X1 U849 ( .A(n751), .B(n750), .ZN(n755) );
  NAND2_X1 U850 ( .A1(G299), .A2(n752), .ZN(n753) );
  XNOR2_X1 U851 ( .A(KEYINPUT28), .B(n753), .ZN(n754) );
  NAND2_X1 U852 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U853 ( .A(n756), .B(KEYINPUT29), .ZN(n763) );
  XNOR2_X1 U854 ( .A(G2078), .B(KEYINPUT91), .ZN(n757) );
  XNOR2_X1 U855 ( .A(n757), .B(KEYINPUT25), .ZN(n963) );
  NOR2_X1 U856 ( .A1(n963), .A2(n758), .ZN(n761) );
  NOR2_X1 U857 ( .A1(n759), .A2(G1961), .ZN(n760) );
  NOR2_X1 U858 ( .A1(n761), .A2(n760), .ZN(n771) );
  NOR2_X1 U859 ( .A1(G301), .A2(n771), .ZN(n762) );
  NOR2_X1 U860 ( .A1(n763), .A2(n762), .ZN(n776) );
  AND2_X1 U861 ( .A1(n764), .A2(G8), .ZN(n765) );
  XNOR2_X2 U862 ( .A(KEYINPUT87), .B(n765), .ZN(n820) );
  NOR2_X1 U863 ( .A1(G1966), .A2(n820), .ZN(n791) );
  NOR2_X1 U864 ( .A1(G2084), .A2(n778), .ZN(n788) );
  NOR2_X1 U865 ( .A1(n791), .A2(n788), .ZN(n766) );
  XOR2_X1 U866 ( .A(KEYINPUT97), .B(n766), .Z(n767) );
  NAND2_X1 U867 ( .A1(n767), .A2(G8), .ZN(n769) );
  NOR2_X1 U868 ( .A1(G168), .A2(n770), .ZN(n773) );
  AND2_X1 U869 ( .A1(G301), .A2(n771), .ZN(n772) );
  NOR2_X1 U870 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U871 ( .A(n774), .B(KEYINPUT31), .ZN(n775) );
  NOR2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U873 ( .A(n777), .B(KEYINPUT99), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n789), .A2(G286), .ZN(n783) );
  NOR2_X1 U875 ( .A1(G1971), .A2(n820), .ZN(n780) );
  NOR2_X1 U876 ( .A1(G2090), .A2(n778), .ZN(n779) );
  NOR2_X1 U877 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U878 ( .A1(n781), .A2(G303), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U880 ( .A(n784), .B(KEYINPUT100), .ZN(n785) );
  NAND2_X1 U881 ( .A1(n785), .A2(G8), .ZN(n787) );
  XNOR2_X1 U882 ( .A(n787), .B(n786), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G8), .A2(n788), .ZN(n793) );
  INV_X1 U884 ( .A(n518), .ZN(n790) );
  NOR2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U886 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n813) );
  NOR2_X1 U888 ( .A1(G1976), .A2(G288), .ZN(n797) );
  NOR2_X1 U889 ( .A1(G1971), .A2(G303), .ZN(n796) );
  NOR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n994) );
  NAND2_X1 U891 ( .A1(n797), .A2(KEYINPUT33), .ZN(n798) );
  NOR2_X1 U892 ( .A1(n798), .A2(n820), .ZN(n801) );
  XOR2_X1 U893 ( .A(KEYINPUT102), .B(G1981), .Z(n799) );
  XNOR2_X1 U894 ( .A(G305), .B(n799), .ZN(n985) );
  INV_X1 U895 ( .A(n985), .ZN(n800) );
  NOR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n805), .A2(KEYINPUT33), .ZN(n803) );
  AND2_X1 U898 ( .A1(n994), .A2(n803), .ZN(n802) );
  NAND2_X1 U899 ( .A1(n813), .A2(n802), .ZN(n810) );
  INV_X1 U900 ( .A(n803), .ZN(n808) );
  INV_X1 U901 ( .A(n820), .ZN(n804) );
  NAND2_X1 U902 ( .A1(G1976), .A2(G288), .ZN(n993) );
  AND2_X1 U903 ( .A1(n804), .A2(n993), .ZN(n806) );
  AND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n816) );
  NOR2_X1 U907 ( .A1(G2090), .A2(G303), .ZN(n811) );
  NAND2_X1 U908 ( .A1(G8), .A2(n811), .ZN(n812) );
  NAND2_X1 U909 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n820), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n823) );
  NOR2_X1 U912 ( .A1(G1981), .A2(G305), .ZN(n817) );
  XOR2_X1 U913 ( .A(n817), .B(KEYINPUT88), .Z(n818) );
  XNOR2_X1 U914 ( .A(KEYINPUT24), .B(n818), .ZN(n819) );
  NOR2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U916 ( .A(n829), .B(n828), .ZN(n844) );
  AND2_X1 U917 ( .A1(n965), .A2(n902), .ZN(n936) );
  INV_X1 U918 ( .A(n830), .ZN(n941) );
  NOR2_X1 U919 ( .A1(G1991), .A2(n901), .ZN(n939) );
  NOR2_X1 U920 ( .A1(G1986), .A2(G290), .ZN(n831) );
  NOR2_X1 U921 ( .A1(n939), .A2(n831), .ZN(n832) );
  XOR2_X1 U922 ( .A(KEYINPUT105), .B(n832), .Z(n833) );
  NOR2_X1 U923 ( .A1(n941), .A2(n833), .ZN(n834) );
  NOR2_X1 U924 ( .A1(n936), .A2(n834), .ZN(n835) );
  XNOR2_X1 U925 ( .A(n835), .B(KEYINPUT39), .ZN(n837) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(n839) );
  NAND2_X1 U927 ( .A1(n909), .A2(n838), .ZN(n948) );
  NAND2_X1 U928 ( .A1(n839), .A2(n948), .ZN(n840) );
  XNOR2_X1 U929 ( .A(KEYINPUT106), .B(n840), .ZN(n842) );
  NAND2_X1 U930 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U931 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U932 ( .A(n845), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n846), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U935 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U937 ( .A1(n849), .A2(n848), .ZN(G188) );
  XOR2_X1 U938 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U940 ( .A(G132), .ZN(G219) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G82), .ZN(G220) );
  NOR2_X1 U944 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  INV_X1 U946 ( .A(n852), .ZN(G319) );
  XNOR2_X1 U947 ( .A(G1961), .B(KEYINPUT41), .ZN(n862) );
  XOR2_X1 U948 ( .A(G1956), .B(G1971), .Z(n854) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1976), .ZN(n853) );
  XNOR2_X1 U950 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U951 ( .A(G1966), .B(G1981), .Z(n856) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U954 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U955 ( .A(KEYINPUT110), .B(G2474), .ZN(n859) );
  XNOR2_X1 U956 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n862), .B(n861), .ZN(G229) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2090), .Z(n864) );
  XNOR2_X1 U959 ( .A(G2078), .B(G2084), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U961 ( .A(n865), .B(G2096), .Z(n867) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U964 ( .A(G2100), .B(KEYINPUT43), .Z(n869) );
  XNOR2_X1 U965 ( .A(G2678), .B(KEYINPUT109), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U967 ( .A(n871), .B(n870), .Z(G227) );
  NAND2_X1 U968 ( .A1(G100), .A2(n891), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G112), .A2(n888), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n879) );
  NAND2_X1 U971 ( .A1(G124), .A2(n609), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT44), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n539), .A2(G136), .ZN(n875) );
  XOR2_X1 U974 ( .A(KEYINPUT111), .B(n875), .Z(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U976 ( .A1(n879), .A2(n878), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G103), .A2(n891), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G139), .A2(n539), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U980 ( .A(KEYINPUT112), .B(n882), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G115), .A2(n888), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G127), .A2(n609), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U985 ( .A1(n887), .A2(n886), .ZN(n949) );
  NAND2_X1 U986 ( .A1(G118), .A2(n888), .ZN(n890) );
  NAND2_X1 U987 ( .A1(G130), .A2(n609), .ZN(n889) );
  NAND2_X1 U988 ( .A1(n890), .A2(n889), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G106), .A2(n891), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G142), .A2(n539), .ZN(n892) );
  NAND2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n894), .Z(n895) );
  NOR2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n949), .B(n897), .ZN(n908) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n899) );
  XNOR2_X1 U996 ( .A(G162), .B(KEYINPUT113), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U998 ( .A(G164), .B(n900), .ZN(n906) );
  XNOR2_X1 U999 ( .A(n901), .B(n938), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(G160), .B(n902), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1004 ( .A(n910), .B(n909), .Z(n911) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n911), .ZN(G395) );
  XOR2_X1 U1006 ( .A(n912), .B(G286), .Z(n915) );
  XNOR2_X1 U1007 ( .A(G171), .B(n913), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n916), .ZN(G397) );
  XOR2_X1 U1010 ( .A(G2430), .B(G2451), .Z(n918) );
  XNOR2_X1 U1011 ( .A(G2446), .B(G2427), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n925) );
  XOR2_X1 U1013 ( .A(G2438), .B(G2435), .Z(n920) );
  XNOR2_X1 U1014 ( .A(G2443), .B(KEYINPUT107), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n920), .B(n919), .ZN(n921) );
  XOR2_X1 U1016 ( .A(n921), .B(G2454), .Z(n923) );
  XNOR2_X1 U1017 ( .A(G1341), .B(G1348), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1019 ( .A(n925), .B(n924), .ZN(n926) );
  NAND2_X1 U1020 ( .A1(n926), .A2(G14), .ZN(n934) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n934), .ZN(n931) );
  XNOR2_X1 U1022 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(G229), .A2(G227), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1025 ( .A(KEYINPUT49), .B(n929), .Z(n930) );
  NOR2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  INV_X1 U1030 ( .A(G108), .ZN(G238) );
  INV_X1 U1031 ( .A(n934), .ZN(G401) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n937), .Z(n957) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n943) );
  XOR2_X1 U1036 ( .A(G160), .B(G2084), .Z(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(n946), .B(KEYINPUT116), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n955) );
  XNOR2_X1 U1042 ( .A(G2072), .B(n949), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G164), .B(G2078), .ZN(n950) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1045 ( .A(KEYINPUT117), .B(n952), .Z(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT50), .B(n953), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(KEYINPUT52), .B(n958), .ZN(n959) );
  NAND2_X1 U1050 ( .A1(n959), .A2(G29), .ZN(n1040) );
  XOR2_X1 U1051 ( .A(G1991), .B(G25), .Z(n960) );
  NAND2_X1 U1052 ( .A1(n960), .A2(G28), .ZN(n973) );
  XNOR2_X1 U1053 ( .A(G2067), .B(G26), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(G33), .B(G2072), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n971) );
  XNOR2_X1 U1056 ( .A(n963), .B(KEYINPUT118), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n964), .B(G27), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(KEYINPUT119), .B(G32), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n966), .B(n965), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n969), .B(KEYINPUT120), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1064 ( .A(KEYINPUT53), .B(n974), .Z(n978) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n975), .B(G34), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(G2084), .B(n976), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G35), .B(G2090), .ZN(n979) );
  NOR2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(n981), .B(KEYINPUT122), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n982), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(KEYINPUT55), .B(n983), .ZN(n984) );
  NAND2_X1 U1074 ( .A1(n984), .A2(G11), .ZN(n1038) );
  XNOR2_X1 U1075 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(n987), .B(KEYINPUT57), .ZN(n1006) );
  XNOR2_X1 U1079 ( .A(G171), .B(G1961), .ZN(n1001) );
  XNOR2_X1 U1080 ( .A(G299), .B(G1956), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n988), .B(G1341), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n999) );
  AND2_X1 U1084 ( .A1(G303), .A2(G1971), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(KEYINPUT123), .B(n997), .ZN(n998) );
  NOR2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(G1348), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1036) );
  INV_X1 U1094 ( .A(G16), .ZN(n1034) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G22), .B(G1971), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT126), .B(n1011), .Z(n1013) );
  XNOR2_X1 U1099 ( .A(G1986), .B(G24), .ZN(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1014), .ZN(n1018) );
  XNOR2_X1 U1102 ( .A(G1966), .B(G21), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G5), .B(G1961), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1030) );
  XNOR2_X1 U1106 ( .A(KEYINPUT59), .B(G1348), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(n1019), .B(G4), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(G1981), .B(G6), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(G19), .B(G1341), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1111 ( .A(KEYINPUT124), .B(n1022), .Z(n1024) );
  XNOR2_X1 U1112 ( .A(G1956), .B(G20), .ZN(n1023) );
  NOR2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1115 ( .A(KEYINPUT60), .B(n1027), .Z(n1028) );
  XNOR2_X1 U1116 ( .A(KEYINPUT125), .B(n1028), .ZN(n1029) );
  NOR2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1118 ( .A(n1031), .B(KEYINPUT61), .Z(n1032) );
  XNOR2_X1 U1119 ( .A(KEYINPUT127), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1122 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1123 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1124 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1125 ( .A(G311), .ZN(G150) );
endmodule

