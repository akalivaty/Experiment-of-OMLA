//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1256, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT64), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n215), .A2(G1), .A3(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n207), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT65), .B(G244), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(G77), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n222), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  NAND2_X1  g0040(.A1(G68), .A2(G77), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n203), .A2(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n242), .B(KEYINPUT66), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  OAI21_X1  g0049(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NOR3_X1   g0053(.A1(new_n252), .A2(new_n253), .A3(new_n213), .ZN(new_n254));
  AND2_X1   g0054(.A1(G1), .A2(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT67), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(G274), .B(new_n251), .C1(new_n254), .C2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n253), .B1(new_n252), .B2(new_n213), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n255), .A2(KEYINPUT67), .A3(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n250), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT68), .B(G226), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n258), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT69), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G222), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(G1698), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  OAI221_X1 g0071(.A(new_n269), .B1(new_n202), .B2(new_n267), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n252), .B1(new_n214), .B2(new_n216), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n264), .A2(new_n265), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n266), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n266), .A2(KEYINPUT70), .A3(new_n274), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(G200), .A3(new_n279), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n214), .A2(new_n216), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT71), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT71), .ZN(new_n289));
  INV_X1    g0089(.A(G58), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(KEYINPUT8), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n207), .A2(G33), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G50), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(new_n290), .A3(new_n201), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n296), .A2(G20), .B1(G150), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n286), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n285), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n206), .A2(G20), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(G50), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G50), .B2(new_n300), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g0106(.A(new_n306), .B(KEYINPUT9), .Z(new_n307));
  OAI211_X1 g0107(.A(new_n283), .B(new_n307), .C1(KEYINPUT74), .C2(KEYINPUT10), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n281), .A2(KEYINPUT74), .A3(new_n282), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n281), .A2(new_n307), .A3(new_n282), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT10), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n280), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n306), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n278), .A2(new_n316), .A3(new_n279), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n308), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  XOR2_X1   g0119(.A(KEYINPUT77), .B(KEYINPUT14), .Z(new_n320));
  INV_X1    g0120(.A(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G33), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n322), .A2(new_n324), .A3(G232), .A4(G1698), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n322), .A2(new_n324), .A3(G226), .A4(new_n268), .ZN(new_n326));
  NAND2_X1  g0126(.A1(G33), .A2(G97), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT75), .A4(new_n327), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n273), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n251), .B1(new_n259), .B2(new_n260), .ZN(new_n334));
  INV_X1    g0134(.A(G274), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n335), .B1(new_n259), .B2(new_n260), .ZN(new_n336));
  AOI22_X1  g0136(.A1(G238), .A2(new_n334), .B1(new_n336), .B2(new_n251), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n332), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n333), .B1(new_n332), .B2(new_n337), .ZN(new_n340));
  OAI211_X1 g0140(.A(G169), .B(new_n320), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n332), .A2(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n343), .A2(G179), .A3(new_n338), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  OAI21_X1  g0146(.A(G169), .B1(new_n339), .B2(new_n340), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n346), .B1(new_n347), .B2(KEYINPUT76), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n316), .B1(new_n343), .B2(new_n338), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n345), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n201), .A2(G20), .ZN(new_n353));
  INV_X1    g0153(.A(new_n297), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n353), .B1(new_n293), .B2(new_n202), .C1(new_n354), .C2(new_n295), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n285), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT11), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT72), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n300), .B(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(new_n285), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n360), .A2(G68), .A3(new_n303), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G13), .ZN(new_n363));
  NOR4_X1   g0163(.A1(new_n353), .A2(KEYINPUT12), .A3(G1), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n359), .A2(new_n201), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(KEYINPUT12), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n352), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G200), .B1(new_n339), .B2(new_n340), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n343), .A2(G190), .A3(new_n338), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT7), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n267), .A2(new_n374), .A3(G20), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n322), .A2(new_n324), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT7), .B1(new_n376), .B2(new_n207), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n290), .A2(new_n201), .ZN(new_n379));
  NOR2_X1   g0179(.A1(G58), .A2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n297), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n378), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT16), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n374), .B1(new_n267), .B2(G20), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n376), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n201), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n386), .B1(new_n389), .B2(new_n383), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(new_n390), .A3(new_n285), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n292), .B1(new_n206), .B2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n302), .B1(new_n301), .B2(new_n292), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n271), .A2(new_n268), .ZN(new_n394));
  INV_X1    g0194(.A(G226), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G1698), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n322), .A2(new_n394), .A3(new_n324), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT78), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(KEYINPUT78), .A3(new_n398), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n273), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G190), .ZN(new_n404));
  AOI22_X1  g0204(.A1(G232), .A2(new_n334), .B1(new_n336), .B2(new_n251), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(G200), .B1(new_n403), .B2(new_n405), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n391), .B(new_n393), .C1(new_n406), .C2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT79), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n405), .A3(new_n404), .ZN(new_n410));
  OAI211_X1 g0210(.A(G232), .B(new_n250), .C1(new_n254), .C2(new_n257), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n258), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n217), .A2(new_n256), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G223), .A2(G1698), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n395), .B2(G1698), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n267), .B1(G33), .B2(G87), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n413), .B1(new_n416), .B2(KEYINPUT78), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n412), .B1(new_n401), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n410), .B1(new_n418), .B2(G200), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n391), .A4(new_n393), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n419), .A2(new_n423), .A3(new_n391), .A4(new_n393), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT80), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(G169), .B1(new_n403), .B2(new_n405), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n313), .B2(new_n418), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n391), .A2(new_n393), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n433), .B1(new_n429), .B2(new_n430), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n409), .A2(KEYINPUT80), .A3(KEYINPUT17), .A4(new_n421), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n427), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n438));
  INV_X1    g0238(.A(G107), .ZN(new_n439));
  INV_X1    g0239(.A(G238), .ZN(new_n440));
  OAI221_X1 g0240(.A(new_n438), .B1(new_n439), .B2(new_n267), .C1(new_n270), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n273), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n334), .A2(new_n223), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n258), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G200), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n404), .B2(new_n444), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G20), .A2(G77), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT15), .B(G87), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n447), .B1(new_n287), .B2(new_n354), .C1(new_n293), .C2(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n285), .B1(new_n202), .B2(new_n359), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n360), .A2(G77), .A3(new_n303), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT73), .ZN(new_n453));
  XNOR2_X1  g0253(.A(new_n452), .B(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n444), .A2(new_n316), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n444), .A2(G179), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NOR4_X1   g0259(.A1(new_n319), .A2(new_n373), .A3(new_n437), .A4(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n363), .A2(G1), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n207), .A2(G107), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n464));
  OR2_X1    g0264(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n465));
  NAND2_X1  g0265(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n461), .A2(new_n462), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n206), .A2(G33), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n302), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n439), .A2(KEYINPUT23), .A3(G20), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT23), .B1(new_n439), .B2(G20), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n322), .A2(new_n324), .A3(new_n207), .A4(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT22), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n267), .A2(new_n478), .A3(new_n207), .A4(G87), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n285), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n481), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n483), .B(new_n475), .C1(new_n477), .C2(new_n479), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n471), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n322), .A2(new_n324), .A3(G257), .A4(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n322), .A2(new_n324), .A3(G250), .A4(new_n268), .ZN(new_n488));
  INV_X1    g0288(.A(G294), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(new_n321), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n273), .ZN(new_n491));
  OR2_X1    g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NAND2_X1  g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G45), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G1), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n259), .A2(new_n260), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G264), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n206), .A2(G45), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n492), .B2(new_n493), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n500), .B(G274), .C1(new_n254), .C2(new_n257), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n491), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G200), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n490), .A2(new_n273), .B1(new_n497), .B2(G264), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(new_n404), .A3(new_n501), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n461), .A2(new_n358), .A3(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n206), .B2(G33), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n286), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n359), .A2(new_n511), .ZN(new_n514));
  AOI21_X1  g0314(.A(G20), .B1(G33), .B2(G283), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n321), .A2(G97), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n515), .A2(new_n516), .B1(G20), .B2(new_n511), .ZN(new_n517));
  AND3_X1   g0317(.A1(new_n517), .A2(new_n285), .A3(KEYINPUT20), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT20), .B1(new_n517), .B2(new_n285), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n513), .B(new_n514), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n322), .A2(new_n324), .A3(G264), .A4(G1698), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n322), .A2(new_n324), .A3(G257), .A4(new_n268), .ZN(new_n522));
  XOR2_X1   g0322(.A(KEYINPUT84), .B(G303), .Z(new_n523));
  OAI211_X1 g0323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n267), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n273), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n497), .A2(G270), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(new_n501), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n520), .B1(new_n527), .B2(G200), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n497), .A2(G270), .B1(new_n336), .B2(new_n500), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(G190), .A3(new_n525), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n486), .A2(new_n507), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n322), .A2(new_n324), .A3(G244), .A4(new_n268), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n267), .A2(KEYINPUT4), .A3(G244), .A4(new_n268), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G283), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n267), .A2(G250), .A3(G1698), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n273), .ZN(new_n539));
  INV_X1    g0339(.A(new_n493), .ZN(new_n540));
  NOR2_X1   g0340(.A1(KEYINPUT5), .A2(G41), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n496), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G257), .B(new_n542), .C1(new_n254), .C2(new_n257), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n501), .A2(new_n543), .A3(KEYINPUT81), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT81), .B1(new_n501), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G200), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n300), .A2(G97), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n470), .B2(G97), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT6), .ZN(new_n550));
  INV_X1    g0350(.A(G97), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n550), .A2(new_n551), .A3(G107), .ZN(new_n552));
  XNOR2_X1  g0352(.A(G97), .B(G107), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  OAI22_X1  g0354(.A1(new_n554), .A2(new_n207), .B1(new_n202), .B2(new_n354), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n439), .B1(new_n387), .B2(new_n388), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n285), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n501), .A2(new_n543), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n273), .B2(new_n538), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(G190), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n501), .A2(new_n543), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n539), .A2(new_n564), .A3(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT82), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n547), .A2(new_n559), .A3(new_n563), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n539), .A2(new_n564), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n316), .A2(new_n568), .B1(new_n549), .B2(new_n557), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n313), .B(new_n539), .C1(new_n544), .C2(new_n545), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n531), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n440), .A2(new_n268), .ZN(new_n574));
  INV_X1    g0374(.A(G244), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G1698), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n322), .A2(new_n574), .A3(new_n324), .A4(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n413), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(G250), .B1(new_n206), .B2(G45), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(new_n335), .B2(new_n496), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n261), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(G200), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n207), .B1(new_n327), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G87), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n551), .A3(new_n439), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n322), .A2(new_n324), .A3(new_n207), .A4(G68), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n584), .B1(new_n293), .B2(new_n551), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n591), .A2(new_n285), .B1(new_n359), .B2(new_n448), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n286), .A2(G87), .A3(new_n300), .A4(new_n469), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n582), .A2(new_n583), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n285), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n359), .A2(new_n448), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n577), .A2(new_n573), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n273), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n261), .A2(new_n580), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n503), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT83), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(G190), .A3(new_n600), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n594), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n316), .B1(new_n578), .B2(new_n581), .ZN(new_n605));
  INV_X1    g0405(.A(new_n448), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n302), .A2(new_n606), .A3(new_n469), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n595), .A3(new_n596), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n598), .A2(new_n273), .B1(new_n261), .B2(new_n580), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n313), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n605), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n604), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n502), .A2(new_n316), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n505), .A2(new_n313), .A3(new_n501), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n485), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n527), .A2(new_n520), .A3(G169), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n520), .A2(G179), .A3(new_n525), .A4(new_n529), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n527), .A2(new_n520), .A3(KEYINPUT21), .A4(G169), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n615), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n572), .A2(new_n612), .A3(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n460), .A2(new_n622), .ZN(G372));
  INV_X1    g0423(.A(KEYINPUT89), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT88), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n619), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n316), .B1(new_n529), .B2(new_n525), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT21), .B1(new_n627), .B2(new_n520), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n618), .A2(KEYINPUT88), .A3(new_n619), .A4(new_n620), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n624), .B1(new_n631), .B2(new_n615), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n485), .A2(new_n613), .A3(new_n614), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT89), .B(new_n633), .C1(new_n629), .C2(new_n630), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n582), .A2(new_n592), .A3(new_n593), .A4(new_n603), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n611), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n611), .A3(KEYINPUT87), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n486), .B2(new_n507), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n565), .B(new_n562), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n558), .B1(G200), .B2(new_n546), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n641), .A2(new_n642), .B1(new_n570), .B2(new_n569), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n632), .A2(new_n634), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n611), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n568), .A2(new_n316), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n648), .A2(new_n570), .A3(new_n558), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n635), .A2(new_n611), .A3(KEYINPUT87), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT87), .B1(new_n635), .B2(new_n611), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT90), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n604), .A2(new_n570), .A3(new_n569), .A4(new_n611), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(new_n654), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n653), .B1(new_n652), .B2(new_n654), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n647), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n646), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n460), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n318), .ZN(new_n664));
  INV_X1    g0464(.A(new_n458), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n368), .B1(new_n372), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n427), .A2(new_n436), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n435), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n308), .A2(new_n312), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n664), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n461), .A2(new_n207), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT91), .Z(new_n673));
  INV_X1    g0473(.A(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n672), .B(KEYINPUT91), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(G213), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(KEYINPUT92), .B(G343), .Z(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n520), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n629), .B2(new_n630), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n528), .A2(new_n530), .ZN(new_n683));
  INV_X1    g0483(.A(new_n681), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n626), .A2(new_n628), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT93), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n486), .A2(new_n507), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n680), .A2(new_n485), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n633), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n615), .A2(new_n680), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n688), .A2(G330), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n685), .A2(new_n680), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n692), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n210), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n587), .A2(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n220), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n640), .A2(new_n643), .A3(new_n621), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n656), .A2(new_n654), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT26), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n708), .A3(new_n611), .ZN(new_n709));
  INV_X1    g0509(.A(new_n680), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(KEYINPUT29), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n680), .B1(new_n646), .B2(new_n661), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(KEYINPUT29), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n609), .A2(G179), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT95), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n546), .A2(new_n715), .A3(new_n502), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n715), .B1(new_n546), .B2(new_n502), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n527), .B(new_n714), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT94), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n505), .A2(new_n539), .A3(new_n564), .A4(new_n609), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n529), .A2(G179), .A3(new_n525), .ZN(new_n723));
  OAI211_X1 g0523(.A(new_n720), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n723), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n505), .A2(new_n609), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n720), .A2(new_n721), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n726), .A3(new_n561), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n710), .B1(new_n719), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n621), .A2(new_n612), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n643), .A3(new_n531), .A4(new_n710), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n731), .B1(new_n733), .B2(KEYINPUT31), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n714), .A2(new_n527), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n546), .A2(new_n502), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT95), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n735), .B1(new_n737), .B2(new_n716), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT31), .B(new_n680), .C1(new_n738), .C2(new_n729), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(G330), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n713), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n704), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n363), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n206), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n699), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n688), .B2(G330), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n749), .B1(G330), .B2(new_n688), .ZN(new_n750));
  INV_X1    g0550(.A(new_n748), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n698), .A2(new_n376), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(G355), .B1(new_n511), .B2(new_n698), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n245), .A2(G45), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n698), .A2(new_n267), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G45), .B2(new_n220), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT96), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n753), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT97), .Z(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n218), .B1(G20), .B2(new_n316), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n751), .B1(new_n758), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n761), .ZN(new_n765));
  NOR4_X1   g0565(.A1(new_n207), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OR2_X1    g0567(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(KEYINPUT98), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT32), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n207), .A2(G179), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n503), .A2(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n207), .A2(new_n313), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n503), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n267), .B1(new_n776), .B2(new_n439), .C1(new_n780), .C2(new_n295), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n777), .A2(new_n775), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n777), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G68), .A2(new_n783), .B1(new_n786), .B2(G77), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(new_n586), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n778), .A2(G200), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n290), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n404), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n207), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n551), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n781), .A2(new_n789), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n773), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(KEYINPUT99), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n797), .A2(KEYINPUT99), .ZN(new_n799));
  INV_X1    g0599(.A(new_n770), .ZN(new_n800));
  INV_X1    g0600(.A(new_n776), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n800), .A2(G329), .B1(G283), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT100), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n790), .A2(G322), .ZN(new_n804));
  INV_X1    g0604(.A(G326), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n780), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n267), .B1(new_n783), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G303), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(new_n809), .B2(new_n788), .C1(new_n810), .C2(new_n785), .ZN(new_n811));
  INV_X1    g0611(.A(new_n794), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n806), .B(new_n811), .C1(G294), .C2(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n798), .B(new_n799), .C1(new_n803), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n762), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n764), .B1(new_n687), .B2(new_n765), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n750), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  AOI22_X1  g0618(.A1(G150), .A2(new_n783), .B1(new_n786), .B2(G159), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n819), .B1(new_n780), .B2(new_n820), .C1(new_n821), .C2(new_n791), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT34), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n800), .A2(G132), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n776), .A2(new_n201), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n267), .B1(new_n788), .B2(new_n295), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G58), .C2(new_n812), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n824), .A2(new_n825), .A3(new_n826), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n780), .A2(new_n809), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n795), .B(new_n831), .C1(G294), .C2(new_n790), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n783), .A2(KEYINPUT101), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G283), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n800), .A2(G311), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n439), .A2(new_n788), .B1(new_n785), .B2(new_n511), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n267), .B(new_n839), .C1(G87), .C2(new_n801), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n832), .A2(new_n837), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n815), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n760), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n762), .A2(new_n843), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n751), .B(new_n842), .C1(new_n202), .C2(new_n844), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT102), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n458), .A2(new_n680), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n454), .A2(new_n680), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n455), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n847), .B1(new_n849), .B2(new_n458), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n846), .B1(new_n760), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n662), .A2(new_n710), .ZN(new_n852));
  INV_X1    g0652(.A(new_n850), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n741), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n655), .A2(new_n657), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n611), .B1(new_n856), .B2(new_n659), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n710), .B(new_n850), .C1(new_n857), .C2(new_n645), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n854), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT103), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT103), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n854), .A2(new_n861), .A3(new_n855), .A4(new_n858), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n860), .A2(KEYINPUT104), .A3(new_n751), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n854), .A2(new_n858), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n741), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n862), .A2(new_n751), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT104), .B1(new_n867), .B2(new_n860), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n851), .B1(new_n866), .B2(new_n868), .ZN(G384));
  NOR2_X1   g0669(.A1(new_n745), .A2(new_n206), .ZN(new_n870));
  INV_X1    g0670(.A(new_n678), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n430), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n437), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT105), .B1(new_n429), .B2(new_n430), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n429), .A2(KEYINPUT105), .A3(new_n430), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n409), .A3(new_n421), .A4(new_n879), .ZN(new_n880));
  AND4_X1   g0680(.A1(new_n431), .A2(new_n409), .A3(new_n421), .A4(new_n872), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(new_n875), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n874), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n874), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n369), .A2(new_n680), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n874), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n431), .A2(new_n408), .A3(new_n872), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n874), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n889), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n887), .B(new_n888), .C1(new_n894), .C2(KEYINPUT39), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n435), .A2(new_n871), .ZN(new_n896));
  INV_X1    g0696(.A(new_n367), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT14), .B1(new_n349), .B2(new_n350), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n347), .A2(KEYINPUT76), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n344), .B(new_n341), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n372), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n897), .B(new_n680), .C1(new_n900), .C2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n680), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n372), .B(new_n903), .C1(new_n352), .C2(new_n367), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n847), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n858), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n885), .A2(new_n886), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n896), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n895), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n460), .B(new_n711), .C1(KEYINPUT29), .C2(new_n712), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n670), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n910), .B(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(G330), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n853), .B1(new_n904), .B2(new_n902), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n739), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n719), .A2(new_n730), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n918), .A2(KEYINPUT106), .A3(KEYINPUT31), .A4(new_n680), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT31), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n622), .B2(new_n710), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n917), .B(new_n919), .C1(new_n921), .C2(new_n731), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT40), .B1(new_n894), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n902), .A2(new_n904), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n850), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n919), .A2(new_n917), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n734), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n908), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n460), .A2(new_n922), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n914), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n933), .B2(new_n932), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n870), .B1(new_n913), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n913), .B2(new_n935), .ZN(new_n937));
  INV_X1    g0737(.A(new_n554), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n938), .A2(KEYINPUT35), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(KEYINPUT35), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n939), .A2(G116), .A3(new_n219), .A4(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT36), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n379), .A2(new_n220), .A3(new_n202), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n201), .A2(G50), .ZN(new_n944));
  OAI211_X1 g0744(.A(G1), .B(new_n363), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n937), .A2(new_n942), .A3(new_n945), .ZN(G367));
  OAI21_X1  g0746(.A(new_n763), .B1(new_n210), .B2(new_n448), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n239), .A2(new_n698), .A3(new_n267), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n748), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(G283), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n376), .B1(new_n776), .B2(new_n551), .C1(new_n950), .C2(new_n785), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n780), .A2(new_n810), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n788), .A2(new_n511), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n951), .B(new_n952), .C1(KEYINPUT46), .C2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(G317), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n954), .B1(new_n489), .B2(new_n835), .C1(new_n955), .C2(new_n770), .ZN(new_n956));
  INV_X1    g0756(.A(new_n523), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n790), .A2(new_n957), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n958), .B1(KEYINPUT46), .B2(new_n953), .C1(new_n439), .C2(new_n794), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n794), .A2(new_n201), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n788), .A2(new_n290), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n785), .A2(new_n295), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(G150), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n963), .B1(new_n821), .B2(new_n780), .C1(new_n964), .C2(new_n791), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n267), .B1(new_n776), .B2(new_n202), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT110), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n967), .B1(new_n820), .B2(new_n770), .C1(new_n771), .C2(new_n835), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n956), .A2(new_n959), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT47), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n949), .B1(new_n970), .B2(new_n762), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n680), .A2(new_n597), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n611), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n638), .A2(new_n639), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n973), .B1(new_n974), .B2(new_n972), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n761), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n699), .B(KEYINPUT41), .Z(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n688), .A2(G330), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n693), .B(new_n695), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT107), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n643), .B1(new_n559), .B2(new_n710), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n649), .A2(new_n680), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n696), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n985), .B1(new_n696), .B2(new_n988), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n984), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT44), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n696), .A2(new_n993), .A3(new_n988), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n696), .B2(new_n988), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n696), .A2(new_n988), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT107), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n992), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT108), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n694), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n694), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n983), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n980), .B1(new_n1005), .B2(new_n742), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT109), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n983), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1004), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1009), .B1(new_n1010), .B2(new_n1002), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n743), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1012), .A2(KEYINPUT109), .A3(new_n980), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n747), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n988), .A2(new_n693), .A3(new_n695), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n571), .B1(new_n986), .B2(new_n615), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n1015), .A2(KEYINPUT42), .B1(new_n1016), .B2(new_n710), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(KEYINPUT42), .B2(new_n1015), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT43), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n975), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n975), .A2(new_n1019), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1020), .B(new_n1021), .Z(new_n1022));
  AOI21_X1  g0822(.A(new_n694), .B1(new_n986), .B2(new_n987), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n978), .B1(new_n1014), .B2(new_n1025), .ZN(G387));
  INV_X1    g0826(.A(new_n701), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n752), .A2(new_n1027), .B1(new_n439), .B2(new_n698), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n236), .A2(new_n495), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n287), .A2(G50), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT50), .Z(new_n1031));
  NAND3_X1  g0831(.A1(new_n701), .A2(new_n495), .A3(new_n241), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n755), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1028), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n751), .B1(new_n1034), .B2(new_n763), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n788), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G77), .A2(new_n1036), .B1(new_n786), .B2(G68), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n376), .B1(new_n801), .B2(G97), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1037), .B(new_n1038), .C1(new_n292), .C2(new_n782), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n812), .A2(new_n606), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n780), .B2(new_n771), .C1(new_n295), .C2(new_n791), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(G150), .C2(new_n800), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n779), .A2(G322), .B1(new_n957), .B2(new_n786), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n955), .B2(new_n791), .C1(new_n835), .C2(new_n810), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n812), .A2(G283), .B1(new_n1036), .B2(G294), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1050), .A2(KEYINPUT49), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n376), .B1(new_n511), .B2(new_n776), .C1(new_n770), .C2(new_n805), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n1050), .B2(KEYINPUT49), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1042), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1035), .B1(new_n693), .B2(new_n765), .C1(new_n1054), .C2(new_n815), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n743), .A2(new_n1009), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n699), .B1(new_n742), .B2(new_n983), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1055), .B1(new_n746), .B2(new_n983), .C1(new_n1056), .C2(new_n1057), .ZN(G393));
  XOR2_X1   g0858(.A(new_n1000), .B(new_n694), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1057), .B2(new_n746), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n763), .B1(new_n551), .B2(new_n210), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n755), .A2(new_n248), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n748), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n812), .A2(G77), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n287), .B2(new_n785), .C1(new_n835), .C2(new_n295), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT111), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G150), .A2(new_n779), .B1(new_n790), .B2(G159), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n376), .B1(new_n801), .B2(G87), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n201), .B2(new_n788), .C1(new_n770), .C2(new_n821), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT112), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G311), .A2(new_n790), .B1(new_n779), .B2(G317), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI21_X1  g0875(.A(new_n376), .B1(new_n776), .B2(new_n439), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n950), .A2(new_n788), .B1(new_n785), .B2(new_n489), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G116), .C2(new_n812), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n836), .A2(new_n957), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n800), .A2(G322), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1075), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1072), .A2(KEYINPUT112), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1073), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1063), .B1(new_n1083), .B2(new_n762), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n765), .B2(new_n988), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n743), .A2(new_n699), .A3(new_n1009), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1060), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(G390));
  OAI21_X1  g0890(.A(new_n887), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n843), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n751), .B1(new_n844), .B2(new_n292), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n267), .B1(new_n776), .B2(new_n295), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n800), .A2(G125), .B1(KEYINPUT116), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n820), .B2(new_n835), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n788), .A2(new_n964), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(KEYINPUT116), .B2(new_n1094), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G159), .A2(new_n812), .B1(new_n779), .B2(G128), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT54), .B(G143), .Z(new_n1101));
  AOI22_X1  g0901(.A1(new_n790), .A2(G132), .B1(new_n786), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1096), .A2(new_n1099), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n827), .B1(new_n800), .B2(G294), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT118), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n376), .B1(new_n785), .B2(new_n551), .C1(new_n586), .C2(new_n788), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1064), .B1(new_n780), .B2(new_n950), .C1(new_n511), .C2(new_n791), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(G107), .C2(new_n836), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1106), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1092), .B(new_n1093), .C1(new_n815), .C2(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n874), .A2(new_n892), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n884), .ZN(new_n1118));
  AOI21_X1  g0918(.A(KEYINPUT39), .B1(new_n1118), .B2(new_n886), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1116), .A2(new_n1119), .B1(new_n907), .B2(new_n888), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n849), .A2(new_n458), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n709), .A2(new_n710), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n906), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT113), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT113), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1122), .A2(new_n1125), .A3(new_n906), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(new_n925), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT114), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n888), .B1(new_n1118), .B2(new_n886), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1128), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1120), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n915), .A2(new_n922), .A3(G330), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n855), .A2(new_n850), .A3(new_n925), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1120), .B(new_n1136), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1115), .B1(new_n1138), .B2(new_n746), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1138), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n741), .A2(new_n905), .A3(new_n853), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n1126), .B2(new_n1124), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n922), .A2(G330), .A3(new_n850), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n905), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n858), .A2(new_n906), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n905), .B1(new_n741), .B2(new_n853), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1133), .A2(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1142), .A2(new_n1144), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n460), .A2(G330), .A3(new_n922), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n911), .A2(new_n670), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT115), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n700), .B1(new_n1140), .B2(new_n1151), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n911), .A2(new_n670), .A3(new_n1149), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1122), .A2(new_n1125), .A3(new_n906), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1125), .B1(new_n1122), .B2(new_n906), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1144), .B(new_n1136), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1147), .A2(new_n1145), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1138), .A2(KEYINPUT115), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1139), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(G378));
  NOR2_X1   g0962(.A1(new_n306), .A2(new_n678), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT55), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(new_n319), .B(new_n1164), .ZN(new_n1165));
  XOR2_X1   g0965(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1166));
  XNOR2_X1  g0966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(new_n760), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n844), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(G33), .A2(G41), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1170), .A2(G50), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n267), .B2(G41), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G41), .B(new_n267), .C1(new_n1036), .C2(G77), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n290), .B2(new_n776), .C1(new_n770), .C2(new_n950), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT119), .Z(new_n1175));
  OAI22_X1  g0975(.A1(new_n551), .A2(new_n782), .B1(new_n785), .B2(new_n448), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n791), .A2(new_n439), .B1(new_n780), .B2(new_n511), .ZN(new_n1177));
  NOR4_X1   g0977(.A1(new_n1175), .A2(new_n960), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1172), .B1(new_n1178), .B2(KEYINPUT58), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1179), .A2(KEYINPUT120), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(KEYINPUT120), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G150), .A2(new_n812), .B1(new_n790), .B2(G128), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1036), .A2(new_n1101), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G132), .A2(new_n783), .B1(new_n786), .B2(G137), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n779), .A2(G125), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  INV_X1    g0987(.A(G124), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1170), .B1(new_n771), .B2(new_n776), .C1(new_n770), .C2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n1186), .B2(KEYINPUT59), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1178), .A2(KEYINPUT58), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1180), .A2(new_n1181), .A3(new_n1191), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n748), .B1(G50), .B2(new_n1169), .C1(new_n1192), .C2(new_n815), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1168), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT38), .B1(new_n874), .B2(new_n882), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n930), .B1(new_n889), .B2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(new_n923), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n437), .A2(new_n873), .B1(new_n880), .B2(new_n891), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n886), .B1(KEYINPUT38), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n930), .B1(new_n929), .B2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(G330), .B1(new_n1197), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n895), .A3(new_n909), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n914), .B1(new_n924), .B2(new_n931), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n910), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n1202), .A2(new_n1204), .A3(new_n1167), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1167), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1194), .B1(new_n1207), .B2(new_n747), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1154), .A2(new_n1155), .A3(new_n905), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n888), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1199), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT114), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1127), .A2(new_n1129), .A3(new_n1128), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1145), .A2(new_n925), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n1210), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1212), .A2(new_n1213), .B1(new_n1215), .B2(new_n1091), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1137), .B(new_n1158), .C1(new_n1216), .C2(new_n1133), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1153), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT122), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT122), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1220), .A3(new_n1153), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1222), .B2(new_n1207), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1205), .A2(new_n1206), .A3(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1217), .A2(new_n1220), .A3(new_n1153), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1220), .B1(new_n1217), .B2(new_n1153), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n699), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1208), .B1(new_n1223), .B2(new_n1229), .ZN(G375));
  NAND2_X1  g1030(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1159), .A2(new_n1231), .A3(new_n980), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n905), .A2(new_n843), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n748), .B1(new_n1169), .B2(G68), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n791), .A2(new_n820), .B1(new_n295), .B2(new_n794), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G132), .B2(new_n779), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n836), .A2(new_n1101), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n800), .A2(G128), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n771), .A2(new_n788), .B1(new_n785), .B2(new_n964), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n376), .B(new_n1239), .C1(G58), .C2(new_n801), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n551), .A2(new_n788), .B1(new_n785), .B2(new_n439), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n267), .B(new_n1242), .C1(G77), .C2(new_n801), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n511), .B2(new_n835), .C1(new_n809), .C2(new_n770), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1040), .B1(new_n780), .B2(new_n489), .C1(new_n950), .C2(new_n791), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1241), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1234), .B1(new_n1246), .B2(new_n762), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1158), .A2(new_n747), .B1(new_n1233), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1232), .A2(new_n1248), .ZN(G381));
  OR4_X1    g1049(.A1(G396), .A2(G390), .A3(G393), .A4(G381), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(G384), .A3(G387), .ZN(new_n1251));
  INV_X1    g1051(.A(G375), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1161), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n679), .A2(G213), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT123), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1252), .A2(new_n1161), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G407), .A2(new_n1256), .A3(G213), .ZN(G409));
  INV_X1    g1057(.A(new_n1254), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1153), .B2(new_n1158), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1153), .A2(new_n1158), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1259), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1264));
  OAI211_X1 g1064(.A(KEYINPUT125), .B(new_n1231), .C1(new_n1264), .C2(new_n1260), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n700), .B1(new_n1262), .B2(KEYINPUT60), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n1248), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT126), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(G384), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G384), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(KEYINPUT126), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1267), .A2(new_n1271), .A3(KEYINPUT126), .A4(new_n1248), .ZN(new_n1274));
  AND2_X1   g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1167), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1202), .A2(new_n1204), .A3(new_n1167), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n980), .A3(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1208), .B1(new_n1281), .B2(KEYINPUT124), .ZN(new_n1282));
  NOR3_X1   g1082(.A1(new_n1205), .A2(new_n1206), .A3(new_n979), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(KEYINPUT124), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1161), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G378), .B(new_n1208), .C1(new_n1223), .C2(new_n1229), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1258), .B(new_n1275), .C1(new_n1286), .C2(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT127), .B1(new_n1288), .B2(KEYINPUT63), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1278), .A2(new_n747), .A3(new_n1279), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1291), .B1(new_n1168), .B2(new_n1193), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n700), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1207), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1224), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1161), .B(new_n1292), .C1(new_n1293), .C2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1283), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT124), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1292), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G378), .B1(new_n1299), .B2(new_n1284), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1254), .B(new_n1290), .C1(new_n1296), .C2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT127), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT63), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1255), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(KEYINPUT63), .A3(new_n1290), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(G393), .B(new_n817), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT109), .B1(new_n1012), .B2(new_n980), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1007), .B(new_n979), .C1(new_n1011), .C2(new_n743), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n746), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1024), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G390), .B1(new_n1312), .B2(new_n978), .ZN(new_n1313));
  AOI211_X1 g1113(.A(new_n977), .B(new_n1089), .C1(new_n1311), .C2(new_n1024), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1308), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G387), .A2(new_n1089), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1312), .A2(new_n978), .A3(G390), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1307), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1315), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1254), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1255), .A2(G2897), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1290), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1258), .A2(G2897), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1323), .B1(new_n1290), .B2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1320), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1289), .A2(new_n1304), .A3(new_n1306), .A4(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1275), .A2(new_n1329), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1301), .A2(new_n1329), .B1(new_n1305), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1290), .A2(new_n1324), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1332), .B1(new_n1290), .B2(new_n1322), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1319), .B1(new_n1305), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1328), .B1(new_n1331), .B2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1327), .A2(new_n1335), .ZN(G405));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1161), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1275), .B1(new_n1338), .B2(new_n1296), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1337), .A2(new_n1290), .A3(new_n1287), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1339), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1328), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1341), .B(new_n1342), .ZN(G402));
endmodule


