//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n581, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT67), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n462), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n461), .B1(new_n463), .B2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n472), .A2(KEYINPUT69), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n464), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n470), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT70), .ZN(G160));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n466), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI221_X1 g059(.A(new_n484), .B1(new_n483), .B2(new_n482), .C1(G112), .C2(new_n473), .ZN(new_n485));
  XOR2_X1   g060(.A(new_n485), .B(KEYINPUT72), .Z(new_n486));
  NOR2_X1   g061(.A1(new_n470), .A2(new_n473), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n470), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT73), .Z(G162));
  NAND4_X1  g067(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT4), .A4(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(G102), .A2(G2104), .ZN(new_n494));
  AOI21_X1  g069(.A(G2105), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n462), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n473), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n462), .A2(G138), .A3(new_n473), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n500), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n507), .A2(KEYINPUT75), .A3(G651), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(KEYINPUT74), .A2(KEYINPUT6), .A3(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n505), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n510), .A2(new_n511), .B1(G88), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n501), .B1(new_n515), .B2(new_n516), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  INV_X1    g097(.A(new_n505), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n524));
  INV_X1    g099(.A(new_n519), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT76), .B(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n524), .B(new_n529), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(new_n530), .B1(G89), .B2(new_n517), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n505), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G651), .B1(new_n519), .B2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n517), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n505), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n519), .B2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n517), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n519), .A2(G53), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n519), .B2(G53), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT79), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n559), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(new_n562), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n515), .A2(new_n516), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n523), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT80), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT80), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n517), .A2(new_n569), .A3(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n505), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n568), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n564), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n578));
  NOR2_X1   g153(.A1(G171), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n541), .A2(KEYINPUT81), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G301));
  NAND2_X1  g157(.A1(new_n517), .A2(G87), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n519), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G288));
  AND2_X1   g161(.A1(new_n517), .A2(G86), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT82), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n505), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(new_n519), .B2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n505), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT84), .B(G47), .Z(new_n600));
  NAND2_X1  g175(.A1(new_n519), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n517), .A2(G85), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT85), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n603), .A2(KEYINPUT85), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(new_n523), .A2(G66), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n514), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n566), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n517), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G54), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n525), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n581), .B2(new_n619), .ZN(G284));
  OAI21_X1  g196(.A(new_n620), .B1(new_n581), .B2(new_n619), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n619), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G168), .B2(new_n619), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(G168), .B2(new_n619), .ZN(G280));
  NOR2_X1   g200(.A1(new_n525), .A2(new_n617), .ZN(new_n626));
  AOI211_X1 g201(.A(new_n626), .B(new_n611), .C1(new_n615), .C2(new_n614), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n548), .A2(new_n619), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n618), .A2(G559), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT86), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n630), .B1(new_n632), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n489), .A2(G135), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n635), .A2(new_n636), .B1(G123), .B2(new_n487), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n637), .B(new_n639), .C1(new_n636), .C2(new_n635), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT90), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2096), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n489), .A2(G2104), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT88), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2430), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT15), .B(G2435), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT14), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n656), .B(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(G14), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2067), .B(G2678), .Z(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT17), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2096), .B(G2100), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n676), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  XOR2_X1   g256(.A(G1961), .B(G1966), .Z(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT93), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n685), .B(new_n686), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(KEYINPUT93), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n681), .A2(new_n682), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(KEYINPUT20), .ZN(new_n694));
  INV_X1    g269(.A(new_n683), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n687), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n691), .A2(new_n693), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1991), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT94), .B(G1986), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n697), .B(new_n703), .ZN(G229));
  INV_X1    g279(.A(G29), .ZN(new_n705));
  NOR2_X1   g280(.A1(G164), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G27), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G2078), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n549), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n710), .B2(G19), .ZN(new_n712));
  INV_X1    g287(.A(G1341), .ZN(new_n713));
  INV_X1    g288(.A(G1961), .ZN(new_n714));
  NAND2_X1  g289(.A1(G171), .A2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G5), .B2(G16), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(G168), .A2(new_n710), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n710), .B2(G21), .ZN(new_n719));
  INV_X1    g294(.A(G1966), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n717), .B1(new_n705), .B2(new_n642), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AOI211_X1 g296(.A(new_n709), .B(new_n721), .C1(new_n720), .C2(new_n719), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n707), .A2(new_n708), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n705), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n705), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n726));
  INV_X1    g301(.A(G2090), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(KEYINPUT29), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(new_n728), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G2090), .ZN(new_n731));
  NAND4_X1  g306(.A1(new_n722), .A2(new_n723), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  OAI22_X1  g307(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT99), .ZN(new_n735));
  INV_X1    g310(.A(G28), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT30), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n735), .B1(new_n736), .B2(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(new_n705), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n737), .B(new_n739), .C1(KEYINPUT30), .C2(new_n736), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G29), .B2(G33), .ZN(new_n742));
  OR3_X1    g317(.A1(new_n741), .A2(G29), .A3(G33), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT25), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n489), .A2(G139), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n745), .B(new_n746), .C1(new_n473), .C2(new_n747), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n742), .B(new_n743), .C1(new_n748), .C2(new_n705), .ZN(new_n749));
  INV_X1    g324(.A(G2072), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n734), .B(new_n751), .C1(new_n750), .C2(new_n749), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n487), .A2(G129), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n489), .A2(G141), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT26), .Z(new_n757));
  NAND4_X1  g332(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT97), .ZN(new_n759));
  MUX2_X1   g334(.A(G32), .B(new_n759), .S(G29), .Z(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1996), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n760), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n705), .A2(G26), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n487), .A2(G128), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n489), .A2(G140), .ZN(new_n766));
  OR2_X1    g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(new_n705), .ZN(new_n771));
  MUX2_X1   g346(.A(new_n764), .B(new_n771), .S(KEYINPUT28), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n710), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n627), .B2(new_n710), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1348), .ZN(new_n776));
  NOR4_X1   g351(.A1(new_n752), .A2(new_n763), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n575), .B1(new_n560), .B2(new_n563), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT23), .B1(new_n778), .B2(new_n710), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n710), .A2(G20), .ZN(new_n780));
  MUX2_X1   g355(.A(new_n779), .B(KEYINPUT23), .S(new_n780), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1956), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(G1956), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT31), .B(G11), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n777), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n732), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n787), .A2(KEYINPUT24), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n705), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G160), .B2(new_n705), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G2084), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n710), .A2(G6), .ZN(new_n793));
  INV_X1    g368(.A(G305), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n710), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT32), .B(G1981), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n710), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n710), .ZN(new_n799));
  INV_X1    g374(.A(G1971), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n710), .A2(G23), .ZN(new_n802));
  INV_X1    g377(.A(G288), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(new_n710), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT33), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1976), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n797), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT34), .Z(new_n808));
  NAND2_X1  g383(.A1(new_n705), .A2(G25), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n489), .A2(G131), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT95), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n811), .A2(new_n812), .B1(G119), .B2(new_n487), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n809), .B1(new_n816), .B2(new_n705), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G24), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n607), .B2(G16), .ZN(new_n821));
  INV_X1    g396(.A(G1986), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n808), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n786), .B(new_n792), .C1(new_n825), .C2(new_n826), .ZN(G150));
  INV_X1    g402(.A(G150), .ZN(G311));
  NAND2_X1  g403(.A1(new_n517), .A2(G93), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n519), .A2(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n829), .B(new_n830), .C1(new_n514), .C2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n548), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n627), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT101), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n840), .B(new_n841), .C1(new_n839), .C2(new_n838), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n832), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT102), .ZN(G145));
  XNOR2_X1  g421(.A(G160), .B(new_n642), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT103), .ZN(new_n848));
  INV_X1    g423(.A(G162), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(KEYINPUT103), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(G162), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n748), .A2(new_n758), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n759), .B2(new_n748), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n857));
  NAND2_X1  g432(.A1(G114), .A2(G2104), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n473), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT4), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n498), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n495), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n769), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n856), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n813), .A2(new_n815), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n473), .A2(G118), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n466), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI221_X1 g445(.A(new_n870), .B1(new_n869), .B2(new_n868), .C1(G106), .C2(G2105), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n489), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n487), .A2(G130), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n867), .A2(new_n874), .ZN(new_n876));
  INV_X1    g451(.A(new_n646), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n875), .B2(new_n876), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(KEYINPUT105), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n878), .B2(new_n879), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n866), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n879), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n865), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n854), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  INV_X1    g463(.A(new_n882), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n889), .A2(new_n880), .A3(new_n865), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(new_n853), .A3(new_n850), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(new_n888), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g469(.A(new_n833), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n632), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(G299), .A2(new_n618), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n778), .A2(new_n627), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT41), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(G299), .A2(new_n618), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n778), .A2(new_n627), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n896), .A2(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT42), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT107), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n606), .ZN(new_n913));
  NAND2_X1  g488(.A1(G303), .A2(new_n803), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(G303), .A2(new_n803), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n913), .B(new_n604), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n914), .B(new_n918), .C1(new_n605), .C2(new_n606), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(G305), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n919), .A3(new_n794), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(KEYINPUT42), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n908), .B(new_n909), .C1(new_n924), .C2(KEYINPUT42), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n912), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n925), .B1(new_n912), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(G868), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n832), .A2(new_n619), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(G295));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n930), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g508(.A1(G286), .A2(G171), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n581), .A2(G286), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n833), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n934), .B(new_n895), .C1(G286), .C2(new_n581), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n933), .B1(new_n907), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n903), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n906), .A2(KEYINPUT108), .A3(new_n937), .A4(new_n938), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n940), .A2(new_n923), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(new_n888), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n897), .A2(new_n898), .A3(new_n905), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(KEYINPUT109), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n903), .A2(new_n899), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n945), .A2(KEYINPUT109), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n941), .B1(new_n949), .B2(new_n939), .ZN(new_n950));
  INV_X1    g525(.A(new_n923), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n944), .A2(KEYINPUT43), .A3(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n951), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n944), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AND4_X1   g533(.A1(new_n958), .A2(new_n952), .A3(new_n888), .A4(new_n943), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n955), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n943), .A2(new_n888), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT43), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n957), .B1(new_n965), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g541(.A1(new_n607), .A2(new_n822), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n863), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G40), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n972), .B1(new_n478), .B2(G2105), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n464), .A2(new_n973), .A3(new_n474), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n971), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n967), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT124), .B(KEYINPUT48), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n978), .B(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n816), .B(new_n818), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n758), .A2(G1996), .ZN(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n769), .B(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n982), .B(new_n984), .C1(new_n759), .C2(G1996), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n980), .B1(new_n977), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n977), .B2(G1996), .ZN(new_n989));
  INV_X1    g564(.A(new_n984), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n976), .B1(new_n758), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n976), .A2(KEYINPUT46), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n816), .A2(new_n818), .ZN(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT123), .Z(new_n997));
  OAI22_X1  g572(.A1(new_n997), .A2(new_n985), .B1(G2067), .B2(new_n769), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n976), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n987), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n592), .ZN(new_n1001));
  OAI21_X1  g576(.A(G1981), .B1(new_n1001), .B2(new_n587), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1002), .B1(G305), .B2(G1981), .ZN(new_n1003));
  NOR2_X1   g578(.A1(KEYINPUT112), .A2(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1384), .B1(new_n861), .B2(new_n862), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n974), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI221_X1 g584(.A(new_n1002), .B1(KEYINPUT112), .B2(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n1012));
  INV_X1    g587(.A(G1976), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1009), .B(new_n1012), .C1(new_n1013), .C2(G288), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1013), .A3(G288), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1011), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1006), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1022), .A2(new_n974), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G2090), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n971), .A2(new_n974), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1029), .B2(new_n800), .ZN(new_n1030));
  INV_X1    g605(.A(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT55), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1021), .A2(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1011), .A2(G1976), .A3(G288), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G305), .A2(G1981), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1009), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1034), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1033), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1021), .A2(new_n1039), .A3(KEYINPUT63), .A4(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT116), .B(G2084), .ZN(new_n1042));
  AND4_X1   g617(.A1(new_n974), .A2(new_n1022), .A3(new_n1024), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n974), .B1(new_n1006), .B2(KEYINPUT45), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT115), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n969), .A2(new_n970), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n974), .B(new_n1047), .C1(new_n1006), .C2(KEYINPUT45), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1043), .B1(new_n1049), .B2(new_n720), .ZN(new_n1050));
  OR3_X1    g625(.A1(new_n1050), .A2(new_n1031), .A3(G286), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1041), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT63), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1035), .B(new_n1038), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1058), .B1(G286), .B2(G8), .ZN(new_n1059));
  AOI211_X1 g634(.A(KEYINPUT119), .B(new_n1031), .C1(new_n531), .C2(new_n533), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1050), .B2(new_n1031), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT120), .B(new_n1061), .C1(new_n1050), .C2(new_n1031), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1064), .A2(KEYINPUT51), .A3(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1050), .A2(new_n1061), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1062), .A2(new_n1063), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n1072));
  OR3_X1    g647(.A1(new_n1049), .A2(new_n1072), .A3(G2078), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1028), .A2(new_n708), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1074), .A2(new_n1072), .B1(new_n714), .B2(new_n1025), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n581), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1066), .A2(new_n1079), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1071), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1041), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1007), .A2(G2067), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1025), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(new_n618), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n618), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1085), .A3(new_n627), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n971), .A2(new_n992), .A3(new_n974), .A4(new_n1027), .ZN(new_n1095));
  XOR2_X1   g670(.A(KEYINPUT58), .B(G1341), .Z(new_n1096));
  NAND2_X1  g671(.A1(new_n1007), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1098), .B2(new_n549), .ZN(new_n1099));
  AOI211_X1 g674(.A(KEYINPUT59), .B(new_n548), .C1(new_n1095), .C2(new_n1097), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1093), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(KEYINPUT57), .B1(new_n561), .B2(new_n557), .ZN(new_n1102));
  AOI22_X1  g677(.A1(G299), .A2(KEYINPUT57), .B1(new_n576), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1956), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1025), .A2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT56), .B(G2072), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n971), .A2(new_n974), .A3(new_n1027), .A4(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT61), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT61), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1103), .A2(new_n1105), .A3(new_n1110), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1092), .A2(new_n1101), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n1103), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1108), .B2(new_n1089), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1084), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1074), .A2(new_n1072), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1025), .A2(new_n714), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n971), .A2(new_n1027), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1072), .B(G2078), .C1(new_n475), .C2(KEYINPUT121), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n475), .A2(KEYINPUT121), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1121), .A2(new_n973), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1119), .A2(G301), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT54), .B1(new_n1125), .B2(KEYINPUT122), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1075), .A2(new_n1127), .A3(G301), .A4(new_n1124), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1077), .A3(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1073), .A2(new_n1075), .A3(G301), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n541), .B1(new_n1075), .B2(new_n1124), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT54), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1088), .A2(new_n618), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT60), .B1(new_n1135), .B2(new_n1089), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1136), .A3(new_n1093), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1116), .B(KEYINPUT118), .C1(new_n1137), .C2(new_n1112), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1118), .A2(new_n1133), .A3(new_n1070), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1081), .A2(new_n1083), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1034), .A2(KEYINPUT113), .ZN(new_n1141));
  XOR2_X1   g716(.A(new_n1141), .B(new_n1040), .Z(new_n1142));
  XNOR2_X1  g717(.A(new_n1021), .B(KEYINPUT114), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1057), .B1(new_n1140), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n986), .A2(new_n967), .ZN(new_n1146));
  NAND2_X1  g721(.A1(G290), .A2(G1986), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n977), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1000), .B1(new_n1145), .B2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g724(.A(G229), .ZN(new_n1151));
  NAND3_X1  g725(.A1(new_n663), .A2(G319), .A3(new_n679), .ZN(new_n1152));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n1153));
  OAI21_X1  g727(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g728(.A(new_n1154), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1155));
  AOI21_X1  g729(.A(new_n958), .B1(new_n944), .B2(new_n955), .ZN(new_n1156));
  OAI211_X1 g730(.A(new_n893), .B(new_n1155), .C1(new_n1156), .C2(new_n959), .ZN(G225));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1158));
  NAND2_X1  g732(.A1(G225), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g733(.A1(new_n964), .A2(KEYINPUT126), .A3(new_n893), .A4(new_n1155), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1159), .A2(new_n1160), .ZN(G308));
endmodule


